module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 ;
  assign n129 = x110 | x111 ;
  assign n130 = x108 | x109 ;
  assign n131 = n129 | n130 ;
  assign n132 = x104 | x105 ;
  assign n133 = x106 | x107 ;
  assign n134 = n132 | n133 ;
  assign n135 = n131 | n134 ;
  assign n136 = x102 | x103 ;
  assign n137 = x100 | x101 ;
  assign n138 = n136 | n137 ;
  assign n139 = x98 | x99 ;
  assign n140 = x96 | x97 ;
  assign n141 = n139 | n140 ;
  assign n142 = n138 | n141 ;
  assign n143 = n135 | n142 ;
  assign n144 = x124 | x125 ;
  assign n145 = x126 | x127 ;
  assign n146 = n144 | n145 ;
  assign n147 = x122 | x123 ;
  assign n148 = x120 | x121 ;
  assign n149 = n147 | n148 ;
  assign n150 = n146 | n149 ;
  assign n151 = x116 | x117 ;
  assign n152 = x118 | x119 ;
  assign n153 = n151 | n152 ;
  assign n154 = x112 | x113 ;
  assign n155 = x114 | x115 ;
  assign n156 = n154 | n155 ;
  assign n157 = n153 | n156 ;
  assign n158 = n150 | n157 ;
  assign n159 = n143 | n158 ;
  assign n160 = x82 | x83 ;
  assign n161 = x80 | x81 ;
  assign n162 = n160 | n161 ;
  assign n163 = x86 | x87 ;
  assign n164 = x84 | x85 ;
  assign n165 = n163 | n164 ;
  assign n166 = n162 | n165 ;
  assign n167 = x88 | x89 ;
  assign n168 = x90 | x91 ;
  assign n169 = n167 | n168 ;
  assign n170 = x92 | x93 ;
  assign n171 = x94 | x95 ;
  assign n172 = n170 | n171 ;
  assign n173 = n169 | n172 ;
  assign n174 = n166 | n173 ;
  assign n175 = x78 | x79 ;
  assign n176 = x76 | x77 ;
  assign n177 = n175 | n176 ;
  assign n178 = x72 | x73 ;
  assign n179 = x74 | x75 ;
  assign n180 = n178 | n179 ;
  assign n181 = n177 | n180 ;
  assign n182 = x70 | x71 ;
  assign n183 = x68 | x69 ;
  assign n184 = n182 | n183 ;
  assign n185 = x66 | x67 ;
  assign n186 = x64 | x65 ;
  assign n187 = n185 | n186 ;
  assign n188 = n184 | n187 ;
  assign n189 = n181 | n188 ;
  assign n190 = n174 | n189 ;
  assign n191 = n159 | n190 ;
  assign n192 = x62 | x63 ;
  assign n193 = x60 | x61 ;
  assign n194 = n192 | n193 ;
  assign n195 = x56 | x57 ;
  assign n196 = x58 | x59 ;
  assign n197 = n195 | n196 ;
  assign n198 = n194 | n197 ;
  assign n199 = x50 | x51 ;
  assign n200 = x48 | x49 ;
  assign n201 = n199 | n200 ;
  assign n202 = x52 | x53 ;
  assign n203 = x54 | x55 ;
  assign n204 = n202 | n203 ;
  assign n205 = n201 | n204 ;
  assign n206 = n198 | n205 ;
  assign n207 = x36 | x37 ;
  assign n208 = x38 | x39 ;
  assign n209 = n207 | n208 ;
  assign n210 = x34 | x35 ;
  assign n211 = x32 | x33 ;
  assign n212 = n210 | n211 ;
  assign n213 = n209 | n212 ;
  assign n214 = x46 | x47 ;
  assign n215 = x44 | x45 ;
  assign n216 = n214 | n215 ;
  assign n217 = x42 | x43 ;
  assign n218 = x40 | x41 ;
  assign n219 = n217 | n218 ;
  assign n220 = n216 | n219 ;
  assign n221 = n213 | n220 ;
  assign n222 = n206 | n221 ;
  assign n223 = n191 | n222 ;
  assign n224 = x28 | x29 ;
  assign n225 = x30 | x31 ;
  assign n226 = n224 | n225 ;
  assign n227 = x24 | x25 ;
  assign n228 = x26 | x27 ;
  assign n229 = n227 | n228 ;
  assign n230 = n226 | n229 ;
  assign n231 = x18 | x19 ;
  assign n232 = x16 | x17 ;
  assign n233 = n231 | n232 ;
  assign n234 = x22 | x23 ;
  assign n235 = x20 | x21 ;
  assign n236 = n234 | n235 ;
  assign n237 = n233 | n236 ;
  assign n238 = n230 | n237 ;
  assign n239 = n223 | n238 ;
  assign n240 = x12 | x13 ;
  assign n241 = x14 | x15 ;
  assign n242 = n240 | n241 ;
  assign n243 = x8 | x9 ;
  assign n244 = x10 | x11 ;
  assign n245 = n243 | n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = x4 | x5 ;
  assign n248 = x6 | x7 ;
  assign n249 = n247 | n248 ;
  assign n250 = x2 | x3 ;
  assign n251 = x0 | x1 ;
  assign n252 = n250 | n251 ;
  assign n253 = n249 | n252 ;
  assign n254 = n246 | n253 ;
  assign n255 = n239 | n254 ;
  assign n256 = x1 & ~n250 ;
  assign n257 = ( x3 & ~n247 ) | ( x3 & n256 ) | ( ~n247 & n256 ) ;
  assign n258 = ( x5 & ~x6 ) | ( x5 & n257 ) | ( ~x6 & n257 ) ;
  assign n259 = x7 | n258 ;
  assign n260 = x9 & ~n244 ;
  assign n261 = ( x11 & ~n240 ) | ( x11 & n260 ) | ( ~n240 & n260 ) ;
  assign n262 = ( x13 & ~x14 ) | ( x13 & n261 ) | ( ~x14 & n261 ) ;
  assign n263 = n246 & ~n262 ;
  assign n264 = ( n259 & n262 ) | ( n259 & ~n263 ) | ( n262 & ~n263 ) ;
  assign n265 = x15 | n264 ;
  assign n266 = ~n239 & n265 ;
  assign n267 = x121 & ~n147 ;
  assign n268 = ( x123 & ~n144 ) | ( x123 & n267 ) | ( ~n144 & n267 ) ;
  assign n269 = ( x125 & ~x126 ) | ( x125 & n268 ) | ( ~x126 & n268 ) ;
  assign n270 = x127 | n269 ;
  assign n271 = x113 & ~n155 ;
  assign n272 = ( x115 & ~n151 ) | ( x115 & n271 ) | ( ~n151 & n271 ) ;
  assign n273 = ( x117 & ~x118 ) | ( x117 & n272 ) | ( ~x118 & n272 ) ;
  assign n274 = x119 | n273 ;
  assign n275 = ~n150 & n274 ;
  assign n276 = n270 | n275 ;
  assign n277 = x25 & ~n228 ;
  assign n278 = ( x27 & ~n224 ) | ( x27 & n277 ) | ( ~n224 & n277 ) ;
  assign n279 = ( x29 & ~x30 ) | ( x29 & n278 ) | ( ~x30 & n278 ) ;
  assign n280 = x31 | n279 ;
  assign n281 = x17 & ~n231 ;
  assign n282 = ( x19 & ~n235 ) | ( x19 & n281 ) | ( ~n235 & n281 ) ;
  assign n283 = ( x21 & ~x22 ) | ( x21 & n282 ) | ( ~x22 & n282 ) ;
  assign n284 = x23 | n283 ;
  assign n285 = ~n230 & n284 ;
  assign n286 = n280 | n285 ;
  assign n287 = ~n223 & n286 ;
  assign n288 = n276 | n287 ;
  assign n289 = n266 | n288 ;
  assign n290 = x65 & ~n185 ;
  assign n291 = ( x67 & ~n183 ) | ( x67 & n290 ) | ( ~n183 & n290 ) ;
  assign n292 = ( x69 & ~x70 ) | ( x69 & n291 ) | ( ~x70 & n291 ) ;
  assign n293 = x71 | n292 ;
  assign n294 = ~n181 & n293 ;
  assign n295 = x73 & ~n179 ;
  assign n296 = ( x75 & ~n176 ) | ( x75 & n295 ) | ( ~n176 & n295 ) ;
  assign n297 = ( x77 & ~x78 ) | ( x77 & n296 ) | ( ~x78 & n296 ) ;
  assign n298 = x79 | n297 ;
  assign n299 = n166 | n298 ;
  assign n300 = n294 | n299 ;
  assign n301 = ( ~x81 & n160 ) | ( ~x81 & n162 ) | ( n160 & n162 ) ;
  assign n302 = ( ~x83 & n164 ) | ( ~x83 & n301 ) | ( n164 & n301 ) ;
  assign n303 = ( ~x85 & n163 ) | ( ~x85 & n302 ) | ( n163 & n302 ) ;
  assign n304 = ( ~x87 & n173 ) | ( ~x87 & n303 ) | ( n173 & n303 ) ;
  assign n305 = n300 & ~n304 ;
  assign n306 = x57 & ~n196 ;
  assign n307 = ( x59 & ~n193 ) | ( x59 & n306 ) | ( ~n193 & n306 ) ;
  assign n308 = ( x61 & ~x62 ) | ( x61 & n307 ) | ( ~x62 & n307 ) ;
  assign n309 = x63 | n308 ;
  assign n310 = ~n190 & n309 ;
  assign n311 = x89 & ~n168 ;
  assign n312 = ( x91 & ~n170 ) | ( x91 & n311 ) | ( ~n170 & n311 ) ;
  assign n313 = ( x93 & ~x94 ) | ( x93 & n312 ) | ( ~x94 & n312 ) ;
  assign n314 = x95 | n313 ;
  assign n315 = n310 | n314 ;
  assign n316 = n305 | n315 ;
  assign n317 = ~n159 & n316 ;
  assign n318 = x33 & ~n210 ;
  assign n319 = ( x35 & ~n207 ) | ( x35 & n318 ) | ( ~n207 & n318 ) ;
  assign n320 = ( x37 & ~x38 ) | ( x37 & n319 ) | ( ~x38 & n319 ) ;
  assign n321 = x39 | n320 ;
  assign n322 = ~n220 & n321 ;
  assign n323 = x41 & ~n217 ;
  assign n324 = ( x43 & ~n215 ) | ( x43 & n323 ) | ( ~n215 & n323 ) ;
  assign n325 = ( x45 & ~x46 ) | ( x45 & n324 ) | ( ~x46 & n324 ) ;
  assign n326 = x47 | n325 ;
  assign n327 = ~n205 & n326 ;
  assign n328 = ( ~n205 & n322 ) | ( ~n205 & n327 ) | ( n322 & n327 ) ;
  assign n329 = x49 & ~n199 ;
  assign n330 = ( x51 & ~n202 ) | ( x51 & n329 ) | ( ~n202 & n329 ) ;
  assign n331 = ( x53 & ~x54 ) | ( x53 & n330 ) | ( ~x54 & n330 ) ;
  assign n332 = x55 | n331 ;
  assign n333 = n328 | n332 ;
  assign n334 = n191 | n198 ;
  assign n335 = n333 & ~n334 ;
  assign n336 = n317 | n335 ;
  assign n337 = n289 | n336 ;
  assign n338 = x97 & ~n139 ;
  assign n339 = ( x99 & ~n137 ) | ( x99 & n338 ) | ( ~n137 & n338 ) ;
  assign n340 = ( x101 & ~x102 ) | ( x101 & n339 ) | ( ~x102 & n339 ) ;
  assign n341 = x103 | n340 ;
  assign n342 = ~n135 & n341 ;
  assign n343 = x105 & ~n133 ;
  assign n344 = ( x107 & ~n130 ) | ( x107 & n343 ) | ( ~n130 & n343 ) ;
  assign n345 = ( x109 & ~x110 ) | ( x109 & n344 ) | ( ~x110 & n344 ) ;
  assign n346 = x111 | n345 ;
  assign n347 = ~n158 & n346 ;
  assign n348 = ( ~n158 & n342 ) | ( ~n158 & n347 ) | ( n342 & n347 ) ;
  assign n349 = n337 | n348 ;
  assign n350 = ~n215 & n217 ;
  assign n351 = n214 | n350 ;
  assign n352 = ~n209 & n210 ;
  assign n353 = ( n208 & ~n220 ) | ( n208 & n352 ) | ( ~n220 & n352 ) ;
  assign n354 = n351 | n353 ;
  assign n355 = ~n206 & n354 ;
  assign n356 = n199 & ~n204 ;
  assign n357 = ( ~n195 & n203 ) | ( ~n195 & n356 ) | ( n203 & n356 ) ;
  assign n358 = n196 | n357 ;
  assign n359 = ~n192 & n193 ;
  assign n360 = ( n192 & n358 ) | ( n192 & ~n359 ) | ( n358 & ~n359 ) ;
  assign n361 = n355 | n360 ;
  assign n362 = ~n191 & n361 ;
  assign n363 = ~n144 & n147 ;
  assign n364 = n145 | n363 ;
  assign n365 = n231 & ~n236 ;
  assign n366 = ( ~n229 & n234 ) | ( ~n229 & n365 ) | ( n234 & n365 ) ;
  assign n367 = ( ~n224 & n228 ) | ( ~n224 & n366 ) | ( n228 & n366 ) ;
  assign n368 = ( n225 & n364 ) | ( n225 & ~n367 ) | ( n364 & ~n367 ) ;
  assign n369 = n367 | n368 ;
  assign n370 = ( ~n223 & n364 ) | ( ~n223 & n369 ) | ( n364 & n369 ) ;
  assign n371 = n362 | n370 ;
  assign n372 = ~n249 & n250 ;
  assign n373 = ( ~n245 & n248 ) | ( ~n245 & n372 ) | ( n248 & n372 ) ;
  assign n374 = ( ~n242 & n244 ) | ( ~n242 & n373 ) | ( n244 & n373 ) ;
  assign n375 = ( ~n239 & n241 ) | ( ~n239 & n374 ) | ( n241 & n374 ) ;
  assign n376 = n371 | n375 ;
  assign n377 = ~n138 & n139 ;
  assign n378 = ( ~n132 & n136 ) | ( ~n132 & n377 ) | ( n136 & n377 ) ;
  assign n379 = n133 | n378 ;
  assign n380 = ~n129 & n130 ;
  assign n381 = ( n129 & n379 ) | ( n129 & ~n380 ) | ( n379 & ~n380 ) ;
  assign n382 = n154 & ~n155 ;
  assign n383 = ( n155 & n381 ) | ( n155 & ~n382 ) | ( n381 & ~n382 ) ;
  assign n384 = n151 & ~n152 ;
  assign n385 = ( n152 & n383 ) | ( n152 & ~n384 ) | ( n383 & ~n384 ) ;
  assign n386 = ~n150 & n385 ;
  assign n387 = n159 & ~n386 ;
  assign n388 = n163 & ~n169 ;
  assign n389 = ( n168 & ~n170 ) | ( n168 & n388 ) | ( ~n170 & n388 ) ;
  assign n390 = n171 | n389 ;
  assign n391 = ~n184 & n185 ;
  assign n392 = ( ~n178 & n182 ) | ( ~n178 & n391 ) | ( n182 & n391 ) ;
  assign n393 = n179 | n392 ;
  assign n394 = ~n175 & n176 ;
  assign n395 = ( n175 & n393 ) | ( n175 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = ~n161 & n395 ;
  assign n397 = n164 | n173 ;
  assign n398 = n160 & ~n397 ;
  assign n399 = ( n396 & ~n397 ) | ( n396 & n398 ) | ( ~n397 & n398 ) ;
  assign n400 = n390 | n399 ;
  assign n401 = n159 | n400 ;
  assign n402 = ( n376 & ~n387 ) | ( n376 & n401 ) | ( ~n387 & n401 ) ;
  assign n403 = ~n149 & n153 ;
  assign n404 = n146 | n403 ;
  assign n405 = ~n135 & n138 ;
  assign n406 = ( n131 & ~n158 ) | ( n131 & n405 ) | ( ~n158 & n405 ) ;
  assign n407 = n404 | n406 ;
  assign n408 = ~n246 & n249 ;
  assign n409 = ( ~n237 & n242 ) | ( ~n237 & n408 ) | ( n242 & n408 ) ;
  assign n410 = ( ~n230 & n236 ) | ( ~n230 & n409 ) | ( n236 & n409 ) ;
  assign n411 = ( ~n223 & n226 ) | ( ~n223 & n410 ) | ( n226 & n410 ) ;
  assign n412 = n407 | n411 ;
  assign n413 = ~n181 & n184 ;
  assign n414 = ( ~n166 & n177 ) | ( ~n166 & n413 ) | ( n177 & n413 ) ;
  assign n415 = ( n165 & ~n169 ) | ( n165 & n414 ) | ( ~n169 & n414 ) ;
  assign n416 = n172 | n415 ;
  assign n417 = n209 & ~n220 ;
  assign n418 = ( ~n201 & n216 ) | ( ~n201 & n417 ) | ( n216 & n417 ) ;
  assign n419 = n204 | n418 ;
  assign n420 = ~n194 & n197 ;
  assign n421 = ( n194 & n419 ) | ( n194 & ~n420 ) | ( n419 & ~n420 ) ;
  assign n422 = ~n190 & n421 ;
  assign n423 = n416 | n422 ;
  assign n424 = ~n159 & n423 ;
  assign n425 = n412 | n424 ;
  assign n426 = ~n238 & n246 ;
  assign n427 = ( ~n213 & n230 ) | ( ~n213 & n426 ) | ( n230 & n426 ) ;
  assign n428 = n220 | n427 ;
  assign n429 = ~n198 & n205 ;
  assign n430 = ( n198 & n428 ) | ( n198 & ~n429 ) | ( n428 & ~n429 ) ;
  assign n431 = ~n191 & n430 ;
  assign n432 = ~n174 & n181 ;
  assign n433 = ( ~n143 & n173 ) | ( ~n143 & n432 ) | ( n173 & n432 ) ;
  assign n434 = ( n135 & ~n157 ) | ( n135 & n433 ) | ( ~n157 & n433 ) ;
  assign n435 = n150 | n434 ;
  assign n436 = n431 | n435 ;
  assign n437 = ~n223 & n238 ;
  assign n438 = ~n190 & n206 ;
  assign n439 = ( ~n143 & n174 ) | ( ~n143 & n438 ) | ( n174 & n438 ) ;
  assign n440 = n158 | n439 ;
  assign n441 = n437 | n440 ;
  assign n442 = ( n159 & ~n190 ) | ( n159 & n223 ) | ( ~n190 & n223 ) ;
  assign y0 = n255 ;
  assign y1 = n349 ;
  assign y2 = n402 ;
  assign y3 = n425 ;
  assign y4 = n436 ;
  assign y5 = n441 ;
  assign y6 = n442 ;
  assign y7 = n191 ;
endmodule
