module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 ;
  assign n513 = x0 & ~x128 ;
  assign n514 = ( x1 & ~x129 ) | ( x1 & n513 ) | ( ~x129 & n513 ) ;
  assign n515 = ( x2 & ~x130 ) | ( x2 & n514 ) | ( ~x130 & n514 ) ;
  assign n516 = ( x3 & ~x131 ) | ( x3 & n515 ) | ( ~x131 & n515 ) ;
  assign n517 = ( x4 & ~x132 ) | ( x4 & n516 ) | ( ~x132 & n516 ) ;
  assign n518 = ( x5 & ~x133 ) | ( x5 & n517 ) | ( ~x133 & n517 ) ;
  assign n519 = ( x6 & ~x134 ) | ( x6 & n518 ) | ( ~x134 & n518 ) ;
  assign n520 = ( x7 & ~x135 ) | ( x7 & n519 ) | ( ~x135 & n519 ) ;
  assign n521 = ( x8 & ~x136 ) | ( x8 & n520 ) | ( ~x136 & n520 ) ;
  assign n522 = ( x9 & ~x137 ) | ( x9 & n521 ) | ( ~x137 & n521 ) ;
  assign n523 = ( x10 & ~x138 ) | ( x10 & n522 ) | ( ~x138 & n522 ) ;
  assign n524 = ( x11 & ~x139 ) | ( x11 & n523 ) | ( ~x139 & n523 ) ;
  assign n525 = ( x12 & ~x140 ) | ( x12 & n524 ) | ( ~x140 & n524 ) ;
  assign n526 = ( x13 & ~x141 ) | ( x13 & n525 ) | ( ~x141 & n525 ) ;
  assign n527 = ( x14 & ~x142 ) | ( x14 & n526 ) | ( ~x142 & n526 ) ;
  assign n528 = ( x15 & ~x143 ) | ( x15 & n527 ) | ( ~x143 & n527 ) ;
  assign n529 = ( x16 & ~x144 ) | ( x16 & n528 ) | ( ~x144 & n528 ) ;
  assign n530 = ( x17 & ~x145 ) | ( x17 & n529 ) | ( ~x145 & n529 ) ;
  assign n531 = ( x18 & ~x146 ) | ( x18 & n530 ) | ( ~x146 & n530 ) ;
  assign n532 = ( x19 & ~x147 ) | ( x19 & n531 ) | ( ~x147 & n531 ) ;
  assign n533 = ( x20 & ~x148 ) | ( x20 & n532 ) | ( ~x148 & n532 ) ;
  assign n534 = ( x21 & ~x149 ) | ( x21 & n533 ) | ( ~x149 & n533 ) ;
  assign n535 = ( x22 & ~x150 ) | ( x22 & n534 ) | ( ~x150 & n534 ) ;
  assign n536 = ( x23 & ~x151 ) | ( x23 & n535 ) | ( ~x151 & n535 ) ;
  assign n537 = ( x24 & ~x152 ) | ( x24 & n536 ) | ( ~x152 & n536 ) ;
  assign n538 = ( x25 & ~x153 ) | ( x25 & n537 ) | ( ~x153 & n537 ) ;
  assign n539 = ( x26 & ~x154 ) | ( x26 & n538 ) | ( ~x154 & n538 ) ;
  assign n540 = ( x27 & ~x155 ) | ( x27 & n539 ) | ( ~x155 & n539 ) ;
  assign n541 = ( x28 & ~x156 ) | ( x28 & n540 ) | ( ~x156 & n540 ) ;
  assign n542 = ( x29 & ~x157 ) | ( x29 & n541 ) | ( ~x157 & n541 ) ;
  assign n543 = ( x30 & ~x158 ) | ( x30 & n542 ) | ( ~x158 & n542 ) ;
  assign n544 = ( x31 & ~x159 ) | ( x31 & n543 ) | ( ~x159 & n543 ) ;
  assign n545 = ( x32 & ~x160 ) | ( x32 & n544 ) | ( ~x160 & n544 ) ;
  assign n546 = ( x33 & ~x161 ) | ( x33 & n545 ) | ( ~x161 & n545 ) ;
  assign n547 = ( x34 & ~x162 ) | ( x34 & n546 ) | ( ~x162 & n546 ) ;
  assign n548 = ( x35 & ~x163 ) | ( x35 & n547 ) | ( ~x163 & n547 ) ;
  assign n549 = ( x36 & ~x164 ) | ( x36 & n548 ) | ( ~x164 & n548 ) ;
  assign n550 = ( x37 & ~x165 ) | ( x37 & n549 ) | ( ~x165 & n549 ) ;
  assign n551 = ( x38 & ~x166 ) | ( x38 & n550 ) | ( ~x166 & n550 ) ;
  assign n552 = ( x39 & ~x167 ) | ( x39 & n551 ) | ( ~x167 & n551 ) ;
  assign n553 = ( x40 & ~x168 ) | ( x40 & n552 ) | ( ~x168 & n552 ) ;
  assign n554 = ( x41 & ~x169 ) | ( x41 & n553 ) | ( ~x169 & n553 ) ;
  assign n555 = ( x42 & ~x170 ) | ( x42 & n554 ) | ( ~x170 & n554 ) ;
  assign n556 = ( x43 & ~x171 ) | ( x43 & n555 ) | ( ~x171 & n555 ) ;
  assign n557 = ( x44 & ~x172 ) | ( x44 & n556 ) | ( ~x172 & n556 ) ;
  assign n558 = ( x45 & ~x173 ) | ( x45 & n557 ) | ( ~x173 & n557 ) ;
  assign n559 = ( x46 & ~x174 ) | ( x46 & n558 ) | ( ~x174 & n558 ) ;
  assign n560 = ( x47 & ~x175 ) | ( x47 & n559 ) | ( ~x175 & n559 ) ;
  assign n561 = ( x48 & ~x176 ) | ( x48 & n560 ) | ( ~x176 & n560 ) ;
  assign n562 = ( x49 & ~x177 ) | ( x49 & n561 ) | ( ~x177 & n561 ) ;
  assign n563 = ( x50 & ~x178 ) | ( x50 & n562 ) | ( ~x178 & n562 ) ;
  assign n564 = ( x51 & ~x179 ) | ( x51 & n563 ) | ( ~x179 & n563 ) ;
  assign n565 = ( x52 & ~x180 ) | ( x52 & n564 ) | ( ~x180 & n564 ) ;
  assign n566 = ( x53 & ~x181 ) | ( x53 & n565 ) | ( ~x181 & n565 ) ;
  assign n567 = ( x54 & ~x182 ) | ( x54 & n566 ) | ( ~x182 & n566 ) ;
  assign n568 = ( x55 & ~x183 ) | ( x55 & n567 ) | ( ~x183 & n567 ) ;
  assign n569 = ( x56 & ~x184 ) | ( x56 & n568 ) | ( ~x184 & n568 ) ;
  assign n570 = ( x57 & ~x185 ) | ( x57 & n569 ) | ( ~x185 & n569 ) ;
  assign n571 = ( x58 & ~x186 ) | ( x58 & n570 ) | ( ~x186 & n570 ) ;
  assign n572 = ( x59 & ~x187 ) | ( x59 & n571 ) | ( ~x187 & n571 ) ;
  assign n573 = ( x60 & ~x188 ) | ( x60 & n572 ) | ( ~x188 & n572 ) ;
  assign n574 = ( x61 & ~x189 ) | ( x61 & n573 ) | ( ~x189 & n573 ) ;
  assign n575 = ( x62 & ~x190 ) | ( x62 & n574 ) | ( ~x190 & n574 ) ;
  assign n576 = ( x63 & ~x191 ) | ( x63 & n575 ) | ( ~x191 & n575 ) ;
  assign n577 = ( x64 & ~x192 ) | ( x64 & n576 ) | ( ~x192 & n576 ) ;
  assign n578 = ( x65 & ~x193 ) | ( x65 & n577 ) | ( ~x193 & n577 ) ;
  assign n579 = ( x66 & ~x194 ) | ( x66 & n578 ) | ( ~x194 & n578 ) ;
  assign n580 = ( x67 & ~x195 ) | ( x67 & n579 ) | ( ~x195 & n579 ) ;
  assign n581 = ( x68 & ~x196 ) | ( x68 & n580 ) | ( ~x196 & n580 ) ;
  assign n582 = ( x69 & ~x197 ) | ( x69 & n581 ) | ( ~x197 & n581 ) ;
  assign n583 = ( x70 & ~x198 ) | ( x70 & n582 ) | ( ~x198 & n582 ) ;
  assign n584 = ( x71 & ~x199 ) | ( x71 & n583 ) | ( ~x199 & n583 ) ;
  assign n585 = ( x72 & ~x200 ) | ( x72 & n584 ) | ( ~x200 & n584 ) ;
  assign n586 = ( x73 & ~x201 ) | ( x73 & n585 ) | ( ~x201 & n585 ) ;
  assign n587 = ( x74 & ~x202 ) | ( x74 & n586 ) | ( ~x202 & n586 ) ;
  assign n588 = ( x75 & ~x203 ) | ( x75 & n587 ) | ( ~x203 & n587 ) ;
  assign n589 = ( x76 & ~x204 ) | ( x76 & n588 ) | ( ~x204 & n588 ) ;
  assign n590 = ( x77 & ~x205 ) | ( x77 & n589 ) | ( ~x205 & n589 ) ;
  assign n591 = ( x78 & ~x206 ) | ( x78 & n590 ) | ( ~x206 & n590 ) ;
  assign n592 = ( x79 & ~x207 ) | ( x79 & n591 ) | ( ~x207 & n591 ) ;
  assign n593 = ( x80 & ~x208 ) | ( x80 & n592 ) | ( ~x208 & n592 ) ;
  assign n594 = ( x81 & ~x209 ) | ( x81 & n593 ) | ( ~x209 & n593 ) ;
  assign n595 = ( x82 & ~x210 ) | ( x82 & n594 ) | ( ~x210 & n594 ) ;
  assign n596 = ( x83 & ~x211 ) | ( x83 & n595 ) | ( ~x211 & n595 ) ;
  assign n597 = ( x84 & ~x212 ) | ( x84 & n596 ) | ( ~x212 & n596 ) ;
  assign n598 = ( x85 & ~x213 ) | ( x85 & n597 ) | ( ~x213 & n597 ) ;
  assign n599 = ( x86 & ~x214 ) | ( x86 & n598 ) | ( ~x214 & n598 ) ;
  assign n600 = ( x87 & ~x215 ) | ( x87 & n599 ) | ( ~x215 & n599 ) ;
  assign n601 = ( x88 & ~x216 ) | ( x88 & n600 ) | ( ~x216 & n600 ) ;
  assign n602 = ( x89 & ~x217 ) | ( x89 & n601 ) | ( ~x217 & n601 ) ;
  assign n603 = ( x90 & ~x218 ) | ( x90 & n602 ) | ( ~x218 & n602 ) ;
  assign n604 = ( x91 & ~x219 ) | ( x91 & n603 ) | ( ~x219 & n603 ) ;
  assign n605 = ( x92 & ~x220 ) | ( x92 & n604 ) | ( ~x220 & n604 ) ;
  assign n606 = ( x93 & ~x221 ) | ( x93 & n605 ) | ( ~x221 & n605 ) ;
  assign n607 = ( x94 & ~x222 ) | ( x94 & n606 ) | ( ~x222 & n606 ) ;
  assign n608 = ( x95 & ~x223 ) | ( x95 & n607 ) | ( ~x223 & n607 ) ;
  assign n609 = ( x96 & ~x224 ) | ( x96 & n608 ) | ( ~x224 & n608 ) ;
  assign n610 = ( x97 & ~x225 ) | ( x97 & n609 ) | ( ~x225 & n609 ) ;
  assign n611 = ( x98 & ~x226 ) | ( x98 & n610 ) | ( ~x226 & n610 ) ;
  assign n612 = ( x99 & ~x227 ) | ( x99 & n611 ) | ( ~x227 & n611 ) ;
  assign n613 = ( x100 & ~x228 ) | ( x100 & n612 ) | ( ~x228 & n612 ) ;
  assign n614 = ( x101 & ~x229 ) | ( x101 & n613 ) | ( ~x229 & n613 ) ;
  assign n615 = ( x102 & ~x230 ) | ( x102 & n614 ) | ( ~x230 & n614 ) ;
  assign n616 = ( x103 & ~x231 ) | ( x103 & n615 ) | ( ~x231 & n615 ) ;
  assign n617 = ( x104 & ~x232 ) | ( x104 & n616 ) | ( ~x232 & n616 ) ;
  assign n618 = ( x105 & ~x233 ) | ( x105 & n617 ) | ( ~x233 & n617 ) ;
  assign n619 = ( x106 & ~x234 ) | ( x106 & n618 ) | ( ~x234 & n618 ) ;
  assign n620 = ( x107 & ~x235 ) | ( x107 & n619 ) | ( ~x235 & n619 ) ;
  assign n621 = ( x108 & ~x236 ) | ( x108 & n620 ) | ( ~x236 & n620 ) ;
  assign n622 = ( x109 & ~x237 ) | ( x109 & n621 ) | ( ~x237 & n621 ) ;
  assign n623 = ( x110 & ~x238 ) | ( x110 & n622 ) | ( ~x238 & n622 ) ;
  assign n624 = ( x111 & ~x239 ) | ( x111 & n623 ) | ( ~x239 & n623 ) ;
  assign n625 = ( x112 & ~x240 ) | ( x112 & n624 ) | ( ~x240 & n624 ) ;
  assign n626 = ( x113 & ~x241 ) | ( x113 & n625 ) | ( ~x241 & n625 ) ;
  assign n627 = ( x114 & ~x242 ) | ( x114 & n626 ) | ( ~x242 & n626 ) ;
  assign n628 = ( x115 & ~x243 ) | ( x115 & n627 ) | ( ~x243 & n627 ) ;
  assign n629 = ( x116 & ~x244 ) | ( x116 & n628 ) | ( ~x244 & n628 ) ;
  assign n630 = ( x117 & ~x245 ) | ( x117 & n629 ) | ( ~x245 & n629 ) ;
  assign n631 = ( x118 & ~x246 ) | ( x118 & n630 ) | ( ~x246 & n630 ) ;
  assign n632 = ( x119 & ~x247 ) | ( x119 & n631 ) | ( ~x247 & n631 ) ;
  assign n633 = ( x120 & ~x248 ) | ( x120 & n632 ) | ( ~x248 & n632 ) ;
  assign n634 = ( x121 & ~x249 ) | ( x121 & n633 ) | ( ~x249 & n633 ) ;
  assign n635 = ( x122 & ~x250 ) | ( x122 & n634 ) | ( ~x250 & n634 ) ;
  assign n636 = ( x123 & ~x251 ) | ( x123 & n635 ) | ( ~x251 & n635 ) ;
  assign n637 = ( x124 & ~x252 ) | ( x124 & n636 ) | ( ~x252 & n636 ) ;
  assign n638 = ( x125 & ~x253 ) | ( x125 & n637 ) | ( ~x253 & n637 ) ;
  assign n639 = ( x126 & ~x254 ) | ( x126 & n638 ) | ( ~x254 & n638 ) ;
  assign n640 = ( ~x127 & x255 ) | ( ~x127 & n639 ) | ( x255 & n639 ) ;
  assign n641 = x0 & n640 ;
  assign n642 = x128 & ~n640 ;
  assign n643 = n641 | n642 ;
  assign n644 = x256 & ~x384 ;
  assign n645 = ( x257 & ~x385 ) | ( x257 & n644 ) | ( ~x385 & n644 ) ;
  assign n646 = ( x258 & ~x386 ) | ( x258 & n645 ) | ( ~x386 & n645 ) ;
  assign n647 = ( x259 & ~x387 ) | ( x259 & n646 ) | ( ~x387 & n646 ) ;
  assign n648 = ( x260 & ~x388 ) | ( x260 & n647 ) | ( ~x388 & n647 ) ;
  assign n649 = ( x261 & ~x389 ) | ( x261 & n648 ) | ( ~x389 & n648 ) ;
  assign n650 = ( x262 & ~x390 ) | ( x262 & n649 ) | ( ~x390 & n649 ) ;
  assign n651 = ( x263 & ~x391 ) | ( x263 & n650 ) | ( ~x391 & n650 ) ;
  assign n652 = ( x264 & ~x392 ) | ( x264 & n651 ) | ( ~x392 & n651 ) ;
  assign n653 = ( x265 & ~x393 ) | ( x265 & n652 ) | ( ~x393 & n652 ) ;
  assign n654 = ( x266 & ~x394 ) | ( x266 & n653 ) | ( ~x394 & n653 ) ;
  assign n655 = ( x267 & ~x395 ) | ( x267 & n654 ) | ( ~x395 & n654 ) ;
  assign n656 = ( x268 & ~x396 ) | ( x268 & n655 ) | ( ~x396 & n655 ) ;
  assign n657 = ( x269 & ~x397 ) | ( x269 & n656 ) | ( ~x397 & n656 ) ;
  assign n658 = ( x270 & ~x398 ) | ( x270 & n657 ) | ( ~x398 & n657 ) ;
  assign n659 = ( x271 & ~x399 ) | ( x271 & n658 ) | ( ~x399 & n658 ) ;
  assign n660 = ( x272 & ~x400 ) | ( x272 & n659 ) | ( ~x400 & n659 ) ;
  assign n661 = ( x273 & ~x401 ) | ( x273 & n660 ) | ( ~x401 & n660 ) ;
  assign n662 = ( x274 & ~x402 ) | ( x274 & n661 ) | ( ~x402 & n661 ) ;
  assign n663 = ( x275 & ~x403 ) | ( x275 & n662 ) | ( ~x403 & n662 ) ;
  assign n664 = ( x276 & ~x404 ) | ( x276 & n663 ) | ( ~x404 & n663 ) ;
  assign n665 = ( x277 & ~x405 ) | ( x277 & n664 ) | ( ~x405 & n664 ) ;
  assign n666 = ( x278 & ~x406 ) | ( x278 & n665 ) | ( ~x406 & n665 ) ;
  assign n667 = ( x279 & ~x407 ) | ( x279 & n666 ) | ( ~x407 & n666 ) ;
  assign n668 = ( x280 & ~x408 ) | ( x280 & n667 ) | ( ~x408 & n667 ) ;
  assign n669 = ( x281 & ~x409 ) | ( x281 & n668 ) | ( ~x409 & n668 ) ;
  assign n670 = ( x282 & ~x410 ) | ( x282 & n669 ) | ( ~x410 & n669 ) ;
  assign n671 = ( x283 & ~x411 ) | ( x283 & n670 ) | ( ~x411 & n670 ) ;
  assign n672 = ( x284 & ~x412 ) | ( x284 & n671 ) | ( ~x412 & n671 ) ;
  assign n673 = ( x285 & ~x413 ) | ( x285 & n672 ) | ( ~x413 & n672 ) ;
  assign n674 = ( x286 & ~x414 ) | ( x286 & n673 ) | ( ~x414 & n673 ) ;
  assign n675 = ( x287 & ~x415 ) | ( x287 & n674 ) | ( ~x415 & n674 ) ;
  assign n676 = ( x288 & ~x416 ) | ( x288 & n675 ) | ( ~x416 & n675 ) ;
  assign n677 = ( x289 & ~x417 ) | ( x289 & n676 ) | ( ~x417 & n676 ) ;
  assign n678 = ( x290 & ~x418 ) | ( x290 & n677 ) | ( ~x418 & n677 ) ;
  assign n679 = ( x291 & ~x419 ) | ( x291 & n678 ) | ( ~x419 & n678 ) ;
  assign n680 = ( x292 & ~x420 ) | ( x292 & n679 ) | ( ~x420 & n679 ) ;
  assign n681 = ( x293 & ~x421 ) | ( x293 & n680 ) | ( ~x421 & n680 ) ;
  assign n682 = ( x294 & ~x422 ) | ( x294 & n681 ) | ( ~x422 & n681 ) ;
  assign n683 = ( x295 & ~x423 ) | ( x295 & n682 ) | ( ~x423 & n682 ) ;
  assign n684 = ( x296 & ~x424 ) | ( x296 & n683 ) | ( ~x424 & n683 ) ;
  assign n685 = ( x297 & ~x425 ) | ( x297 & n684 ) | ( ~x425 & n684 ) ;
  assign n686 = ( x298 & ~x426 ) | ( x298 & n685 ) | ( ~x426 & n685 ) ;
  assign n687 = ( x299 & ~x427 ) | ( x299 & n686 ) | ( ~x427 & n686 ) ;
  assign n688 = ( x300 & ~x428 ) | ( x300 & n687 ) | ( ~x428 & n687 ) ;
  assign n689 = ( x301 & ~x429 ) | ( x301 & n688 ) | ( ~x429 & n688 ) ;
  assign n690 = ( x302 & ~x430 ) | ( x302 & n689 ) | ( ~x430 & n689 ) ;
  assign n691 = ( x303 & ~x431 ) | ( x303 & n690 ) | ( ~x431 & n690 ) ;
  assign n692 = ( x304 & ~x432 ) | ( x304 & n691 ) | ( ~x432 & n691 ) ;
  assign n693 = ( x305 & ~x433 ) | ( x305 & n692 ) | ( ~x433 & n692 ) ;
  assign n694 = ( x306 & ~x434 ) | ( x306 & n693 ) | ( ~x434 & n693 ) ;
  assign n695 = ( x307 & ~x435 ) | ( x307 & n694 ) | ( ~x435 & n694 ) ;
  assign n696 = ( x308 & ~x436 ) | ( x308 & n695 ) | ( ~x436 & n695 ) ;
  assign n697 = ( x309 & ~x437 ) | ( x309 & n696 ) | ( ~x437 & n696 ) ;
  assign n698 = ( x310 & ~x438 ) | ( x310 & n697 ) | ( ~x438 & n697 ) ;
  assign n699 = ( x311 & ~x439 ) | ( x311 & n698 ) | ( ~x439 & n698 ) ;
  assign n700 = ( x312 & ~x440 ) | ( x312 & n699 ) | ( ~x440 & n699 ) ;
  assign n701 = ( x313 & ~x441 ) | ( x313 & n700 ) | ( ~x441 & n700 ) ;
  assign n702 = ( x314 & ~x442 ) | ( x314 & n701 ) | ( ~x442 & n701 ) ;
  assign n703 = ( x315 & ~x443 ) | ( x315 & n702 ) | ( ~x443 & n702 ) ;
  assign n704 = ( x316 & ~x444 ) | ( x316 & n703 ) | ( ~x444 & n703 ) ;
  assign n705 = ( x317 & ~x445 ) | ( x317 & n704 ) | ( ~x445 & n704 ) ;
  assign n706 = ( x318 & ~x446 ) | ( x318 & n705 ) | ( ~x446 & n705 ) ;
  assign n707 = ( x319 & ~x447 ) | ( x319 & n706 ) | ( ~x447 & n706 ) ;
  assign n708 = ( x320 & ~x448 ) | ( x320 & n707 ) | ( ~x448 & n707 ) ;
  assign n709 = ( x321 & ~x449 ) | ( x321 & n708 ) | ( ~x449 & n708 ) ;
  assign n710 = ( x322 & ~x450 ) | ( x322 & n709 ) | ( ~x450 & n709 ) ;
  assign n711 = ( x323 & ~x451 ) | ( x323 & n710 ) | ( ~x451 & n710 ) ;
  assign n712 = ( x324 & ~x452 ) | ( x324 & n711 ) | ( ~x452 & n711 ) ;
  assign n713 = ( x325 & ~x453 ) | ( x325 & n712 ) | ( ~x453 & n712 ) ;
  assign n714 = ( x326 & ~x454 ) | ( x326 & n713 ) | ( ~x454 & n713 ) ;
  assign n715 = ( x327 & ~x455 ) | ( x327 & n714 ) | ( ~x455 & n714 ) ;
  assign n716 = ( x328 & ~x456 ) | ( x328 & n715 ) | ( ~x456 & n715 ) ;
  assign n717 = ( x329 & ~x457 ) | ( x329 & n716 ) | ( ~x457 & n716 ) ;
  assign n718 = ( x330 & ~x458 ) | ( x330 & n717 ) | ( ~x458 & n717 ) ;
  assign n719 = ( x331 & ~x459 ) | ( x331 & n718 ) | ( ~x459 & n718 ) ;
  assign n720 = ( x332 & ~x460 ) | ( x332 & n719 ) | ( ~x460 & n719 ) ;
  assign n721 = ( x333 & ~x461 ) | ( x333 & n720 ) | ( ~x461 & n720 ) ;
  assign n722 = ( x334 & ~x462 ) | ( x334 & n721 ) | ( ~x462 & n721 ) ;
  assign n723 = ( x335 & ~x463 ) | ( x335 & n722 ) | ( ~x463 & n722 ) ;
  assign n724 = ( x336 & ~x464 ) | ( x336 & n723 ) | ( ~x464 & n723 ) ;
  assign n725 = ( x337 & ~x465 ) | ( x337 & n724 ) | ( ~x465 & n724 ) ;
  assign n726 = ( x338 & ~x466 ) | ( x338 & n725 ) | ( ~x466 & n725 ) ;
  assign n727 = ( x339 & ~x467 ) | ( x339 & n726 ) | ( ~x467 & n726 ) ;
  assign n728 = ( x340 & ~x468 ) | ( x340 & n727 ) | ( ~x468 & n727 ) ;
  assign n729 = ( x341 & ~x469 ) | ( x341 & n728 ) | ( ~x469 & n728 ) ;
  assign n730 = ( x342 & ~x470 ) | ( x342 & n729 ) | ( ~x470 & n729 ) ;
  assign n731 = ( x343 & ~x471 ) | ( x343 & n730 ) | ( ~x471 & n730 ) ;
  assign n732 = ( x344 & ~x472 ) | ( x344 & n731 ) | ( ~x472 & n731 ) ;
  assign n733 = ( x345 & ~x473 ) | ( x345 & n732 ) | ( ~x473 & n732 ) ;
  assign n734 = ( x346 & ~x474 ) | ( x346 & n733 ) | ( ~x474 & n733 ) ;
  assign n735 = ( x347 & ~x475 ) | ( x347 & n734 ) | ( ~x475 & n734 ) ;
  assign n736 = ( x348 & ~x476 ) | ( x348 & n735 ) | ( ~x476 & n735 ) ;
  assign n737 = ( x349 & ~x477 ) | ( x349 & n736 ) | ( ~x477 & n736 ) ;
  assign n738 = ( x350 & ~x478 ) | ( x350 & n737 ) | ( ~x478 & n737 ) ;
  assign n739 = ( x351 & ~x479 ) | ( x351 & n738 ) | ( ~x479 & n738 ) ;
  assign n740 = ( x352 & ~x480 ) | ( x352 & n739 ) | ( ~x480 & n739 ) ;
  assign n741 = ( x353 & ~x481 ) | ( x353 & n740 ) | ( ~x481 & n740 ) ;
  assign n742 = ( x354 & ~x482 ) | ( x354 & n741 ) | ( ~x482 & n741 ) ;
  assign n743 = ( x355 & ~x483 ) | ( x355 & n742 ) | ( ~x483 & n742 ) ;
  assign n744 = ( x356 & ~x484 ) | ( x356 & n743 ) | ( ~x484 & n743 ) ;
  assign n745 = ( x357 & ~x485 ) | ( x357 & n744 ) | ( ~x485 & n744 ) ;
  assign n746 = ( x358 & ~x486 ) | ( x358 & n745 ) | ( ~x486 & n745 ) ;
  assign n747 = ( x359 & ~x487 ) | ( x359 & n746 ) | ( ~x487 & n746 ) ;
  assign n748 = ( x360 & ~x488 ) | ( x360 & n747 ) | ( ~x488 & n747 ) ;
  assign n749 = ( x361 & ~x489 ) | ( x361 & n748 ) | ( ~x489 & n748 ) ;
  assign n750 = ( x362 & ~x490 ) | ( x362 & n749 ) | ( ~x490 & n749 ) ;
  assign n751 = ( x363 & ~x491 ) | ( x363 & n750 ) | ( ~x491 & n750 ) ;
  assign n752 = ( x364 & ~x492 ) | ( x364 & n751 ) | ( ~x492 & n751 ) ;
  assign n753 = ( x365 & ~x493 ) | ( x365 & n752 ) | ( ~x493 & n752 ) ;
  assign n754 = ( x366 & ~x494 ) | ( x366 & n753 ) | ( ~x494 & n753 ) ;
  assign n755 = ( x367 & ~x495 ) | ( x367 & n754 ) | ( ~x495 & n754 ) ;
  assign n756 = ( x368 & ~x496 ) | ( x368 & n755 ) | ( ~x496 & n755 ) ;
  assign n757 = ( x369 & ~x497 ) | ( x369 & n756 ) | ( ~x497 & n756 ) ;
  assign n758 = ( x370 & ~x498 ) | ( x370 & n757 ) | ( ~x498 & n757 ) ;
  assign n759 = ( x371 & ~x499 ) | ( x371 & n758 ) | ( ~x499 & n758 ) ;
  assign n760 = ( x372 & ~x500 ) | ( x372 & n759 ) | ( ~x500 & n759 ) ;
  assign n761 = ( x373 & ~x501 ) | ( x373 & n760 ) | ( ~x501 & n760 ) ;
  assign n762 = ( x374 & ~x502 ) | ( x374 & n761 ) | ( ~x502 & n761 ) ;
  assign n763 = ( x375 & ~x503 ) | ( x375 & n762 ) | ( ~x503 & n762 ) ;
  assign n764 = ( x376 & ~x504 ) | ( x376 & n763 ) | ( ~x504 & n763 ) ;
  assign n765 = ( x377 & ~x505 ) | ( x377 & n764 ) | ( ~x505 & n764 ) ;
  assign n766 = ( x378 & ~x506 ) | ( x378 & n765 ) | ( ~x506 & n765 ) ;
  assign n767 = ( x379 & ~x507 ) | ( x379 & n766 ) | ( ~x507 & n766 ) ;
  assign n768 = ( x380 & ~x508 ) | ( x380 & n767 ) | ( ~x508 & n767 ) ;
  assign n769 = ( x381 & ~x509 ) | ( x381 & n768 ) | ( ~x509 & n768 ) ;
  assign n770 = ( x382 & ~x510 ) | ( x382 & n769 ) | ( ~x510 & n769 ) ;
  assign n771 = ( ~x383 & x511 ) | ( ~x383 & n770 ) | ( x511 & n770 ) ;
  assign n772 = x375 & n771 ;
  assign n773 = x503 & ~n771 ;
  assign n774 = n772 | n773 ;
  assign n775 = x119 & n640 ;
  assign n776 = x247 & ~n640 ;
  assign n777 = n775 | n776 ;
  assign n778 = x368 & n771 ;
  assign n779 = x496 & ~n771 ;
  assign n780 = n778 | n779 ;
  assign n781 = x112 & n640 ;
  assign n782 = x240 & ~n640 ;
  assign n783 = n781 | n782 ;
  assign n784 = x349 & n771 ;
  assign n785 = x477 & ~n771 ;
  assign n786 = n784 | n785 ;
  assign n787 = x93 & n640 ;
  assign n788 = x221 & ~n640 ;
  assign n789 = n787 | n788 ;
  assign n790 = x345 & n771 ;
  assign n791 = x473 & ~n771 ;
  assign n792 = n790 | n791 ;
  assign n793 = x89 & n640 ;
  assign n794 = x217 & ~n640 ;
  assign n795 = n793 | n794 ;
  assign n796 = x330 & n771 ;
  assign n797 = x458 & ~n771 ;
  assign n798 = n796 | n797 ;
  assign n799 = x74 & n640 ;
  assign n800 = x202 & ~n640 ;
  assign n801 = n799 | n800 ;
  assign n802 = x260 & n771 ;
  assign n803 = x388 & ~n771 ;
  assign n804 = n802 | n803 ;
  assign n805 = x4 & n640 ;
  assign n806 = x132 & ~n640 ;
  assign n807 = n805 | n806 ;
  assign n808 = x1 & n640 ;
  assign n809 = x129 & ~n640 ;
  assign n810 = n808 | n809 ;
  assign n811 = x257 & n771 ;
  assign n812 = x385 & ~n771 ;
  assign n813 = n811 | n812 ;
  assign n814 = x256 & n771 ;
  assign n815 = x384 & ~n771 ;
  assign n816 = n814 | n815 ;
  assign n817 = n643 & ~n816 ;
  assign n818 = ( n810 & ~n813 ) | ( n810 & n817 ) | ( ~n813 & n817 ) ;
  assign n819 = x258 & n771 ;
  assign n820 = x386 & ~n771 ;
  assign n821 = n819 | n820 ;
  assign n822 = x2 & n640 ;
  assign n823 = x130 & ~n640 ;
  assign n824 = n822 | n823 ;
  assign n825 = ( n818 & ~n821 ) | ( n818 & n824 ) | ( ~n821 & n824 ) ;
  assign n826 = x3 & n640 ;
  assign n827 = x131 & ~n640 ;
  assign n828 = n826 | n827 ;
  assign n829 = x259 & n771 ;
  assign n830 = x387 & ~n771 ;
  assign n831 = n829 | n830 ;
  assign n832 = ( n825 & n828 ) | ( n825 & ~n831 ) | ( n828 & ~n831 ) ;
  assign n833 = ( ~n804 & n807 ) | ( ~n804 & n832 ) | ( n807 & n832 ) ;
  assign n834 = x5 & n640 ;
  assign n835 = x133 & ~n640 ;
  assign n836 = n834 | n835 ;
  assign n837 = x261 & n771 ;
  assign n838 = x389 & ~n771 ;
  assign n839 = n837 | n838 ;
  assign n840 = ( n833 & n836 ) | ( n833 & ~n839 ) | ( n836 & ~n839 ) ;
  assign n841 = x6 & n640 ;
  assign n842 = x134 & ~n640 ;
  assign n843 = n841 | n842 ;
  assign n844 = x262 & n771 ;
  assign n845 = x390 & ~n771 ;
  assign n846 = n844 | n845 ;
  assign n847 = ( n840 & n843 ) | ( n840 & ~n846 ) | ( n843 & ~n846 ) ;
  assign n848 = x263 & n771 ;
  assign n849 = x391 & ~n771 ;
  assign n850 = n848 | n849 ;
  assign n851 = x7 & n640 ;
  assign n852 = x135 & ~n640 ;
  assign n853 = n851 | n852 ;
  assign n854 = ( n847 & ~n850 ) | ( n847 & n853 ) | ( ~n850 & n853 ) ;
  assign n855 = x264 & n771 ;
  assign n856 = x392 & ~n771 ;
  assign n857 = n855 | n856 ;
  assign n858 = x8 & n640 ;
  assign n859 = x136 & ~n640 ;
  assign n860 = n858 | n859 ;
  assign n861 = ( n854 & ~n857 ) | ( n854 & n860 ) | ( ~n857 & n860 ) ;
  assign n862 = x9 & n640 ;
  assign n863 = x137 & ~n640 ;
  assign n864 = n862 | n863 ;
  assign n865 = x265 & n771 ;
  assign n866 = x393 & ~n771 ;
  assign n867 = n865 | n866 ;
  assign n868 = ( n861 & n864 ) | ( n861 & ~n867 ) | ( n864 & ~n867 ) ;
  assign n869 = x10 & n640 ;
  assign n870 = x138 & ~n640 ;
  assign n871 = n869 | n870 ;
  assign n872 = x266 & n771 ;
  assign n873 = x394 & ~n771 ;
  assign n874 = n872 | n873 ;
  assign n875 = ( n868 & n871 ) | ( n868 & ~n874 ) | ( n871 & ~n874 ) ;
  assign n876 = x267 & n771 ;
  assign n877 = x395 & ~n771 ;
  assign n878 = n876 | n877 ;
  assign n879 = x11 & n640 ;
  assign n880 = x139 & ~n640 ;
  assign n881 = n879 | n880 ;
  assign n882 = ( n875 & ~n878 ) | ( n875 & n881 ) | ( ~n878 & n881 ) ;
  assign n883 = x12 & n640 ;
  assign n884 = x140 & ~n640 ;
  assign n885 = n883 | n884 ;
  assign n886 = x268 & n771 ;
  assign n887 = x396 & ~n771 ;
  assign n888 = n886 | n887 ;
  assign n889 = ( n882 & n885 ) | ( n882 & ~n888 ) | ( n885 & ~n888 ) ;
  assign n890 = x269 & n771 ;
  assign n891 = x397 & ~n771 ;
  assign n892 = n890 | n891 ;
  assign n893 = x13 & n640 ;
  assign n894 = x141 & ~n640 ;
  assign n895 = n893 | n894 ;
  assign n896 = ( n889 & ~n892 ) | ( n889 & n895 ) | ( ~n892 & n895 ) ;
  assign n897 = x270 & n771 ;
  assign n898 = x398 & ~n771 ;
  assign n899 = n897 | n898 ;
  assign n900 = x14 & n640 ;
  assign n901 = x142 & ~n640 ;
  assign n902 = n900 | n901 ;
  assign n903 = ( n896 & ~n899 ) | ( n896 & n902 ) | ( ~n899 & n902 ) ;
  assign n904 = x15 & n640 ;
  assign n905 = x143 & ~n640 ;
  assign n906 = n904 | n905 ;
  assign n907 = x271 & n771 ;
  assign n908 = x399 & ~n771 ;
  assign n909 = n907 | n908 ;
  assign n910 = ( n903 & n906 ) | ( n903 & ~n909 ) | ( n906 & ~n909 ) ;
  assign n911 = x272 & n771 ;
  assign n912 = x400 & ~n771 ;
  assign n913 = n911 | n912 ;
  assign n914 = x16 & n640 ;
  assign n915 = x144 & ~n640 ;
  assign n916 = n914 | n915 ;
  assign n917 = ( n910 & ~n913 ) | ( n910 & n916 ) | ( ~n913 & n916 ) ;
  assign n918 = x273 & n771 ;
  assign n919 = x401 & ~n771 ;
  assign n920 = n918 | n919 ;
  assign n921 = x17 & n640 ;
  assign n922 = x145 & ~n640 ;
  assign n923 = n921 | n922 ;
  assign n924 = ( n917 & ~n920 ) | ( n917 & n923 ) | ( ~n920 & n923 ) ;
  assign n925 = x18 & n640 ;
  assign n926 = x146 & ~n640 ;
  assign n927 = n925 | n926 ;
  assign n928 = x274 & n771 ;
  assign n929 = x402 & ~n771 ;
  assign n930 = n928 | n929 ;
  assign n931 = ( n924 & n927 ) | ( n924 & ~n930 ) | ( n927 & ~n930 ) ;
  assign n932 = x19 & n640 ;
  assign n933 = x147 & ~n640 ;
  assign n934 = n932 | n933 ;
  assign n935 = x275 & n771 ;
  assign n936 = x403 & ~n771 ;
  assign n937 = n935 | n936 ;
  assign n938 = ( n931 & n934 ) | ( n931 & ~n937 ) | ( n934 & ~n937 ) ;
  assign n939 = x276 & n771 ;
  assign n940 = x404 & ~n771 ;
  assign n941 = n939 | n940 ;
  assign n942 = x20 & n640 ;
  assign n943 = x148 & ~n640 ;
  assign n944 = n942 | n943 ;
  assign n945 = ( n938 & ~n941 ) | ( n938 & n944 ) | ( ~n941 & n944 ) ;
  assign n946 = x21 & n640 ;
  assign n947 = x149 & ~n640 ;
  assign n948 = n946 | n947 ;
  assign n949 = x277 & n771 ;
  assign n950 = x405 & ~n771 ;
  assign n951 = n949 | n950 ;
  assign n952 = ( n945 & n948 ) | ( n945 & ~n951 ) | ( n948 & ~n951 ) ;
  assign n953 = x278 & n771 ;
  assign n954 = x406 & ~n771 ;
  assign n955 = n953 | n954 ;
  assign n956 = x22 & n640 ;
  assign n957 = x150 & ~n640 ;
  assign n958 = n956 | n957 ;
  assign n959 = ( n952 & ~n955 ) | ( n952 & n958 ) | ( ~n955 & n958 ) ;
  assign n960 = x279 & n771 ;
  assign n961 = x407 & ~n771 ;
  assign n962 = n960 | n961 ;
  assign n963 = x23 & n640 ;
  assign n964 = x151 & ~n640 ;
  assign n965 = n963 | n964 ;
  assign n966 = ( n959 & ~n962 ) | ( n959 & n965 ) | ( ~n962 & n965 ) ;
  assign n967 = x280 & n771 ;
  assign n968 = x408 & ~n771 ;
  assign n969 = n967 | n968 ;
  assign n970 = x24 & n640 ;
  assign n971 = x152 & ~n640 ;
  assign n972 = n970 | n971 ;
  assign n973 = ( n966 & ~n969 ) | ( n966 & n972 ) | ( ~n969 & n972 ) ;
  assign n974 = x281 & n771 ;
  assign n975 = x409 & ~n771 ;
  assign n976 = n974 | n975 ;
  assign n977 = x25 & n640 ;
  assign n978 = x153 & ~n640 ;
  assign n979 = n977 | n978 ;
  assign n980 = ( n973 & ~n976 ) | ( n973 & n979 ) | ( ~n976 & n979 ) ;
  assign n981 = x26 & n640 ;
  assign n982 = x154 & ~n640 ;
  assign n983 = n981 | n982 ;
  assign n984 = x282 & n771 ;
  assign n985 = x410 & ~n771 ;
  assign n986 = n984 | n985 ;
  assign n987 = ( n980 & n983 ) | ( n980 & ~n986 ) | ( n983 & ~n986 ) ;
  assign n988 = x283 & n771 ;
  assign n989 = x411 & ~n771 ;
  assign n990 = n988 | n989 ;
  assign n991 = x27 & n640 ;
  assign n992 = x155 & ~n640 ;
  assign n993 = n991 | n992 ;
  assign n994 = ( n987 & ~n990 ) | ( n987 & n993 ) | ( ~n990 & n993 ) ;
  assign n995 = x284 & n771 ;
  assign n996 = x412 & ~n771 ;
  assign n997 = n995 | n996 ;
  assign n998 = x28 & n640 ;
  assign n999 = x156 & ~n640 ;
  assign n1000 = n998 | n999 ;
  assign n1001 = ( n994 & ~n997 ) | ( n994 & n1000 ) | ( ~n997 & n1000 ) ;
  assign n1002 = x29 & n640 ;
  assign n1003 = x157 & ~n640 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = x285 & n771 ;
  assign n1006 = x413 & ~n771 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = ( n1001 & n1004 ) | ( n1001 & ~n1007 ) | ( n1004 & ~n1007 ) ;
  assign n1009 = x30 & n640 ;
  assign n1010 = x158 & ~n640 ;
  assign n1011 = n1009 | n1010 ;
  assign n1012 = x286 & n771 ;
  assign n1013 = x414 & ~n771 ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = ( n1008 & n1011 ) | ( n1008 & ~n1014 ) | ( n1011 & ~n1014 ) ;
  assign n1016 = x287 & n771 ;
  assign n1017 = x415 & ~n771 ;
  assign n1018 = n1016 | n1017 ;
  assign n1019 = x31 & n640 ;
  assign n1020 = x159 & ~n640 ;
  assign n1021 = n1019 | n1020 ;
  assign n1022 = ( n1015 & ~n1018 ) | ( n1015 & n1021 ) | ( ~n1018 & n1021 ) ;
  assign n1023 = x288 & n771 ;
  assign n1024 = x416 & ~n771 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = x32 & n640 ;
  assign n1027 = x160 & ~n640 ;
  assign n1028 = n1026 | n1027 ;
  assign n1029 = ( n1022 & ~n1025 ) | ( n1022 & n1028 ) | ( ~n1025 & n1028 ) ;
  assign n1030 = x33 & n640 ;
  assign n1031 = x161 & ~n640 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = x289 & n771 ;
  assign n1034 = x417 & ~n771 ;
  assign n1035 = n1033 | n1034 ;
  assign n1036 = ( n1029 & n1032 ) | ( n1029 & ~n1035 ) | ( n1032 & ~n1035 ) ;
  assign n1037 = x290 & n771 ;
  assign n1038 = x418 & ~n771 ;
  assign n1039 = n1037 | n1038 ;
  assign n1040 = x34 & n640 ;
  assign n1041 = x162 & ~n640 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = ( n1036 & ~n1039 ) | ( n1036 & n1042 ) | ( ~n1039 & n1042 ) ;
  assign n1044 = x35 & n640 ;
  assign n1045 = x163 & ~n640 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = x291 & n771 ;
  assign n1048 = x419 & ~n771 ;
  assign n1049 = n1047 | n1048 ;
  assign n1050 = ( n1043 & n1046 ) | ( n1043 & ~n1049 ) | ( n1046 & ~n1049 ) ;
  assign n1051 = x292 & n771 ;
  assign n1052 = x420 & ~n771 ;
  assign n1053 = n1051 | n1052 ;
  assign n1054 = x36 & n640 ;
  assign n1055 = x164 & ~n640 ;
  assign n1056 = n1054 | n1055 ;
  assign n1057 = ( n1050 & ~n1053 ) | ( n1050 & n1056 ) | ( ~n1053 & n1056 ) ;
  assign n1058 = x293 & n771 ;
  assign n1059 = x421 & ~n771 ;
  assign n1060 = n1058 | n1059 ;
  assign n1061 = x37 & n640 ;
  assign n1062 = x165 & ~n640 ;
  assign n1063 = n1061 | n1062 ;
  assign n1064 = ( n1057 & ~n1060 ) | ( n1057 & n1063 ) | ( ~n1060 & n1063 ) ;
  assign n1065 = x294 & n771 ;
  assign n1066 = x422 & ~n771 ;
  assign n1067 = n1065 | n1066 ;
  assign n1068 = x38 & n640 ;
  assign n1069 = x166 & ~n640 ;
  assign n1070 = n1068 | n1069 ;
  assign n1071 = ( n1064 & ~n1067 ) | ( n1064 & n1070 ) | ( ~n1067 & n1070 ) ;
  assign n1072 = x39 & n640 ;
  assign n1073 = x167 & ~n640 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = x295 & n771 ;
  assign n1076 = x423 & ~n771 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = ( n1071 & n1074 ) | ( n1071 & ~n1077 ) | ( n1074 & ~n1077 ) ;
  assign n1079 = x296 & n771 ;
  assign n1080 = x424 & ~n771 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = x40 & n640 ;
  assign n1083 = x168 & ~n640 ;
  assign n1084 = n1082 | n1083 ;
  assign n1085 = ( n1078 & ~n1081 ) | ( n1078 & n1084 ) | ( ~n1081 & n1084 ) ;
  assign n1086 = x297 & n771 ;
  assign n1087 = x425 & ~n771 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = x41 & n640 ;
  assign n1090 = x169 & ~n640 ;
  assign n1091 = n1089 | n1090 ;
  assign n1092 = ( n1085 & ~n1088 ) | ( n1085 & n1091 ) | ( ~n1088 & n1091 ) ;
  assign n1093 = x42 & n640 ;
  assign n1094 = x170 & ~n640 ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = x298 & n771 ;
  assign n1097 = x426 & ~n771 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = ( n1092 & n1095 ) | ( n1092 & ~n1098 ) | ( n1095 & ~n1098 ) ;
  assign n1100 = x43 & n640 ;
  assign n1101 = x171 & ~n640 ;
  assign n1102 = n1100 | n1101 ;
  assign n1103 = x299 & n771 ;
  assign n1104 = x427 & ~n771 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = ( n1099 & n1102 ) | ( n1099 & ~n1105 ) | ( n1102 & ~n1105 ) ;
  assign n1107 = x44 & n640 ;
  assign n1108 = x172 & ~n640 ;
  assign n1109 = n1107 | n1108 ;
  assign n1110 = x300 & n771 ;
  assign n1111 = x428 & ~n771 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = ( n1106 & n1109 ) | ( n1106 & ~n1112 ) | ( n1109 & ~n1112 ) ;
  assign n1114 = x301 & n771 ;
  assign n1115 = x429 & ~n771 ;
  assign n1116 = n1114 | n1115 ;
  assign n1117 = x45 & n640 ;
  assign n1118 = x173 & ~n640 ;
  assign n1119 = n1117 | n1118 ;
  assign n1120 = ( n1113 & ~n1116 ) | ( n1113 & n1119 ) | ( ~n1116 & n1119 ) ;
  assign n1121 = x302 & n771 ;
  assign n1122 = x430 & ~n771 ;
  assign n1123 = n1121 | n1122 ;
  assign n1124 = x46 & n640 ;
  assign n1125 = x174 & ~n640 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = ( n1120 & ~n1123 ) | ( n1120 & n1126 ) | ( ~n1123 & n1126 ) ;
  assign n1128 = x47 & n640 ;
  assign n1129 = x175 & ~n640 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = x303 & n771 ;
  assign n1132 = x431 & ~n771 ;
  assign n1133 = n1131 | n1132 ;
  assign n1134 = ( n1127 & n1130 ) | ( n1127 & ~n1133 ) | ( n1130 & ~n1133 ) ;
  assign n1135 = x304 & n771 ;
  assign n1136 = x432 & ~n771 ;
  assign n1137 = n1135 | n1136 ;
  assign n1138 = x48 & n640 ;
  assign n1139 = x176 & ~n640 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = ( n1134 & ~n1137 ) | ( n1134 & n1140 ) | ( ~n1137 & n1140 ) ;
  assign n1142 = x305 & n771 ;
  assign n1143 = x433 & ~n771 ;
  assign n1144 = n1142 | n1143 ;
  assign n1145 = x49 & n640 ;
  assign n1146 = x177 & ~n640 ;
  assign n1147 = n1145 | n1146 ;
  assign n1148 = ( n1141 & ~n1144 ) | ( n1141 & n1147 ) | ( ~n1144 & n1147 ) ;
  assign n1149 = x50 & n640 ;
  assign n1150 = x178 & ~n640 ;
  assign n1151 = n1149 | n1150 ;
  assign n1152 = x306 & n771 ;
  assign n1153 = x434 & ~n771 ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = ( n1148 & n1151 ) | ( n1148 & ~n1154 ) | ( n1151 & ~n1154 ) ;
  assign n1156 = x307 & n771 ;
  assign n1157 = x435 & ~n771 ;
  assign n1158 = n1156 | n1157 ;
  assign n1159 = x51 & n640 ;
  assign n1160 = x179 & ~n640 ;
  assign n1161 = n1159 | n1160 ;
  assign n1162 = ( n1155 & ~n1158 ) | ( n1155 & n1161 ) | ( ~n1158 & n1161 ) ;
  assign n1163 = x308 & n771 ;
  assign n1164 = x436 & ~n771 ;
  assign n1165 = n1163 | n1164 ;
  assign n1166 = x52 & n640 ;
  assign n1167 = x180 & ~n640 ;
  assign n1168 = n1166 | n1167 ;
  assign n1169 = ( n1162 & ~n1165 ) | ( n1162 & n1168 ) | ( ~n1165 & n1168 ) ;
  assign n1170 = x53 & n640 ;
  assign n1171 = x181 & ~n640 ;
  assign n1172 = n1170 | n1171 ;
  assign n1173 = x309 & n771 ;
  assign n1174 = x437 & ~n771 ;
  assign n1175 = n1173 | n1174 ;
  assign n1176 = ( n1169 & n1172 ) | ( n1169 & ~n1175 ) | ( n1172 & ~n1175 ) ;
  assign n1177 = x310 & n771 ;
  assign n1178 = x438 & ~n771 ;
  assign n1179 = n1177 | n1178 ;
  assign n1180 = x54 & n640 ;
  assign n1181 = x182 & ~n640 ;
  assign n1182 = n1180 | n1181 ;
  assign n1183 = ( n1176 & ~n1179 ) | ( n1176 & n1182 ) | ( ~n1179 & n1182 ) ;
  assign n1184 = x311 & n771 ;
  assign n1185 = x439 & ~n771 ;
  assign n1186 = n1184 | n1185 ;
  assign n1187 = x55 & n640 ;
  assign n1188 = x183 & ~n640 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = ( n1183 & ~n1186 ) | ( n1183 & n1189 ) | ( ~n1186 & n1189 ) ;
  assign n1191 = x56 & n640 ;
  assign n1192 = x184 & ~n640 ;
  assign n1193 = n1191 | n1192 ;
  assign n1194 = x312 & n771 ;
  assign n1195 = x440 & ~n771 ;
  assign n1196 = n1194 | n1195 ;
  assign n1197 = ( n1190 & n1193 ) | ( n1190 & ~n1196 ) | ( n1193 & ~n1196 ) ;
  assign n1198 = x57 & n640 ;
  assign n1199 = x185 & ~n640 ;
  assign n1200 = n1198 | n1199 ;
  assign n1201 = x313 & n771 ;
  assign n1202 = x441 & ~n771 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = ( n1197 & n1200 ) | ( n1197 & ~n1203 ) | ( n1200 & ~n1203 ) ;
  assign n1205 = x58 & n640 ;
  assign n1206 = x186 & ~n640 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = x314 & n771 ;
  assign n1209 = x442 & ~n771 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = ( n1204 & n1207 ) | ( n1204 & ~n1210 ) | ( n1207 & ~n1210 ) ;
  assign n1212 = x315 & n771 ;
  assign n1213 = x443 & ~n771 ;
  assign n1214 = n1212 | n1213 ;
  assign n1215 = x59 & n640 ;
  assign n1216 = x187 & ~n640 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = ( n1211 & ~n1214 ) | ( n1211 & n1217 ) | ( ~n1214 & n1217 ) ;
  assign n1219 = x60 & n640 ;
  assign n1220 = x188 & ~n640 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = x316 & n771 ;
  assign n1223 = x444 & ~n771 ;
  assign n1224 = n1222 | n1223 ;
  assign n1225 = ( n1218 & n1221 ) | ( n1218 & ~n1224 ) | ( n1221 & ~n1224 ) ;
  assign n1226 = x317 & n771 ;
  assign n1227 = x445 & ~n771 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = x61 & n640 ;
  assign n1230 = x189 & ~n640 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = ( n1225 & ~n1228 ) | ( n1225 & n1231 ) | ( ~n1228 & n1231 ) ;
  assign n1233 = x62 & n640 ;
  assign n1234 = x190 & ~n640 ;
  assign n1235 = n1233 | n1234 ;
  assign n1236 = x318 & n771 ;
  assign n1237 = x446 & ~n771 ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = ( n1232 & n1235 ) | ( n1232 & ~n1238 ) | ( n1235 & ~n1238 ) ;
  assign n1240 = x319 & n771 ;
  assign n1241 = x447 & ~n771 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = x63 & n640 ;
  assign n1244 = x191 & ~n640 ;
  assign n1245 = n1243 | n1244 ;
  assign n1246 = ( n1239 & ~n1242 ) | ( n1239 & n1245 ) | ( ~n1242 & n1245 ) ;
  assign n1247 = x64 & n640 ;
  assign n1248 = x192 & ~n640 ;
  assign n1249 = n1247 | n1248 ;
  assign n1250 = x320 & n771 ;
  assign n1251 = x448 & ~n771 ;
  assign n1252 = n1250 | n1251 ;
  assign n1253 = ( n1246 & n1249 ) | ( n1246 & ~n1252 ) | ( n1249 & ~n1252 ) ;
  assign n1254 = x321 & n771 ;
  assign n1255 = x449 & ~n771 ;
  assign n1256 = n1254 | n1255 ;
  assign n1257 = x65 & n640 ;
  assign n1258 = x193 & ~n640 ;
  assign n1259 = n1257 | n1258 ;
  assign n1260 = ( n1253 & ~n1256 ) | ( n1253 & n1259 ) | ( ~n1256 & n1259 ) ;
  assign n1261 = x322 & n771 ;
  assign n1262 = x450 & ~n771 ;
  assign n1263 = n1261 | n1262 ;
  assign n1264 = x66 & n640 ;
  assign n1265 = x194 & ~n640 ;
  assign n1266 = n1264 | n1265 ;
  assign n1267 = ( n1260 & ~n1263 ) | ( n1260 & n1266 ) | ( ~n1263 & n1266 ) ;
  assign n1268 = x67 & n640 ;
  assign n1269 = x195 & ~n640 ;
  assign n1270 = n1268 | n1269 ;
  assign n1271 = x323 & n771 ;
  assign n1272 = x451 & ~n771 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = ( n1267 & n1270 ) | ( n1267 & ~n1273 ) | ( n1270 & ~n1273 ) ;
  assign n1275 = x324 & n771 ;
  assign n1276 = x452 & ~n771 ;
  assign n1277 = n1275 | n1276 ;
  assign n1278 = x68 & n640 ;
  assign n1279 = x196 & ~n640 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = ( n1274 & ~n1277 ) | ( n1274 & n1280 ) | ( ~n1277 & n1280 ) ;
  assign n1282 = x325 & n771 ;
  assign n1283 = x453 & ~n771 ;
  assign n1284 = n1282 | n1283 ;
  assign n1285 = x69 & n640 ;
  assign n1286 = x197 & ~n640 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = ( n1281 & ~n1284 ) | ( n1281 & n1287 ) | ( ~n1284 & n1287 ) ;
  assign n1289 = x326 & n771 ;
  assign n1290 = x454 & ~n771 ;
  assign n1291 = n1289 | n1290 ;
  assign n1292 = x70 & n640 ;
  assign n1293 = x198 & ~n640 ;
  assign n1294 = n1292 | n1293 ;
  assign n1295 = ( n1288 & ~n1291 ) | ( n1288 & n1294 ) | ( ~n1291 & n1294 ) ;
  assign n1296 = x71 & n640 ;
  assign n1297 = x199 & ~n640 ;
  assign n1298 = n1296 | n1297 ;
  assign n1299 = x327 & n771 ;
  assign n1300 = x455 & ~n771 ;
  assign n1301 = n1299 | n1300 ;
  assign n1302 = ( n1295 & n1298 ) | ( n1295 & ~n1301 ) | ( n1298 & ~n1301 ) ;
  assign n1303 = x328 & n771 ;
  assign n1304 = x456 & ~n771 ;
  assign n1305 = n1303 | n1304 ;
  assign n1306 = x72 & n640 ;
  assign n1307 = x200 & ~n640 ;
  assign n1308 = n1306 | n1307 ;
  assign n1309 = ( n1302 & ~n1305 ) | ( n1302 & n1308 ) | ( ~n1305 & n1308 ) ;
  assign n1310 = x73 & n640 ;
  assign n1311 = x201 & ~n640 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = x329 & n771 ;
  assign n1314 = x457 & ~n771 ;
  assign n1315 = n1313 | n1314 ;
  assign n1316 = ( n1309 & n1312 ) | ( n1309 & ~n1315 ) | ( n1312 & ~n1315 ) ;
  assign n1317 = ( ~n798 & n801 ) | ( ~n798 & n1316 ) | ( n801 & n1316 ) ;
  assign n1318 = x75 & n640 ;
  assign n1319 = x203 & ~n640 ;
  assign n1320 = n1318 | n1319 ;
  assign n1321 = x331 & n771 ;
  assign n1322 = x459 & ~n771 ;
  assign n1323 = n1321 | n1322 ;
  assign n1324 = ( n1317 & n1320 ) | ( n1317 & ~n1323 ) | ( n1320 & ~n1323 ) ;
  assign n1325 = x76 & n640 ;
  assign n1326 = x204 & ~n640 ;
  assign n1327 = n1325 | n1326 ;
  assign n1328 = x332 & n771 ;
  assign n1329 = x460 & ~n771 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = ( n1324 & n1327 ) | ( n1324 & ~n1330 ) | ( n1327 & ~n1330 ) ;
  assign n1332 = x333 & n771 ;
  assign n1333 = x461 & ~n771 ;
  assign n1334 = n1332 | n1333 ;
  assign n1335 = x77 & n640 ;
  assign n1336 = x205 & ~n640 ;
  assign n1337 = n1335 | n1336 ;
  assign n1338 = ( n1331 & ~n1334 ) | ( n1331 & n1337 ) | ( ~n1334 & n1337 ) ;
  assign n1339 = x78 & n640 ;
  assign n1340 = x206 & ~n640 ;
  assign n1341 = n1339 | n1340 ;
  assign n1342 = x334 & n771 ;
  assign n1343 = x462 & ~n771 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = ( n1338 & n1341 ) | ( n1338 & ~n1344 ) | ( n1341 & ~n1344 ) ;
  assign n1346 = x335 & n771 ;
  assign n1347 = x463 & ~n771 ;
  assign n1348 = n1346 | n1347 ;
  assign n1349 = x79 & n640 ;
  assign n1350 = x207 & ~n640 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = ( n1345 & ~n1348 ) | ( n1345 & n1351 ) | ( ~n1348 & n1351 ) ;
  assign n1353 = x336 & n771 ;
  assign n1354 = x464 & ~n771 ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = x80 & n640 ;
  assign n1357 = x208 & ~n640 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = ( n1352 & ~n1355 ) | ( n1352 & n1358 ) | ( ~n1355 & n1358 ) ;
  assign n1360 = x81 & n640 ;
  assign n1361 = x209 & ~n640 ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = x337 & n771 ;
  assign n1364 = x465 & ~n771 ;
  assign n1365 = n1363 | n1364 ;
  assign n1366 = ( n1359 & n1362 ) | ( n1359 & ~n1365 ) | ( n1362 & ~n1365 ) ;
  assign n1367 = x82 & n640 ;
  assign n1368 = x210 & ~n640 ;
  assign n1369 = n1367 | n1368 ;
  assign n1370 = x338 & n771 ;
  assign n1371 = x466 & ~n771 ;
  assign n1372 = n1370 | n1371 ;
  assign n1373 = ( n1366 & n1369 ) | ( n1366 & ~n1372 ) | ( n1369 & ~n1372 ) ;
  assign n1374 = x83 & n640 ;
  assign n1375 = x211 & ~n640 ;
  assign n1376 = n1374 | n1375 ;
  assign n1377 = x339 & n771 ;
  assign n1378 = x467 & ~n771 ;
  assign n1379 = n1377 | n1378 ;
  assign n1380 = ( n1373 & n1376 ) | ( n1373 & ~n1379 ) | ( n1376 & ~n1379 ) ;
  assign n1381 = x340 & n771 ;
  assign n1382 = x468 & ~n771 ;
  assign n1383 = n1381 | n1382 ;
  assign n1384 = x84 & n640 ;
  assign n1385 = x212 & ~n640 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = ( n1380 & ~n1383 ) | ( n1380 & n1386 ) | ( ~n1383 & n1386 ) ;
  assign n1388 = x85 & n640 ;
  assign n1389 = x213 & ~n640 ;
  assign n1390 = n1388 | n1389 ;
  assign n1391 = x341 & n771 ;
  assign n1392 = x469 & ~n771 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = ( n1387 & n1390 ) | ( n1387 & ~n1393 ) | ( n1390 & ~n1393 ) ;
  assign n1395 = x342 & n771 ;
  assign n1396 = x470 & ~n771 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = x86 & n640 ;
  assign n1399 = x214 & ~n640 ;
  assign n1400 = n1398 | n1399 ;
  assign n1401 = ( n1394 & ~n1397 ) | ( n1394 & n1400 ) | ( ~n1397 & n1400 ) ;
  assign n1402 = x343 & n771 ;
  assign n1403 = x471 & ~n771 ;
  assign n1404 = n1402 | n1403 ;
  assign n1405 = x87 & n640 ;
  assign n1406 = x215 & ~n640 ;
  assign n1407 = n1405 | n1406 ;
  assign n1408 = ( n1401 & ~n1404 ) | ( n1401 & n1407 ) | ( ~n1404 & n1407 ) ;
  assign n1409 = x88 & n640 ;
  assign n1410 = x216 & ~n640 ;
  assign n1411 = n1409 | n1410 ;
  assign n1412 = x344 & n771 ;
  assign n1413 = x472 & ~n771 ;
  assign n1414 = n1412 | n1413 ;
  assign n1415 = ( n1408 & n1411 ) | ( n1408 & ~n1414 ) | ( n1411 & ~n1414 ) ;
  assign n1416 = ( ~n792 & n795 ) | ( ~n792 & n1415 ) | ( n795 & n1415 ) ;
  assign n1417 = x90 & n640 ;
  assign n1418 = x218 & ~n640 ;
  assign n1419 = n1417 | n1418 ;
  assign n1420 = x346 & n771 ;
  assign n1421 = x474 & ~n771 ;
  assign n1422 = n1420 | n1421 ;
  assign n1423 = ( n1416 & n1419 ) | ( n1416 & ~n1422 ) | ( n1419 & ~n1422 ) ;
  assign n1424 = x91 & n640 ;
  assign n1425 = x219 & ~n640 ;
  assign n1426 = n1424 | n1425 ;
  assign n1427 = x347 & n771 ;
  assign n1428 = x475 & ~n771 ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = ( n1423 & n1426 ) | ( n1423 & ~n1429 ) | ( n1426 & ~n1429 ) ;
  assign n1431 = x348 & n771 ;
  assign n1432 = x476 & ~n771 ;
  assign n1433 = n1431 | n1432 ;
  assign n1434 = x92 & n640 ;
  assign n1435 = x220 & ~n640 ;
  assign n1436 = n1434 | n1435 ;
  assign n1437 = ( n1430 & ~n1433 ) | ( n1430 & n1436 ) | ( ~n1433 & n1436 ) ;
  assign n1438 = ( ~n786 & n789 ) | ( ~n786 & n1437 ) | ( n789 & n1437 ) ;
  assign n1439 = x350 & n771 ;
  assign n1440 = x478 & ~n771 ;
  assign n1441 = n1439 | n1440 ;
  assign n1442 = x94 & n640 ;
  assign n1443 = x222 & ~n640 ;
  assign n1444 = n1442 | n1443 ;
  assign n1445 = ( n1438 & ~n1441 ) | ( n1438 & n1444 ) | ( ~n1441 & n1444 ) ;
  assign n1446 = x95 & n640 ;
  assign n1447 = x223 & ~n640 ;
  assign n1448 = n1446 | n1447 ;
  assign n1449 = x351 & n771 ;
  assign n1450 = x479 & ~n771 ;
  assign n1451 = n1449 | n1450 ;
  assign n1452 = ( n1445 & n1448 ) | ( n1445 & ~n1451 ) | ( n1448 & ~n1451 ) ;
  assign n1453 = x96 & n640 ;
  assign n1454 = x224 & ~n640 ;
  assign n1455 = n1453 | n1454 ;
  assign n1456 = x352 & n771 ;
  assign n1457 = x480 & ~n771 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = ( n1452 & n1455 ) | ( n1452 & ~n1458 ) | ( n1455 & ~n1458 ) ;
  assign n1460 = x353 & n771 ;
  assign n1461 = x481 & ~n771 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = x97 & n640 ;
  assign n1464 = x225 & ~n640 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = ( n1459 & ~n1462 ) | ( n1459 & n1465 ) | ( ~n1462 & n1465 ) ;
  assign n1467 = x98 & n640 ;
  assign n1468 = x226 & ~n640 ;
  assign n1469 = n1467 | n1468 ;
  assign n1470 = x354 & n771 ;
  assign n1471 = x482 & ~n771 ;
  assign n1472 = n1470 | n1471 ;
  assign n1473 = ( n1466 & n1469 ) | ( n1466 & ~n1472 ) | ( n1469 & ~n1472 ) ;
  assign n1474 = x355 & n771 ;
  assign n1475 = x483 & ~n771 ;
  assign n1476 = n1474 | n1475 ;
  assign n1477 = x99 & n640 ;
  assign n1478 = x227 & ~n640 ;
  assign n1479 = n1477 | n1478 ;
  assign n1480 = ( n1473 & ~n1476 ) | ( n1473 & n1479 ) | ( ~n1476 & n1479 ) ;
  assign n1481 = x356 & n771 ;
  assign n1482 = x484 & ~n771 ;
  assign n1483 = n1481 | n1482 ;
  assign n1484 = x100 & n640 ;
  assign n1485 = x228 & ~n640 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = ( n1480 & ~n1483 ) | ( n1480 & n1486 ) | ( ~n1483 & n1486 ) ;
  assign n1488 = x101 & n640 ;
  assign n1489 = x229 & ~n640 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = x357 & n771 ;
  assign n1492 = x485 & ~n771 ;
  assign n1493 = n1491 | n1492 ;
  assign n1494 = ( n1487 & n1490 ) | ( n1487 & ~n1493 ) | ( n1490 & ~n1493 ) ;
  assign n1495 = x358 & n771 ;
  assign n1496 = x486 & ~n771 ;
  assign n1497 = n1495 | n1496 ;
  assign n1498 = x102 & n640 ;
  assign n1499 = x230 & ~n640 ;
  assign n1500 = n1498 | n1499 ;
  assign n1501 = ( n1494 & ~n1497 ) | ( n1494 & n1500 ) | ( ~n1497 & n1500 ) ;
  assign n1502 = x359 & n771 ;
  assign n1503 = x487 & ~n771 ;
  assign n1504 = n1502 | n1503 ;
  assign n1505 = x103 & n640 ;
  assign n1506 = x231 & ~n640 ;
  assign n1507 = n1505 | n1506 ;
  assign n1508 = ( n1501 & ~n1504 ) | ( n1501 & n1507 ) | ( ~n1504 & n1507 ) ;
  assign n1509 = x360 & n771 ;
  assign n1510 = x488 & ~n771 ;
  assign n1511 = n1509 | n1510 ;
  assign n1512 = x104 & n640 ;
  assign n1513 = x232 & ~n640 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = ( n1508 & ~n1511 ) | ( n1508 & n1514 ) | ( ~n1511 & n1514 ) ;
  assign n1516 = x361 & n771 ;
  assign n1517 = x489 & ~n771 ;
  assign n1518 = n1516 | n1517 ;
  assign n1519 = x105 & n640 ;
  assign n1520 = x233 & ~n640 ;
  assign n1521 = n1519 | n1520 ;
  assign n1522 = ( n1515 & ~n1518 ) | ( n1515 & n1521 ) | ( ~n1518 & n1521 ) ;
  assign n1523 = x362 & n771 ;
  assign n1524 = x490 & ~n771 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = x106 & n640 ;
  assign n1527 = x234 & ~n640 ;
  assign n1528 = n1526 | n1527 ;
  assign n1529 = ( n1522 & ~n1525 ) | ( n1522 & n1528 ) | ( ~n1525 & n1528 ) ;
  assign n1530 = x107 & n640 ;
  assign n1531 = x235 & ~n640 ;
  assign n1532 = n1530 | n1531 ;
  assign n1533 = x363 & n771 ;
  assign n1534 = x491 & ~n771 ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = ( n1529 & n1532 ) | ( n1529 & ~n1535 ) | ( n1532 & ~n1535 ) ;
  assign n1537 = x364 & n771 ;
  assign n1538 = x492 & ~n771 ;
  assign n1539 = n1537 | n1538 ;
  assign n1540 = x108 & n640 ;
  assign n1541 = x236 & ~n640 ;
  assign n1542 = n1540 | n1541 ;
  assign n1543 = ( n1536 & ~n1539 ) | ( n1536 & n1542 ) | ( ~n1539 & n1542 ) ;
  assign n1544 = x109 & n640 ;
  assign n1545 = x237 & ~n640 ;
  assign n1546 = n1544 | n1545 ;
  assign n1547 = x365 & n771 ;
  assign n1548 = x493 & ~n771 ;
  assign n1549 = n1547 | n1548 ;
  assign n1550 = ( n1543 & n1546 ) | ( n1543 & ~n1549 ) | ( n1546 & ~n1549 ) ;
  assign n1551 = x366 & n771 ;
  assign n1552 = x494 & ~n771 ;
  assign n1553 = n1551 | n1552 ;
  assign n1554 = x110 & n640 ;
  assign n1555 = x238 & ~n640 ;
  assign n1556 = n1554 | n1555 ;
  assign n1557 = ( n1550 & ~n1553 ) | ( n1550 & n1556 ) | ( ~n1553 & n1556 ) ;
  assign n1558 = x111 & n640 ;
  assign n1559 = x239 & ~n640 ;
  assign n1560 = n1558 | n1559 ;
  assign n1561 = x367 & n771 ;
  assign n1562 = x495 & ~n771 ;
  assign n1563 = n1561 | n1562 ;
  assign n1564 = ( n1557 & n1560 ) | ( n1557 & ~n1563 ) | ( n1560 & ~n1563 ) ;
  assign n1565 = ( ~n780 & n783 ) | ( ~n780 & n1564 ) | ( n783 & n1564 ) ;
  assign n1566 = x113 & n640 ;
  assign n1567 = x241 & ~n640 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = x369 & n771 ;
  assign n1570 = x497 & ~n771 ;
  assign n1571 = n1569 | n1570 ;
  assign n1572 = ( n1565 & n1568 ) | ( n1565 & ~n1571 ) | ( n1568 & ~n1571 ) ;
  assign n1573 = x114 & n640 ;
  assign n1574 = x242 & ~n640 ;
  assign n1575 = n1573 | n1574 ;
  assign n1576 = x370 & n771 ;
  assign n1577 = x498 & ~n771 ;
  assign n1578 = n1576 | n1577 ;
  assign n1579 = ( n1572 & n1575 ) | ( n1572 & ~n1578 ) | ( n1575 & ~n1578 ) ;
  assign n1580 = x371 & n771 ;
  assign n1581 = x499 & ~n771 ;
  assign n1582 = n1580 | n1581 ;
  assign n1583 = x115 & n640 ;
  assign n1584 = x243 & ~n640 ;
  assign n1585 = n1583 | n1584 ;
  assign n1586 = ( n1579 & ~n1582 ) | ( n1579 & n1585 ) | ( ~n1582 & n1585 ) ;
  assign n1587 = x372 & n771 ;
  assign n1588 = x500 & ~n771 ;
  assign n1589 = n1587 | n1588 ;
  assign n1590 = x116 & n640 ;
  assign n1591 = x244 & ~n640 ;
  assign n1592 = n1590 | n1591 ;
  assign n1593 = ( n1586 & ~n1589 ) | ( n1586 & n1592 ) | ( ~n1589 & n1592 ) ;
  assign n1594 = x117 & n640 ;
  assign n1595 = x245 & ~n640 ;
  assign n1596 = n1594 | n1595 ;
  assign n1597 = x373 & n771 ;
  assign n1598 = x501 & ~n771 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = ( n1593 & n1596 ) | ( n1593 & ~n1599 ) | ( n1596 & ~n1599 ) ;
  assign n1601 = x118 & n640 ;
  assign n1602 = x246 & ~n640 ;
  assign n1603 = n1601 | n1602 ;
  assign n1604 = x374 & n771 ;
  assign n1605 = x502 & ~n771 ;
  assign n1606 = n1604 | n1605 ;
  assign n1607 = ( n1600 & n1603 ) | ( n1600 & ~n1606 ) | ( n1603 & ~n1606 ) ;
  assign n1608 = ( ~n774 & n777 ) | ( ~n774 & n1607 ) | ( n777 & n1607 ) ;
  assign n1609 = x120 & n640 ;
  assign n1610 = x248 & ~n640 ;
  assign n1611 = n1609 | n1610 ;
  assign n1612 = x376 & n771 ;
  assign n1613 = x504 & ~n771 ;
  assign n1614 = n1612 | n1613 ;
  assign n1615 = ( n1608 & n1611 ) | ( n1608 & ~n1614 ) | ( n1611 & ~n1614 ) ;
  assign n1616 = x121 & n640 ;
  assign n1617 = x249 & ~n640 ;
  assign n1618 = n1616 | n1617 ;
  assign n1619 = x377 & n771 ;
  assign n1620 = x505 & ~n771 ;
  assign n1621 = n1619 | n1620 ;
  assign n1622 = ( n1615 & n1618 ) | ( n1615 & ~n1621 ) | ( n1618 & ~n1621 ) ;
  assign n1623 = x122 & n640 ;
  assign n1624 = x250 & ~n640 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = x378 & n771 ;
  assign n1627 = x506 & ~n771 ;
  assign n1628 = n1626 | n1627 ;
  assign n1629 = ( n1622 & n1625 ) | ( n1622 & ~n1628 ) | ( n1625 & ~n1628 ) ;
  assign n1630 = x379 & n771 ;
  assign n1631 = x507 & ~n771 ;
  assign n1632 = n1630 | n1631 ;
  assign n1633 = x123 & n640 ;
  assign n1634 = x251 & ~n640 ;
  assign n1635 = n1633 | n1634 ;
  assign n1636 = ( n1629 & ~n1632 ) | ( n1629 & n1635 ) | ( ~n1632 & n1635 ) ;
  assign n1637 = x124 & n640 ;
  assign n1638 = x252 & ~n640 ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = x380 & n771 ;
  assign n1641 = x508 & ~n771 ;
  assign n1642 = n1640 | n1641 ;
  assign n1643 = ( n1636 & n1639 ) | ( n1636 & ~n1642 ) | ( n1639 & ~n1642 ) ;
  assign n1644 = x125 & n640 ;
  assign n1645 = x253 & ~n640 ;
  assign n1646 = n1644 | n1645 ;
  assign n1647 = x381 & n771 ;
  assign n1648 = x509 & ~n771 ;
  assign n1649 = n1647 | n1648 ;
  assign n1650 = ( n1643 & n1646 ) | ( n1643 & ~n1649 ) | ( n1646 & ~n1649 ) ;
  assign n1651 = x126 & n640 ;
  assign n1652 = x254 & ~n640 ;
  assign n1653 = n1651 | n1652 ;
  assign n1654 = x382 & n771 ;
  assign n1655 = x510 & ~n771 ;
  assign n1656 = n1654 | n1655 ;
  assign n1657 = ( n1650 & n1653 ) | ( n1650 & ~n1656 ) | ( n1653 & ~n1656 ) ;
  assign n1658 = x127 & x255 ;
  assign n1659 = x383 & x511 ;
  assign n1660 = ( n1657 & ~n1658 ) | ( n1657 & n1659 ) | ( ~n1658 & n1659 ) ;
  assign n1661 = ~n643 & n1660 ;
  assign n1662 = n816 | n1660 ;
  assign n1663 = ~n1661 & n1662 ;
  assign n1664 = ~n810 & n1660 ;
  assign n1665 = n813 | n1660 ;
  assign n1666 = ~n1664 & n1665 ;
  assign n1667 = n821 | n1660 ;
  assign n1668 = ~n824 & n1660 ;
  assign n1669 = n1667 & ~n1668 ;
  assign n1670 = ~n828 & n1660 ;
  assign n1671 = n831 | n1660 ;
  assign n1672 = ~n1670 & n1671 ;
  assign n1673 = n804 | n1660 ;
  assign n1674 = ~n807 & n1660 ;
  assign n1675 = n1673 & ~n1674 ;
  assign n1676 = ~n836 & n1660 ;
  assign n1677 = n839 | n1660 ;
  assign n1678 = ~n1676 & n1677 ;
  assign n1679 = ~n843 & n1660 ;
  assign n1680 = n846 | n1660 ;
  assign n1681 = ~n1679 & n1680 ;
  assign n1682 = n850 | n1660 ;
  assign n1683 = ~n853 & n1660 ;
  assign n1684 = n1682 & ~n1683 ;
  assign n1685 = n857 | n1660 ;
  assign n1686 = ~n860 & n1660 ;
  assign n1687 = n1685 & ~n1686 ;
  assign n1688 = ~n864 & n1660 ;
  assign n1689 = n867 | n1660 ;
  assign n1690 = ~n1688 & n1689 ;
  assign n1691 = ~n871 & n1660 ;
  assign n1692 = n874 | n1660 ;
  assign n1693 = ~n1691 & n1692 ;
  assign n1694 = n878 | n1660 ;
  assign n1695 = ~n881 & n1660 ;
  assign n1696 = n1694 & ~n1695 ;
  assign n1697 = ~n885 & n1660 ;
  assign n1698 = n888 | n1660 ;
  assign n1699 = ~n1697 & n1698 ;
  assign n1700 = n892 | n1660 ;
  assign n1701 = ~n895 & n1660 ;
  assign n1702 = n1700 & ~n1701 ;
  assign n1703 = n899 | n1660 ;
  assign n1704 = ~n902 & n1660 ;
  assign n1705 = n1703 & ~n1704 ;
  assign n1706 = ~n906 & n1660 ;
  assign n1707 = n909 | n1660 ;
  assign n1708 = ~n1706 & n1707 ;
  assign n1709 = n913 | n1660 ;
  assign n1710 = ~n916 & n1660 ;
  assign n1711 = n1709 & ~n1710 ;
  assign n1712 = n920 | n1660 ;
  assign n1713 = ~n923 & n1660 ;
  assign n1714 = n1712 & ~n1713 ;
  assign n1715 = ~n927 & n1660 ;
  assign n1716 = n930 | n1660 ;
  assign n1717 = ~n1715 & n1716 ;
  assign n1718 = ~n934 & n1660 ;
  assign n1719 = n937 | n1660 ;
  assign n1720 = ~n1718 & n1719 ;
  assign n1721 = n941 | n1660 ;
  assign n1722 = ~n944 & n1660 ;
  assign n1723 = n1721 & ~n1722 ;
  assign n1724 = ~n948 & n1660 ;
  assign n1725 = n951 | n1660 ;
  assign n1726 = ~n1724 & n1725 ;
  assign n1727 = n955 | n1660 ;
  assign n1728 = ~n958 & n1660 ;
  assign n1729 = n1727 & ~n1728 ;
  assign n1730 = n962 | n1660 ;
  assign n1731 = ~n965 & n1660 ;
  assign n1732 = n1730 & ~n1731 ;
  assign n1733 = n969 | n1660 ;
  assign n1734 = ~n972 & n1660 ;
  assign n1735 = n1733 & ~n1734 ;
  assign n1736 = n976 | n1660 ;
  assign n1737 = ~n979 & n1660 ;
  assign n1738 = n1736 & ~n1737 ;
  assign n1739 = ~n983 & n1660 ;
  assign n1740 = n986 | n1660 ;
  assign n1741 = ~n1739 & n1740 ;
  assign n1742 = n990 | n1660 ;
  assign n1743 = ~n993 & n1660 ;
  assign n1744 = n1742 & ~n1743 ;
  assign n1745 = n997 | n1660 ;
  assign n1746 = ~n1000 & n1660 ;
  assign n1747 = n1745 & ~n1746 ;
  assign n1748 = ~n1004 & n1660 ;
  assign n1749 = n1007 | n1660 ;
  assign n1750 = ~n1748 & n1749 ;
  assign n1751 = ~n1011 & n1660 ;
  assign n1752 = n1014 | n1660 ;
  assign n1753 = ~n1751 & n1752 ;
  assign n1754 = n1018 | n1660 ;
  assign n1755 = ~n1021 & n1660 ;
  assign n1756 = n1754 & ~n1755 ;
  assign n1757 = n1025 | n1660 ;
  assign n1758 = ~n1028 & n1660 ;
  assign n1759 = n1757 & ~n1758 ;
  assign n1760 = ~n1032 & n1660 ;
  assign n1761 = n1035 | n1660 ;
  assign n1762 = ~n1760 & n1761 ;
  assign n1763 = n1039 | n1660 ;
  assign n1764 = ~n1042 & n1660 ;
  assign n1765 = n1763 & ~n1764 ;
  assign n1766 = ~n1046 & n1660 ;
  assign n1767 = n1049 | n1660 ;
  assign n1768 = ~n1766 & n1767 ;
  assign n1769 = n1053 | n1660 ;
  assign n1770 = ~n1056 & n1660 ;
  assign n1771 = n1769 & ~n1770 ;
  assign n1772 = n1060 | n1660 ;
  assign n1773 = ~n1063 & n1660 ;
  assign n1774 = n1772 & ~n1773 ;
  assign n1775 = n1067 | n1660 ;
  assign n1776 = ~n1070 & n1660 ;
  assign n1777 = n1775 & ~n1776 ;
  assign n1778 = ~n1074 & n1660 ;
  assign n1779 = n1077 | n1660 ;
  assign n1780 = ~n1778 & n1779 ;
  assign n1781 = n1081 | n1660 ;
  assign n1782 = ~n1084 & n1660 ;
  assign n1783 = n1781 & ~n1782 ;
  assign n1784 = n1088 | n1660 ;
  assign n1785 = ~n1091 & n1660 ;
  assign n1786 = n1784 & ~n1785 ;
  assign n1787 = ~n1095 & n1660 ;
  assign n1788 = n1098 | n1660 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = ~n1102 & n1660 ;
  assign n1791 = n1105 | n1660 ;
  assign n1792 = ~n1790 & n1791 ;
  assign n1793 = ~n1109 & n1660 ;
  assign n1794 = n1112 | n1660 ;
  assign n1795 = ~n1793 & n1794 ;
  assign n1796 = n1116 | n1660 ;
  assign n1797 = ~n1119 & n1660 ;
  assign n1798 = n1796 & ~n1797 ;
  assign n1799 = n1123 | n1660 ;
  assign n1800 = ~n1126 & n1660 ;
  assign n1801 = n1799 & ~n1800 ;
  assign n1802 = ~n1130 & n1660 ;
  assign n1803 = n1133 | n1660 ;
  assign n1804 = ~n1802 & n1803 ;
  assign n1805 = n1137 | n1660 ;
  assign n1806 = ~n1140 & n1660 ;
  assign n1807 = n1805 & ~n1806 ;
  assign n1808 = n1144 | n1660 ;
  assign n1809 = ~n1147 & n1660 ;
  assign n1810 = n1808 & ~n1809 ;
  assign n1811 = ~n1151 & n1660 ;
  assign n1812 = n1154 | n1660 ;
  assign n1813 = ~n1811 & n1812 ;
  assign n1814 = n1158 | n1660 ;
  assign n1815 = ~n1161 & n1660 ;
  assign n1816 = n1814 & ~n1815 ;
  assign n1817 = n1165 | n1660 ;
  assign n1818 = ~n1168 & n1660 ;
  assign n1819 = n1817 & ~n1818 ;
  assign n1820 = ~n1172 & n1660 ;
  assign n1821 = n1175 | n1660 ;
  assign n1822 = ~n1820 & n1821 ;
  assign n1823 = n1179 | n1660 ;
  assign n1824 = ~n1182 & n1660 ;
  assign n1825 = n1823 & ~n1824 ;
  assign n1826 = n1186 | n1660 ;
  assign n1827 = ~n1189 & n1660 ;
  assign n1828 = n1826 & ~n1827 ;
  assign n1829 = ~n1193 & n1660 ;
  assign n1830 = n1196 | n1660 ;
  assign n1831 = ~n1829 & n1830 ;
  assign n1832 = ~n1200 & n1660 ;
  assign n1833 = n1203 | n1660 ;
  assign n1834 = ~n1832 & n1833 ;
  assign n1835 = ~n1207 & n1660 ;
  assign n1836 = n1210 | n1660 ;
  assign n1837 = ~n1835 & n1836 ;
  assign n1838 = n1214 | n1660 ;
  assign n1839 = ~n1217 & n1660 ;
  assign n1840 = n1838 & ~n1839 ;
  assign n1841 = ~n1221 & n1660 ;
  assign n1842 = n1224 | n1660 ;
  assign n1843 = ~n1841 & n1842 ;
  assign n1844 = n1228 | n1660 ;
  assign n1845 = ~n1231 & n1660 ;
  assign n1846 = n1844 & ~n1845 ;
  assign n1847 = ~n1235 & n1660 ;
  assign n1848 = n1238 | n1660 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1850 = n1242 | n1660 ;
  assign n1851 = ~n1245 & n1660 ;
  assign n1852 = n1850 & ~n1851 ;
  assign n1853 = ~n1249 & n1660 ;
  assign n1854 = n1252 | n1660 ;
  assign n1855 = ~n1853 & n1854 ;
  assign n1856 = n1256 | n1660 ;
  assign n1857 = ~n1259 & n1660 ;
  assign n1858 = n1856 & ~n1857 ;
  assign n1859 = n1263 | n1660 ;
  assign n1860 = ~n1266 & n1660 ;
  assign n1861 = n1859 & ~n1860 ;
  assign n1862 = ~n1270 & n1660 ;
  assign n1863 = n1273 | n1660 ;
  assign n1864 = ~n1862 & n1863 ;
  assign n1865 = n1277 | n1660 ;
  assign n1866 = ~n1280 & n1660 ;
  assign n1867 = n1865 & ~n1866 ;
  assign n1868 = n1284 | n1660 ;
  assign n1869 = ~n1287 & n1660 ;
  assign n1870 = n1868 & ~n1869 ;
  assign n1871 = n1291 | n1660 ;
  assign n1872 = ~n1294 & n1660 ;
  assign n1873 = n1871 & ~n1872 ;
  assign n1874 = ~n1298 & n1660 ;
  assign n1875 = n1301 | n1660 ;
  assign n1876 = ~n1874 & n1875 ;
  assign n1877 = n1305 | n1660 ;
  assign n1878 = ~n1308 & n1660 ;
  assign n1879 = n1877 & ~n1878 ;
  assign n1880 = ~n1312 & n1660 ;
  assign n1881 = n1315 | n1660 ;
  assign n1882 = ~n1880 & n1881 ;
  assign n1883 = n798 | n1660 ;
  assign n1884 = ~n801 & n1660 ;
  assign n1885 = n1883 & ~n1884 ;
  assign n1886 = ~n1320 & n1660 ;
  assign n1887 = n1323 | n1660 ;
  assign n1888 = ~n1886 & n1887 ;
  assign n1889 = ~n1327 & n1660 ;
  assign n1890 = n1330 | n1660 ;
  assign n1891 = ~n1889 & n1890 ;
  assign n1892 = n1334 | n1660 ;
  assign n1893 = ~n1337 & n1660 ;
  assign n1894 = n1892 & ~n1893 ;
  assign n1895 = ~n1341 & n1660 ;
  assign n1896 = n1344 | n1660 ;
  assign n1897 = ~n1895 & n1896 ;
  assign n1898 = n1348 | n1660 ;
  assign n1899 = ~n1351 & n1660 ;
  assign n1900 = n1898 & ~n1899 ;
  assign n1901 = n1355 | n1660 ;
  assign n1902 = ~n1358 & n1660 ;
  assign n1903 = n1901 & ~n1902 ;
  assign n1904 = ~n1362 & n1660 ;
  assign n1905 = n1365 | n1660 ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = ~n1369 & n1660 ;
  assign n1908 = n1372 | n1660 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1910 = ~n1376 & n1660 ;
  assign n1911 = n1379 | n1660 ;
  assign n1912 = ~n1910 & n1911 ;
  assign n1913 = n1383 | n1660 ;
  assign n1914 = ~n1386 & n1660 ;
  assign n1915 = n1913 & ~n1914 ;
  assign n1916 = ~n1390 & n1660 ;
  assign n1917 = n1393 | n1660 ;
  assign n1918 = ~n1916 & n1917 ;
  assign n1919 = n1397 | n1660 ;
  assign n1920 = ~n1400 & n1660 ;
  assign n1921 = n1919 & ~n1920 ;
  assign n1922 = n1404 | n1660 ;
  assign n1923 = ~n1407 & n1660 ;
  assign n1924 = n1922 & ~n1923 ;
  assign n1925 = ~n1411 & n1660 ;
  assign n1926 = n1414 | n1660 ;
  assign n1927 = ~n1925 & n1926 ;
  assign n1928 = n792 | n1660 ;
  assign n1929 = ~n795 & n1660 ;
  assign n1930 = n1928 & ~n1929 ;
  assign n1931 = ~n1419 & n1660 ;
  assign n1932 = n1422 | n1660 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1934 = ~n1426 & n1660 ;
  assign n1935 = n1429 | n1660 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = n1433 | n1660 ;
  assign n1938 = ~n1436 & n1660 ;
  assign n1939 = n1937 & ~n1938 ;
  assign n1940 = n786 | n1660 ;
  assign n1941 = ~n789 & n1660 ;
  assign n1942 = n1940 & ~n1941 ;
  assign n1943 = n1441 | n1660 ;
  assign n1944 = ~n1444 & n1660 ;
  assign n1945 = n1943 & ~n1944 ;
  assign n1946 = ~n1448 & n1660 ;
  assign n1947 = n1451 | n1660 ;
  assign n1948 = ~n1946 & n1947 ;
  assign n1949 = ~n1455 & n1660 ;
  assign n1950 = n1458 | n1660 ;
  assign n1951 = ~n1949 & n1950 ;
  assign n1952 = n1462 | n1660 ;
  assign n1953 = ~n1465 & n1660 ;
  assign n1954 = n1952 & ~n1953 ;
  assign n1955 = ~n1469 & n1660 ;
  assign n1956 = n1472 | n1660 ;
  assign n1957 = ~n1955 & n1956 ;
  assign n1958 = n1476 | n1660 ;
  assign n1959 = ~n1479 & n1660 ;
  assign n1960 = n1958 & ~n1959 ;
  assign n1961 = n1483 | n1660 ;
  assign n1962 = ~n1486 & n1660 ;
  assign n1963 = n1961 & ~n1962 ;
  assign n1964 = ~n1490 & n1660 ;
  assign n1965 = n1493 | n1660 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1967 = n1497 | n1660 ;
  assign n1968 = ~n1500 & n1660 ;
  assign n1969 = n1967 & ~n1968 ;
  assign n1970 = n1504 | n1660 ;
  assign n1971 = ~n1507 & n1660 ;
  assign n1972 = n1970 & ~n1971 ;
  assign n1973 = n1511 | n1660 ;
  assign n1974 = ~n1514 & n1660 ;
  assign n1975 = n1973 & ~n1974 ;
  assign n1976 = n1518 | n1660 ;
  assign n1977 = ~n1521 & n1660 ;
  assign n1978 = n1976 & ~n1977 ;
  assign n1979 = n1525 | n1660 ;
  assign n1980 = ~n1528 & n1660 ;
  assign n1981 = n1979 & ~n1980 ;
  assign n1982 = ~n1532 & n1660 ;
  assign n1983 = n1535 | n1660 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = n1539 | n1660 ;
  assign n1986 = ~n1542 & n1660 ;
  assign n1987 = n1985 & ~n1986 ;
  assign n1988 = ~n1546 & n1660 ;
  assign n1989 = n1549 | n1660 ;
  assign n1990 = ~n1988 & n1989 ;
  assign n1991 = n1553 | n1660 ;
  assign n1992 = ~n1556 & n1660 ;
  assign n1993 = n1991 & ~n1992 ;
  assign n1994 = ~n1560 & n1660 ;
  assign n1995 = n1563 | n1660 ;
  assign n1996 = ~n1994 & n1995 ;
  assign n1997 = n780 | n1660 ;
  assign n1998 = ~n783 & n1660 ;
  assign n1999 = n1997 & ~n1998 ;
  assign n2000 = ~n1568 & n1660 ;
  assign n2001 = n1571 | n1660 ;
  assign n2002 = ~n2000 & n2001 ;
  assign n2003 = ~n1575 & n1660 ;
  assign n2004 = n1578 | n1660 ;
  assign n2005 = ~n2003 & n2004 ;
  assign n2006 = n1582 | n1660 ;
  assign n2007 = ~n1585 & n1660 ;
  assign n2008 = n2006 & ~n2007 ;
  assign n2009 = n1589 | n1660 ;
  assign n2010 = ~n1592 & n1660 ;
  assign n2011 = n2009 & ~n2010 ;
  assign n2012 = ~n1596 & n1660 ;
  assign n2013 = n1599 | n1660 ;
  assign n2014 = ~n2012 & n2013 ;
  assign n2015 = ~n1603 & n1660 ;
  assign n2016 = n1606 | n1660 ;
  assign n2017 = ~n2015 & n2016 ;
  assign n2018 = n774 | n1660 ;
  assign n2019 = ~n777 & n1660 ;
  assign n2020 = n2018 & ~n2019 ;
  assign n2021 = ~n1611 & n1660 ;
  assign n2022 = n1614 | n1660 ;
  assign n2023 = ~n2021 & n2022 ;
  assign n2024 = ~n1618 & n1660 ;
  assign n2025 = n1621 | n1660 ;
  assign n2026 = ~n2024 & n2025 ;
  assign n2027 = ~n1625 & n1660 ;
  assign n2028 = n1628 | n1660 ;
  assign n2029 = ~n2027 & n2028 ;
  assign n2030 = n1632 | n1660 ;
  assign n2031 = ~n1635 & n1660 ;
  assign n2032 = n2030 & ~n2031 ;
  assign n2033 = ~n1639 & n1660 ;
  assign n2034 = n1642 | n1660 ;
  assign n2035 = ~n2033 & n2034 ;
  assign n2036 = ~n1646 & n1660 ;
  assign n2037 = n1649 | n1660 ;
  assign n2038 = ~n2036 & n2037 ;
  assign n2039 = ~n1653 & n1660 ;
  assign n2040 = n1656 | n1660 ;
  assign n2041 = ~n2039 & n2040 ;
  assign n2042 = n1658 & n1659 ;
  assign n2043 = ~n640 & n1660 ;
  assign n2044 = n771 | n1660 ;
  assign n2045 = ~n2043 & n2044 ;
  assign y0 = n1663 ;
  assign y1 = n1666 ;
  assign y2 = n1669 ;
  assign y3 = n1672 ;
  assign y4 = n1675 ;
  assign y5 = n1678 ;
  assign y6 = n1681 ;
  assign y7 = n1684 ;
  assign y8 = n1687 ;
  assign y9 = n1690 ;
  assign y10 = n1693 ;
  assign y11 = n1696 ;
  assign y12 = n1699 ;
  assign y13 = n1702 ;
  assign y14 = n1705 ;
  assign y15 = n1708 ;
  assign y16 = n1711 ;
  assign y17 = n1714 ;
  assign y18 = n1717 ;
  assign y19 = n1720 ;
  assign y20 = n1723 ;
  assign y21 = n1726 ;
  assign y22 = n1729 ;
  assign y23 = n1732 ;
  assign y24 = n1735 ;
  assign y25 = n1738 ;
  assign y26 = n1741 ;
  assign y27 = n1744 ;
  assign y28 = n1747 ;
  assign y29 = n1750 ;
  assign y30 = n1753 ;
  assign y31 = n1756 ;
  assign y32 = n1759 ;
  assign y33 = n1762 ;
  assign y34 = n1765 ;
  assign y35 = n1768 ;
  assign y36 = n1771 ;
  assign y37 = n1774 ;
  assign y38 = n1777 ;
  assign y39 = n1780 ;
  assign y40 = n1783 ;
  assign y41 = n1786 ;
  assign y42 = n1789 ;
  assign y43 = n1792 ;
  assign y44 = n1795 ;
  assign y45 = n1798 ;
  assign y46 = n1801 ;
  assign y47 = n1804 ;
  assign y48 = n1807 ;
  assign y49 = n1810 ;
  assign y50 = n1813 ;
  assign y51 = n1816 ;
  assign y52 = n1819 ;
  assign y53 = n1822 ;
  assign y54 = n1825 ;
  assign y55 = n1828 ;
  assign y56 = n1831 ;
  assign y57 = n1834 ;
  assign y58 = n1837 ;
  assign y59 = n1840 ;
  assign y60 = n1843 ;
  assign y61 = n1846 ;
  assign y62 = n1849 ;
  assign y63 = n1852 ;
  assign y64 = n1855 ;
  assign y65 = n1858 ;
  assign y66 = n1861 ;
  assign y67 = n1864 ;
  assign y68 = n1867 ;
  assign y69 = n1870 ;
  assign y70 = n1873 ;
  assign y71 = n1876 ;
  assign y72 = n1879 ;
  assign y73 = n1882 ;
  assign y74 = n1885 ;
  assign y75 = n1888 ;
  assign y76 = n1891 ;
  assign y77 = n1894 ;
  assign y78 = n1897 ;
  assign y79 = n1900 ;
  assign y80 = n1903 ;
  assign y81 = n1906 ;
  assign y82 = n1909 ;
  assign y83 = n1912 ;
  assign y84 = n1915 ;
  assign y85 = n1918 ;
  assign y86 = n1921 ;
  assign y87 = n1924 ;
  assign y88 = n1927 ;
  assign y89 = n1930 ;
  assign y90 = n1933 ;
  assign y91 = n1936 ;
  assign y92 = n1939 ;
  assign y93 = n1942 ;
  assign y94 = n1945 ;
  assign y95 = n1948 ;
  assign y96 = n1951 ;
  assign y97 = n1954 ;
  assign y98 = n1957 ;
  assign y99 = n1960 ;
  assign y100 = n1963 ;
  assign y101 = n1966 ;
  assign y102 = n1969 ;
  assign y103 = n1972 ;
  assign y104 = n1975 ;
  assign y105 = n1978 ;
  assign y106 = n1981 ;
  assign y107 = n1984 ;
  assign y108 = n1987 ;
  assign y109 = n1990 ;
  assign y110 = n1993 ;
  assign y111 = n1996 ;
  assign y112 = n1999 ;
  assign y113 = n2002 ;
  assign y114 = n2005 ;
  assign y115 = n2008 ;
  assign y116 = n2011 ;
  assign y117 = n2014 ;
  assign y118 = n2017 ;
  assign y119 = n2020 ;
  assign y120 = n2023 ;
  assign y121 = n2026 ;
  assign y122 = n2029 ;
  assign y123 = n2032 ;
  assign y124 = n2035 ;
  assign y125 = n2038 ;
  assign y126 = n2041 ;
  assign y127 = n2042 ;
  assign y128 = ~n2045 ;
  assign y129 = ~n1660 ;
endmodule
