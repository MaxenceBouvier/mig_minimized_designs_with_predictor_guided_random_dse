module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 ;
  assign n65 = ~x0 & x1 ;
  assign n66 = ~x1 & x2 ;
  assign n67 = x1 & ~x2 ;
  assign n68 = ( x0 & n66 ) | ( x0 & n67 ) | ( n66 & n67 ) ;
  assign n69 = x0 & x3 ;
  assign n70 = x2 & n69 ;
  assign n71 = x2 & ~n65 ;
  assign n72 = ~x2 & n69 ;
  assign n73 = ( ~n70 & n71 ) | ( ~n70 & n72 ) | ( n71 & n72 ) ;
  assign n74 = x2 & x3 ;
  assign n75 = ~x0 & n74 ;
  assign n76 = x0 & x4 ;
  assign n77 = ( x1 & x2 ) | ( x1 & x3 ) | ( x2 & x3 ) ;
  assign n78 = ~n76 & n77 ;
  assign n79 = n76 & ~n77 ;
  assign n80 = ( ~n75 & n78 ) | ( ~n75 & n79 ) | ( n78 & n79 ) ;
  assign n81 = x2 & n76 ;
  assign n82 = ( x3 & ~n66 ) | ( x3 & n81 ) | ( ~n66 & n81 ) ;
  assign n83 = x0 & x5 ;
  assign n84 = x1 & x4 ;
  assign n85 = ~n69 & n84 ;
  assign n86 = ( n82 & n83 ) | ( n82 & n85 ) | ( n83 & n85 ) ;
  assign n87 = ( ~n82 & n83 ) | ( ~n82 & n85 ) | ( n83 & n85 ) ;
  assign n88 = ( n82 & ~n86 ) | ( n82 & n87 ) | ( ~n86 & n87 ) ;
  assign n89 = x3 & x4 ;
  assign n90 = ( x2 & x4 ) | ( x2 & n74 ) | ( x4 & n74 ) ;
  assign n91 = ~n89 & n90 ;
  assign n92 = x1 & x5 ;
  assign n93 = x0 & x6 ;
  assign n94 = ( n91 & n92 ) | ( n91 & n93 ) | ( n92 & n93 ) ;
  assign n95 = ( ~n91 & n92 ) | ( ~n91 & n93 ) | ( n92 & n93 ) ;
  assign n96 = ( n91 & ~n94 ) | ( n91 & n95 ) | ( ~n94 & n95 ) ;
  assign n97 = x3 & n76 ;
  assign n98 = n92 & n97 ;
  assign n99 = n96 & n98 ;
  assign n100 = ( n82 & n83 ) | ( n82 & n84 ) | ( n83 & n84 ) ;
  assign n101 = ( n96 & ~n98 ) | ( n96 & n100 ) | ( ~n98 & n100 ) ;
  assign n102 = n96 & n100 ;
  assign n103 = ( n99 & n101 ) | ( n99 & ~n102 ) | ( n101 & ~n102 ) ;
  assign n104 = x2 & x5 ;
  assign n105 = ~x6 & n84 ;
  assign n106 = n104 & n105 ;
  assign n107 = ( n74 & n93 ) | ( n74 & ~n96 ) | ( n93 & ~n96 ) ;
  assign n108 = x1 & x6 ;
  assign n109 = x4 & ~n108 ;
  assign n110 = x4 & ~n104 ;
  assign n111 = x4 | n108 ;
  assign n112 = ( n109 & ~n110 ) | ( n109 & n111 ) | ( ~n110 & n111 ) ;
  assign n113 = ( n106 & n107 ) | ( n106 & n112 ) | ( n107 & n112 ) ;
  assign n114 = n107 | n112 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = x0 & x7 ;
  assign n117 = ( n89 & ~n104 ) | ( n89 & n116 ) | ( ~n104 & n116 ) ;
  assign n118 = ( n89 & n104 ) | ( n89 & n116 ) | ( n104 & n116 ) ;
  assign n119 = ( n104 & n117 ) | ( n104 & ~n118 ) | ( n117 & ~n118 ) ;
  assign n120 = ( n98 & n100 ) | ( n98 & n102 ) | ( n100 & n102 ) ;
  assign n121 = ( n115 & n119 ) | ( n115 & n120 ) | ( n119 & n120 ) ;
  assign n122 = ( ~n115 & n119 ) | ( ~n115 & n120 ) | ( n119 & n120 ) ;
  assign n123 = ( n115 & ~n121 ) | ( n115 & n122 ) | ( ~n121 & n122 ) ;
  assign n124 = ( x2 & ~x6 ) | ( x2 & n84 ) | ( ~x6 & n84 ) ;
  assign n125 = x0 & x8 ;
  assign n126 = x2 | n84 ;
  assign n127 = ( ~n124 & n125 ) | ( ~n124 & n126 ) | ( n125 & n126 ) ;
  assign n128 = ( n124 & n125 ) | ( n124 & n126 ) | ( n125 & n126 ) ;
  assign n129 = ( n124 & n127 ) | ( n124 & ~n128 ) | ( n127 & ~n128 ) ;
  assign n130 = x1 & x7 ;
  assign n131 = x3 & x5 ;
  assign n132 = n130 | n131 ;
  assign n133 = x3 & x7 ;
  assign n134 = n92 & n133 ;
  assign n135 = n132 & ~n134 ;
  assign n136 = ( n118 & ~n129 ) | ( n118 & n135 ) | ( ~n129 & n135 ) ;
  assign n137 = ( n118 & n129 ) | ( n118 & n135 ) | ( n129 & n135 ) ;
  assign n138 = ( n129 & n136 ) | ( n129 & ~n137 ) | ( n136 & ~n137 ) ;
  assign n139 = ( ~n113 & n121 ) | ( ~n113 & n138 ) | ( n121 & n138 ) ;
  assign n140 = ( n113 & n121 ) | ( n113 & n138 ) | ( n121 & n138 ) ;
  assign n141 = ( n113 & n139 ) | ( n113 & ~n140 ) | ( n139 & ~n140 ) ;
  assign n142 = ( x2 & n84 ) | ( x2 & n125 ) | ( n84 & n125 ) ;
  assign n143 = x6 & n142 ;
  assign n144 = x0 & x9 ;
  assign n145 = x1 & x8 ;
  assign n146 = x5 & ~n134 ;
  assign n147 = ( ~n144 & n145 ) | ( ~n144 & n146 ) | ( n145 & n146 ) ;
  assign n148 = ( n144 & n145 ) | ( n144 & n146 ) | ( n145 & n146 ) ;
  assign n149 = ( n144 & n147 ) | ( n144 & ~n148 ) | ( n147 & ~n148 ) ;
  assign n150 = x4 & x5 ;
  assign n151 = x3 & x6 ;
  assign n152 = x2 & x7 ;
  assign n153 = ( ~n150 & n151 ) | ( ~n150 & n152 ) | ( n151 & n152 ) ;
  assign n154 = ( n150 & n151 ) | ( n150 & n152 ) | ( n151 & n152 ) ;
  assign n155 = ( n150 & n153 ) | ( n150 & ~n154 ) | ( n153 & ~n154 ) ;
  assign n156 = ( ~n143 & n149 ) | ( ~n143 & n155 ) | ( n149 & n155 ) ;
  assign n157 = ( n143 & n149 ) | ( n143 & n155 ) | ( n149 & n155 ) ;
  assign n158 = ( n143 & n156 ) | ( n143 & ~n157 ) | ( n156 & ~n157 ) ;
  assign n159 = ( n137 & ~n140 ) | ( n137 & n158 ) | ( ~n140 & n158 ) ;
  assign n160 = ( n137 & n140 ) | ( n137 & n158 ) | ( n140 & n158 ) ;
  assign n161 = ( n140 & n159 ) | ( n140 & ~n160 ) | ( n159 & ~n160 ) ;
  assign n162 = ( n134 & n144 ) | ( n134 & ~n149 ) | ( n144 & ~n149 ) ;
  assign n163 = x0 & x10 ;
  assign n164 = x2 & x8 ;
  assign n165 = ( ~n133 & n163 ) | ( ~n133 & n164 ) | ( n163 & n164 ) ;
  assign n166 = ( n133 & n163 ) | ( n133 & n164 ) | ( n163 & n164 ) ;
  assign n167 = ( n133 & n165 ) | ( n133 & ~n166 ) | ( n165 & ~n166 ) ;
  assign n168 = x8 & n92 ;
  assign n169 = x1 & x9 ;
  assign n170 = x4 & x6 ;
  assign n171 = n169 | n170 ;
  assign n172 = x6 & x9 ;
  assign n173 = n84 & n172 ;
  assign n174 = n171 & ~n173 ;
  assign n175 = ( n154 & ~n168 ) | ( n154 & n174 ) | ( ~n168 & n174 ) ;
  assign n176 = ( n154 & n168 ) | ( n154 & n174 ) | ( n168 & n174 ) ;
  assign n177 = ( n168 & n175 ) | ( n168 & ~n176 ) | ( n175 & ~n176 ) ;
  assign n178 = ( n162 & n167 ) | ( n162 & n177 ) | ( n167 & n177 ) ;
  assign n179 = ( ~n162 & n167 ) | ( ~n162 & n177 ) | ( n167 & n177 ) ;
  assign n180 = ( n162 & ~n178 ) | ( n162 & n179 ) | ( ~n178 & n179 ) ;
  assign n181 = ( n157 & n160 ) | ( n157 & n180 ) | ( n160 & n180 ) ;
  assign n182 = ( n157 & ~n160 ) | ( n157 & n180 ) | ( ~n160 & n180 ) ;
  assign n183 = ( n160 & ~n181 ) | ( n160 & n182 ) | ( ~n181 & n182 ) ;
  assign n184 = x3 & x8 ;
  assign n185 = x9 & ~n184 ;
  assign n186 = ( x2 & n173 ) | ( x2 & n185 ) | ( n173 & n185 ) ;
  assign n187 = x8 & x9 ;
  assign n188 = x3 & n187 ;
  assign n189 = ( x2 & n173 ) | ( x2 & n188 ) | ( n173 & n188 ) ;
  assign n190 = ( n184 & n186 ) | ( n184 & ~n189 ) | ( n186 & ~n189 ) ;
  assign n191 = ~x1 & x6 ;
  assign n192 = ( x1 & x6 ) | ( x1 & x10 ) | ( x6 & x10 ) ;
  assign n193 = x6 & x10 ;
  assign n194 = ( n191 & n192 ) | ( n191 & ~n193 ) | ( n192 & ~n193 ) ;
  assign n195 = ( n166 & ~n190 ) | ( n166 & n194 ) | ( ~n190 & n194 ) ;
  assign n196 = ( n166 & n190 ) | ( n166 & n194 ) | ( n190 & n194 ) ;
  assign n197 = ( n190 & n195 ) | ( n190 & ~n196 ) | ( n195 & ~n196 ) ;
  assign n198 = x4 & x7 ;
  assign n199 = x0 & x11 ;
  assign n200 = x5 & x6 ;
  assign n201 = ( ~n198 & n199 ) | ( ~n198 & n200 ) | ( n199 & n200 ) ;
  assign n202 = ( n198 & n199 ) | ( n198 & n200 ) | ( n199 & n200 ) ;
  assign n203 = ( n198 & n201 ) | ( n198 & ~n202 ) | ( n201 & ~n202 ) ;
  assign n204 = ( n176 & ~n197 ) | ( n176 & n203 ) | ( ~n197 & n203 ) ;
  assign n205 = ( n176 & n197 ) | ( n176 & n203 ) | ( n197 & n203 ) ;
  assign n206 = ( n197 & n204 ) | ( n197 & ~n205 ) | ( n204 & ~n205 ) ;
  assign n207 = ( n178 & ~n181 ) | ( n178 & n206 ) | ( ~n181 & n206 ) ;
  assign n208 = ( n178 & n181 ) | ( n178 & n206 ) | ( n181 & n206 ) ;
  assign n209 = ( n181 & n207 ) | ( n181 & ~n208 ) | ( n207 & ~n208 ) ;
  assign n210 = x2 & x10 ;
  assign n211 = x0 & x12 ;
  assign n212 = x3 & x9 ;
  assign n213 = ( ~n210 & n211 ) | ( ~n210 & n212 ) | ( n211 & n212 ) ;
  assign n214 = ( n210 & n211 ) | ( n210 & n212 ) | ( n211 & n212 ) ;
  assign n215 = ( n210 & n213 ) | ( n210 & ~n214 ) | ( n213 & ~n214 ) ;
  assign n216 = ( n189 & n202 ) | ( n189 & n215 ) | ( n202 & n215 ) ;
  assign n217 = ( ~n189 & n202 ) | ( ~n189 & n215 ) | ( n202 & n215 ) ;
  assign n218 = ( n189 & ~n216 ) | ( n189 & n217 ) | ( ~n216 & n217 ) ;
  assign n219 = x7 & x11 ;
  assign n220 = n92 & n219 ;
  assign n221 = ( ~x1 & x11 ) | ( ~x1 & n220 ) | ( x11 & n220 ) ;
  assign n222 = x7 & ~n220 ;
  assign n223 = x5 & n222 ;
  assign n224 = ( x11 & ~n221 ) | ( x11 & n223 ) | ( ~n221 & n223 ) ;
  assign n225 = x10 & n108 ;
  assign n226 = x4 & x8 ;
  assign n227 = ( n224 & n225 ) | ( n224 & n226 ) | ( n225 & n226 ) ;
  assign n228 = ( ~n224 & n225 ) | ( ~n224 & n226 ) | ( n225 & n226 ) ;
  assign n229 = ( n224 & ~n227 ) | ( n224 & n228 ) | ( ~n227 & n228 ) ;
  assign n230 = ( n196 & n218 ) | ( n196 & n229 ) | ( n218 & n229 ) ;
  assign n231 = ( ~n196 & n218 ) | ( ~n196 & n229 ) | ( n218 & n229 ) ;
  assign n232 = ( n196 & ~n230 ) | ( n196 & n231 ) | ( ~n230 & n231 ) ;
  assign n233 = ( n205 & n208 ) | ( n205 & n232 ) | ( n208 & n232 ) ;
  assign n234 = ( n205 & ~n208 ) | ( n205 & n232 ) | ( ~n208 & n232 ) ;
  assign n235 = ( n208 & ~n233 ) | ( n208 & n234 ) | ( ~n233 & n234 ) ;
  assign n236 = x6 & x7 ;
  assign n237 = x2 & x11 ;
  assign n238 = x5 & x8 ;
  assign n239 = ( ~n236 & n237 ) | ( ~n236 & n238 ) | ( n237 & n238 ) ;
  assign n240 = ( n236 & n237 ) | ( n236 & n238 ) | ( n237 & n238 ) ;
  assign n241 = ( n236 & n239 ) | ( n236 & ~n240 ) | ( n239 & ~n240 ) ;
  assign n242 = x0 & x13 ;
  assign n243 = x3 & x10 ;
  assign n244 = x4 & x9 ;
  assign n245 = ( ~n242 & n243 ) | ( ~n242 & n244 ) | ( n243 & n244 ) ;
  assign n246 = ( n242 & n243 ) | ( n242 & n244 ) | ( n243 & n244 ) ;
  assign n247 = ( n242 & n245 ) | ( n242 & ~n246 ) | ( n245 & ~n246 ) ;
  assign n248 = ( ~n227 & n241 ) | ( ~n227 & n247 ) | ( n241 & n247 ) ;
  assign n249 = ( n227 & n241 ) | ( n227 & n247 ) | ( n241 & n247 ) ;
  assign n250 = ( n227 & n248 ) | ( n227 & ~n249 ) | ( n248 & ~n249 ) ;
  assign n251 = x1 & x12 ;
  assign n252 = ( n214 & ~n222 ) | ( n214 & n251 ) | ( ~n222 & n251 ) ;
  assign n253 = ( ~n214 & n222 ) | ( ~n214 & n251 ) | ( n222 & n251 ) ;
  assign n254 = ( ~n251 & n252 ) | ( ~n251 & n253 ) | ( n252 & n253 ) ;
  assign n255 = ( n216 & ~n230 ) | ( n216 & n254 ) | ( ~n230 & n254 ) ;
  assign n256 = ( n216 & n230 ) | ( n216 & n254 ) | ( n230 & n254 ) ;
  assign n257 = ( n230 & n255 ) | ( n230 & ~n256 ) | ( n255 & ~n256 ) ;
  assign n258 = ( n233 & ~n250 ) | ( n233 & n257 ) | ( ~n250 & n257 ) ;
  assign n259 = ( n233 & n250 ) | ( n233 & n257 ) | ( n250 & n257 ) ;
  assign n260 = ( n250 & n258 ) | ( n250 & ~n259 ) | ( n258 & ~n259 ) ;
  assign n261 = ( n214 & n220 ) | ( n214 & ~n254 ) | ( n220 & ~n254 ) ;
  assign n262 = x7 & n251 ;
  assign n263 = x4 & x10 ;
  assign n264 = x5 & x9 ;
  assign n265 = ( ~n262 & n263 ) | ( ~n262 & n264 ) | ( n263 & n264 ) ;
  assign n266 = ( n262 & n263 ) | ( n262 & n264 ) | ( n263 & n264 ) ;
  assign n267 = ( n262 & n265 ) | ( n262 & ~n266 ) | ( n265 & ~n266 ) ;
  assign n268 = x0 & x14 ;
  assign n269 = x2 & x12 ;
  assign n270 = x3 & x11 ;
  assign n271 = ( ~n268 & n269 ) | ( ~n268 & n270 ) | ( n269 & n270 ) ;
  assign n272 = ( n268 & n269 ) | ( n268 & n270 ) | ( n269 & n270 ) ;
  assign n273 = ( n268 & n271 ) | ( n268 & ~n272 ) | ( n271 & ~n272 ) ;
  assign n274 = ( ~n261 & n267 ) | ( ~n261 & n273 ) | ( n267 & n273 ) ;
  assign n275 = ( n261 & n267 ) | ( n261 & n273 ) | ( n267 & n273 ) ;
  assign n276 = ( n261 & n274 ) | ( n261 & ~n275 ) | ( n274 & ~n275 ) ;
  assign n277 = x6 & x8 ;
  assign n278 = x1 & x13 ;
  assign n279 = n277 | n278 ;
  assign n280 = x8 & x13 ;
  assign n281 = n108 & n280 ;
  assign n282 = n279 & ~n281 ;
  assign n283 = ( ~n240 & n246 ) | ( ~n240 & n282 ) | ( n246 & n282 ) ;
  assign n284 = ( n240 & n246 ) | ( n240 & n282 ) | ( n246 & n282 ) ;
  assign n285 = ( n240 & n283 ) | ( n240 & ~n284 ) | ( n283 & ~n284 ) ;
  assign n286 = ( n249 & ~n276 ) | ( n249 & n285 ) | ( ~n276 & n285 ) ;
  assign n287 = ( n249 & n276 ) | ( n249 & n285 ) | ( n276 & n285 ) ;
  assign n288 = ( n276 & n286 ) | ( n276 & ~n287 ) | ( n286 & ~n287 ) ;
  assign n289 = ( n256 & n259 ) | ( n256 & n288 ) | ( n259 & n288 ) ;
  assign n290 = ( n256 & ~n259 ) | ( n256 & n288 ) | ( ~n259 & n288 ) ;
  assign n291 = ( n259 & ~n289 ) | ( n259 & n290 ) | ( ~n289 & n290 ) ;
  assign n292 = x8 & ~n281 ;
  assign n293 = x4 & x11 ;
  assign n294 = x1 & x14 ;
  assign n295 = ( ~n292 & n293 ) | ( ~n292 & n294 ) | ( n293 & n294 ) ;
  assign n296 = ( n292 & n293 ) | ( n292 & n294 ) | ( n293 & n294 ) ;
  assign n297 = ( n292 & n295 ) | ( n292 & ~n296 ) | ( n295 & ~n296 ) ;
  assign n298 = x7 & x8 ;
  assign n299 = x2 & x13 ;
  assign n300 = ( ~n172 & n298 ) | ( ~n172 & n299 ) | ( n298 & n299 ) ;
  assign n301 = ( n172 & n298 ) | ( n172 & n299 ) | ( n298 & n299 ) ;
  assign n302 = ( n172 & n300 ) | ( n172 & ~n301 ) | ( n300 & ~n301 ) ;
  assign n303 = ( n284 & ~n297 ) | ( n284 & n302 ) | ( ~n297 & n302 ) ;
  assign n304 = ( n284 & n297 ) | ( n284 & n302 ) | ( n297 & n302 ) ;
  assign n305 = ( n297 & n303 ) | ( n297 & ~n304 ) | ( n303 & ~n304 ) ;
  assign n306 = x3 & x12 ;
  assign n307 = x5 & x10 ;
  assign n308 = x0 & x15 ;
  assign n309 = ( ~n306 & n307 ) | ( ~n306 & n308 ) | ( n307 & n308 ) ;
  assign n310 = ( n306 & n307 ) | ( n306 & n308 ) | ( n307 & n308 ) ;
  assign n311 = ( n306 & n309 ) | ( n306 & ~n310 ) | ( n309 & ~n310 ) ;
  assign n312 = ( ~n266 & n272 ) | ( ~n266 & n311 ) | ( n272 & n311 ) ;
  assign n313 = ( n266 & n272 ) | ( n266 & n311 ) | ( n272 & n311 ) ;
  assign n314 = ( n266 & n312 ) | ( n266 & ~n313 ) | ( n312 & ~n313 ) ;
  assign n315 = ( ~n275 & n305 ) | ( ~n275 & n314 ) | ( n305 & n314 ) ;
  assign n316 = ( n275 & n305 ) | ( n275 & n314 ) | ( n305 & n314 ) ;
  assign n317 = ( n275 & n315 ) | ( n275 & ~n316 ) | ( n315 & ~n316 ) ;
  assign n318 = ( n287 & n289 ) | ( n287 & n317 ) | ( n289 & n317 ) ;
  assign n319 = ( n287 & ~n289 ) | ( n287 & n317 ) | ( ~n289 & n317 ) ;
  assign n320 = ( n289 & ~n318 ) | ( n289 & n319 ) | ( ~n318 & n319 ) ;
  assign n321 = x8 & n294 ;
  assign n322 = ( n281 & n296 ) | ( n281 & ~n321 ) | ( n296 & ~n321 ) ;
  assign n323 = x5 & x11 ;
  assign n324 = x0 & x16 ;
  assign n325 = ( ~n193 & n323 ) | ( ~n193 & n324 ) | ( n323 & n324 ) ;
  assign n326 = ( n193 & n323 ) | ( n193 & n324 ) | ( n323 & n324 ) ;
  assign n327 = ( n193 & n325 ) | ( n193 & ~n326 ) | ( n325 & ~n326 ) ;
  assign n328 = ( n310 & ~n322 ) | ( n310 & n327 ) | ( ~n322 & n327 ) ;
  assign n329 = ( n310 & n322 ) | ( n310 & n327 ) | ( n322 & n327 ) ;
  assign n330 = ( n322 & n328 ) | ( n322 & ~n329 ) | ( n328 & ~n329 ) ;
  assign n331 = x1 & x15 ;
  assign n332 = x7 & x9 ;
  assign n333 = n331 | n332 ;
  assign n334 = x9 & x15 ;
  assign n335 = n130 & n334 ;
  assign n336 = n333 & ~n335 ;
  assign n337 = ( n301 & n321 ) | ( n301 & n336 ) | ( n321 & n336 ) ;
  assign n338 = ( n301 & ~n321 ) | ( n301 & n336 ) | ( ~n321 & n336 ) ;
  assign n339 = ( n321 & ~n337 ) | ( n321 & n338 ) | ( ~n337 & n338 ) ;
  assign n340 = x4 & x12 ;
  assign n341 = x3 & x13 ;
  assign n342 = x2 & x14 ;
  assign n343 = ( ~n340 & n341 ) | ( ~n340 & n342 ) | ( n341 & n342 ) ;
  assign n344 = ( n340 & n341 ) | ( n340 & n342 ) | ( n341 & n342 ) ;
  assign n345 = ( n340 & n343 ) | ( n340 & ~n344 ) | ( n343 & ~n344 ) ;
  assign n346 = ( n313 & n339 ) | ( n313 & n345 ) | ( n339 & n345 ) ;
  assign n347 = ( ~n313 & n339 ) | ( ~n313 & n345 ) | ( n339 & n345 ) ;
  assign n348 = ( n313 & ~n346 ) | ( n313 & n347 ) | ( ~n346 & n347 ) ;
  assign n349 = ( n304 & n330 ) | ( n304 & n348 ) | ( n330 & n348 ) ;
  assign n350 = ( n304 & ~n330 ) | ( n304 & n348 ) | ( ~n330 & n348 ) ;
  assign n351 = ( n330 & ~n349 ) | ( n330 & n350 ) | ( ~n349 & n350 ) ;
  assign n352 = ( n316 & n318 ) | ( n316 & n351 ) | ( n318 & n351 ) ;
  assign n353 = ( n316 & ~n318 ) | ( n316 & n351 ) | ( ~n318 & n351 ) ;
  assign n354 = ( n318 & ~n352 ) | ( n318 & n353 ) | ( ~n352 & n353 ) ;
  assign n355 = x1 & x16 ;
  assign n356 = x9 | n355 ;
  assign n357 = x16 & n169 ;
  assign n358 = n356 & ~n357 ;
  assign n359 = ( n326 & ~n344 ) | ( n326 & n358 ) | ( ~n344 & n358 ) ;
  assign n360 = ( n326 & n344 ) | ( n326 & n358 ) | ( n344 & n358 ) ;
  assign n361 = ( n344 & n359 ) | ( n344 & ~n360 ) | ( n359 & ~n360 ) ;
  assign n362 = ( ~n329 & n337 ) | ( ~n329 & n361 ) | ( n337 & n361 ) ;
  assign n363 = ( n329 & n337 ) | ( n329 & n361 ) | ( n337 & n361 ) ;
  assign n364 = ( n329 & n362 ) | ( n329 & ~n363 ) | ( n362 & ~n363 ) ;
  assign n365 = x0 & x17 ;
  assign n366 = x5 & x12 ;
  assign n367 = ( ~n335 & n365 ) | ( ~n335 & n366 ) | ( n365 & n366 ) ;
  assign n368 = ( n335 & n365 ) | ( n335 & n366 ) | ( n365 & n366 ) ;
  assign n369 = ( n335 & n367 ) | ( n335 & ~n368 ) | ( n367 & ~n368 ) ;
  assign n370 = x2 & x15 ;
  assign n371 = x6 & x11 ;
  assign n372 = x4 & x13 ;
  assign n373 = ( ~n370 & n371 ) | ( ~n370 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( n370 & n371 ) | ( n370 & n372 ) | ( n371 & n372 ) ;
  assign n375 = ( n370 & n373 ) | ( n370 & ~n374 ) | ( n373 & ~n374 ) ;
  assign n376 = x3 & x14 ;
  assign n377 = x7 & x10 ;
  assign n378 = ( ~n187 & n376 ) | ( ~n187 & n377 ) | ( n376 & n377 ) ;
  assign n379 = ( n187 & n376 ) | ( n187 & n377 ) | ( n376 & n377 ) ;
  assign n380 = ( n187 & n378 ) | ( n187 & ~n379 ) | ( n378 & ~n379 ) ;
  assign n381 = ( ~n369 & n375 ) | ( ~n369 & n380 ) | ( n375 & n380 ) ;
  assign n382 = ( n369 & n375 ) | ( n369 & n380 ) | ( n375 & n380 ) ;
  assign n383 = ( n369 & n381 ) | ( n369 & ~n382 ) | ( n381 & ~n382 ) ;
  assign n384 = ( n346 & n364 ) | ( n346 & n383 ) | ( n364 & n383 ) ;
  assign n385 = ( n346 & ~n364 ) | ( n346 & n383 ) | ( ~n364 & n383 ) ;
  assign n386 = ( n364 & ~n384 ) | ( n364 & n385 ) | ( ~n384 & n385 ) ;
  assign n387 = ( n349 & ~n352 ) | ( n349 & n386 ) | ( ~n352 & n386 ) ;
  assign n388 = ( n349 & n352 ) | ( n349 & n386 ) | ( n352 & n386 ) ;
  assign n389 = ( n352 & n387 ) | ( n352 & ~n388 ) | ( n387 & ~n388 ) ;
  assign n390 = ( ~n368 & n374 ) | ( ~n368 & n379 ) | ( n374 & n379 ) ;
  assign n391 = ( n368 & n374 ) | ( n368 & n379 ) | ( n374 & n379 ) ;
  assign n392 = ( n368 & n390 ) | ( n368 & ~n391 ) | ( n390 & ~n391 ) ;
  assign n393 = ( n360 & n382 ) | ( n360 & n392 ) | ( n382 & n392 ) ;
  assign n394 = ( n360 & n382 ) | ( n360 & ~n392 ) | ( n382 & ~n392 ) ;
  assign n395 = ( n392 & ~n393 ) | ( n392 & n394 ) | ( ~n393 & n394 ) ;
  assign n396 = x1 & x17 ;
  assign n397 = x8 & x10 ;
  assign n398 = n396 | n397 ;
  assign n399 = x10 & x17 ;
  assign n400 = n145 & n399 ;
  assign n401 = n398 & ~n400 ;
  assign n402 = x6 & x12 ;
  assign n403 = ( n357 & n401 ) | ( n357 & n402 ) | ( n401 & n402 ) ;
  assign n404 = ( n357 & ~n401 ) | ( n357 & n402 ) | ( ~n401 & n402 ) ;
  assign n405 = ( n401 & ~n403 ) | ( n401 & n404 ) | ( ~n403 & n404 ) ;
  assign n406 = x2 & x16 ;
  assign n407 = x4 & x14 ;
  assign n408 = x3 & x15 ;
  assign n409 = ( ~n406 & n407 ) | ( ~n406 & n408 ) | ( n407 & n408 ) ;
  assign n410 = ( n406 & n407 ) | ( n406 & n408 ) | ( n407 & n408 ) ;
  assign n411 = ( n406 & n409 ) | ( n406 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = x5 & x13 ;
  assign n413 = x0 & x18 ;
  assign n414 = ( ~n219 & n412 ) | ( ~n219 & n413 ) | ( n412 & n413 ) ;
  assign n415 = ( n219 & n412 ) | ( n219 & n413 ) | ( n412 & n413 ) ;
  assign n416 = ( n219 & n414 ) | ( n219 & ~n415 ) | ( n414 & ~n415 ) ;
  assign n417 = ( n405 & n411 ) | ( n405 & n416 ) | ( n411 & n416 ) ;
  assign n418 = ( ~n405 & n411 ) | ( ~n405 & n416 ) | ( n411 & n416 ) ;
  assign n419 = ( n405 & ~n417 ) | ( n405 & n418 ) | ( ~n417 & n418 ) ;
  assign n420 = ( ~n363 & n395 ) | ( ~n363 & n419 ) | ( n395 & n419 ) ;
  assign n421 = ( n363 & n395 ) | ( n363 & n419 ) | ( n395 & n419 ) ;
  assign n422 = ( n363 & n420 ) | ( n363 & ~n421 ) | ( n420 & ~n421 ) ;
  assign n423 = ( n384 & n388 ) | ( n384 & n422 ) | ( n388 & n422 ) ;
  assign n424 = ( n384 & ~n388 ) | ( n384 & n422 ) | ( ~n388 & n422 ) ;
  assign n425 = ( n388 & ~n423 ) | ( n388 & n424 ) | ( ~n423 & n424 ) ;
  assign n426 = x9 & x10 ;
  assign n427 = x3 & x16 ;
  assign n428 = x8 & x11 ;
  assign n429 = ( ~n426 & n427 ) | ( ~n426 & n428 ) | ( n427 & n428 ) ;
  assign n430 = ( n426 & n427 ) | ( n426 & n428 ) | ( n427 & n428 ) ;
  assign n431 = ( n426 & n429 ) | ( n426 & ~n430 ) | ( n429 & ~n430 ) ;
  assign n432 = ( ~n403 & n415 ) | ( ~n403 & n431 ) | ( n415 & n431 ) ;
  assign n433 = ( n403 & n415 ) | ( n403 & n431 ) | ( n415 & n431 ) ;
  assign n434 = ( n403 & n432 ) | ( n403 & ~n433 ) | ( n432 & ~n433 ) ;
  assign n435 = ~x1 & x10 ;
  assign n436 = ( x1 & x10 ) | ( x1 & x18 ) | ( x10 & x18 ) ;
  assign n437 = x10 & x18 ;
  assign n438 = ( n435 & n436 ) | ( n435 & ~n437 ) | ( n436 & ~n437 ) ;
  assign n439 = ( n400 & n410 ) | ( n400 & n438 ) | ( n410 & n438 ) ;
  assign n440 = ( n400 & ~n410 ) | ( n400 & n438 ) | ( ~n410 & n438 ) ;
  assign n441 = ( n410 & ~n439 ) | ( n410 & n440 ) | ( ~n439 & n440 ) ;
  assign n442 = ( ~n417 & n434 ) | ( ~n417 & n441 ) | ( n434 & n441 ) ;
  assign n443 = ( n417 & n434 ) | ( n417 & n441 ) | ( n434 & n441 ) ;
  assign n444 = ( n417 & n442 ) | ( n417 & ~n443 ) | ( n442 & ~n443 ) ;
  assign n445 = x6 & x13 ;
  assign n446 = x5 & x14 ;
  assign n447 = x7 & x12 ;
  assign n448 = ( ~n445 & n446 ) | ( ~n445 & n447 ) | ( n446 & n447 ) ;
  assign n449 = ( n445 & n446 ) | ( n445 & n447 ) | ( n446 & n447 ) ;
  assign n450 = ( n445 & n448 ) | ( n445 & ~n449 ) | ( n448 & ~n449 ) ;
  assign n451 = x0 & x19 ;
  assign n452 = x4 & x15 ;
  assign n453 = x2 & x17 ;
  assign n454 = ( ~n451 & n452 ) | ( ~n451 & n453 ) | ( n452 & n453 ) ;
  assign n455 = ( n451 & n452 ) | ( n451 & n453 ) | ( n452 & n453 ) ;
  assign n456 = ( n451 & n454 ) | ( n451 & ~n455 ) | ( n454 & ~n455 ) ;
  assign n457 = ( ~n391 & n450 ) | ( ~n391 & n456 ) | ( n450 & n456 ) ;
  assign n458 = ( n391 & n450 ) | ( n391 & n456 ) | ( n450 & n456 ) ;
  assign n459 = ( n391 & n457 ) | ( n391 & ~n458 ) | ( n457 & ~n458 ) ;
  assign n460 = ( n393 & n444 ) | ( n393 & n459 ) | ( n444 & n459 ) ;
  assign n461 = ( n393 & ~n444 ) | ( n393 & n459 ) | ( ~n444 & n459 ) ;
  assign n462 = ( n444 & ~n460 ) | ( n444 & n461 ) | ( ~n460 & n461 ) ;
  assign n463 = ( n421 & ~n423 ) | ( n421 & n462 ) | ( ~n423 & n462 ) ;
  assign n464 = ( n421 & n423 ) | ( n421 & n462 ) | ( n423 & n462 ) ;
  assign n465 = ( n423 & n463 ) | ( n423 & ~n464 ) | ( n463 & ~n464 ) ;
  assign n466 = x1 & n437 ;
  assign n467 = x0 & x20 ;
  assign n468 = x7 & x13 ;
  assign n469 = ( ~n466 & n467 ) | ( ~n466 & n468 ) | ( n467 & n468 ) ;
  assign n470 = ( n466 & n467 ) | ( n466 & n468 ) | ( n467 & n468 ) ;
  assign n471 = ( n466 & n469 ) | ( n466 & ~n470 ) | ( n469 & ~n470 ) ;
  assign n472 = x8 & x12 ;
  assign n473 = x5 & x15 ;
  assign n474 = x6 & x14 ;
  assign n475 = ( ~n472 & n473 ) | ( ~n472 & n474 ) | ( n473 & n474 ) ;
  assign n476 = ( n472 & n473 ) | ( n472 & n474 ) | ( n473 & n474 ) ;
  assign n477 = ( n472 & n475 ) | ( n472 & ~n476 ) | ( n475 & ~n476 ) ;
  assign n478 = ( n449 & ~n471 ) | ( n449 & n477 ) | ( ~n471 & n477 ) ;
  assign n479 = ( n449 & n471 ) | ( n449 & n477 ) | ( n471 & n477 ) ;
  assign n480 = ( n471 & n478 ) | ( n471 & ~n479 ) | ( n478 & ~n479 ) ;
  assign n481 = x1 & x19 ;
  assign n482 = x9 & x11 ;
  assign n483 = n481 & n482 ;
  assign n484 = n481 | n482 ;
  assign n485 = ~n483 & n484 ;
  assign n486 = ( ~n430 & n455 ) | ( ~n430 & n485 ) | ( n455 & n485 ) ;
  assign n487 = ( n430 & n455 ) | ( n430 & n485 ) | ( n455 & n485 ) ;
  assign n488 = ( n430 & n486 ) | ( n430 & ~n487 ) | ( n486 & ~n487 ) ;
  assign n489 = ( ~n458 & n480 ) | ( ~n458 & n488 ) | ( n480 & n488 ) ;
  assign n490 = ( n458 & n480 ) | ( n458 & n488 ) | ( n480 & n488 ) ;
  assign n491 = ( n458 & n489 ) | ( n458 & ~n490 ) | ( n489 & ~n490 ) ;
  assign n492 = x2 & x18 ;
  assign n493 = x4 & x16 ;
  assign n494 = x3 & x17 ;
  assign n495 = ( ~n492 & n493 ) | ( ~n492 & n494 ) | ( n493 & n494 ) ;
  assign n496 = ( n492 & n493 ) | ( n492 & n494 ) | ( n493 & n494 ) ;
  assign n497 = ( n492 & n495 ) | ( n492 & ~n496 ) | ( n495 & ~n496 ) ;
  assign n498 = ( n433 & n439 ) | ( n433 & ~n497 ) | ( n439 & ~n497 ) ;
  assign n499 = ( n433 & n439 ) | ( n433 & n497 ) | ( n439 & n497 ) ;
  assign n500 = ( n497 & n498 ) | ( n497 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = ( n443 & n491 ) | ( n443 & n500 ) | ( n491 & n500 ) ;
  assign n502 = ( n443 & ~n491 ) | ( n443 & n500 ) | ( ~n491 & n500 ) ;
  assign n503 = ( n491 & ~n501 ) | ( n491 & n502 ) | ( ~n501 & n502 ) ;
  assign n504 = ( n460 & n464 ) | ( n460 & n503 ) | ( n464 & n503 ) ;
  assign n505 = ( n460 & ~n464 ) | ( n460 & n503 ) | ( ~n464 & n503 ) ;
  assign n506 = ( n464 & ~n504 ) | ( n464 & n505 ) | ( ~n504 & n505 ) ;
  assign n507 = ( ~n470 & n476 ) | ( ~n470 & n496 ) | ( n476 & n496 ) ;
  assign n508 = ( n470 & n476 ) | ( n470 & n496 ) | ( n476 & n496 ) ;
  assign n509 = ( n470 & n507 ) | ( n470 & ~n508 ) | ( n507 & ~n508 ) ;
  assign n510 = x3 & x18 ;
  assign n511 = x2 & x19 ;
  assign n512 = x5 & x16 ;
  assign n513 = ( ~n510 & n511 ) | ( ~n510 & n512 ) | ( n511 & n512 ) ;
  assign n514 = ( n510 & n511 ) | ( n510 & n512 ) | ( n511 & n512 ) ;
  assign n515 = ( n510 & n513 ) | ( n510 & ~n514 ) | ( n513 & ~n514 ) ;
  assign n516 = x7 & x14 ;
  assign n517 = x6 & x15 ;
  assign n518 = ( ~n280 & n516 ) | ( ~n280 & n517 ) | ( n516 & n517 ) ;
  assign n519 = ( n280 & n516 ) | ( n280 & n517 ) | ( n516 & n517 ) ;
  assign n520 = ( n280 & n518 ) | ( n280 & ~n519 ) | ( n518 & ~n519 ) ;
  assign n521 = x9 & x12 ;
  assign n522 = x10 & x11 ;
  assign n523 = x4 & x17 ;
  assign n524 = ( ~n521 & n522 ) | ( ~n521 & n523 ) | ( n522 & n523 ) ;
  assign n525 = ( n521 & n522 ) | ( n521 & n523 ) | ( n522 & n523 ) ;
  assign n526 = ( n521 & n524 ) | ( n521 & ~n525 ) | ( n524 & ~n525 ) ;
  assign n527 = ( ~n515 & n520 ) | ( ~n515 & n526 ) | ( n520 & n526 ) ;
  assign n528 = ( n515 & n520 ) | ( n515 & n526 ) | ( n520 & n526 ) ;
  assign n529 = ( n515 & n527 ) | ( n515 & ~n528 ) | ( n527 & ~n528 ) ;
  assign n530 = ( ~n499 & n509 ) | ( ~n499 & n529 ) | ( n509 & n529 ) ;
  assign n531 = ( n499 & n509 ) | ( n499 & n529 ) | ( n509 & n529 ) ;
  assign n532 = ( n499 & n530 ) | ( n499 & ~n531 ) | ( n530 & ~n531 ) ;
  assign n533 = x9 & x19 ;
  assign n534 = x1 & x20 ;
  assign n535 = x11 & n534 ;
  assign n536 = ~n533 & n535 ;
  assign n537 = x11 | n534 ;
  assign n538 = ~n536 & n537 ;
  assign n539 = x0 & x21 ;
  assign n540 = n538 | n539 ;
  assign n541 = ~x20 & n483 ;
  assign n542 = ( ~n538 & n539 ) | ( ~n538 & n541 ) | ( n539 & n541 ) ;
  assign n543 = n539 | n541 ;
  assign n544 = ( n540 & n542 ) | ( n540 & ~n543 ) | ( n542 & ~n543 ) ;
  assign n545 = ( ~n479 & n487 ) | ( ~n479 & n544 ) | ( n487 & n544 ) ;
  assign n546 = ( n479 & n487 ) | ( n479 & n544 ) | ( n487 & n544 ) ;
  assign n547 = ( n479 & n545 ) | ( n479 & ~n546 ) | ( n545 & ~n546 ) ;
  assign n548 = ( n490 & n532 ) | ( n490 & n547 ) | ( n532 & n547 ) ;
  assign n549 = ( n490 & ~n532 ) | ( n490 & n547 ) | ( ~n532 & n547 ) ;
  assign n550 = ( n532 & ~n548 ) | ( n532 & n549 ) | ( ~n548 & n549 ) ;
  assign n551 = ( n501 & ~n504 ) | ( n501 & n550 ) | ( ~n504 & n550 ) ;
  assign n552 = ( n501 & n504 ) | ( n501 & n550 ) | ( n504 & n550 ) ;
  assign n553 = ( n504 & n551 ) | ( n504 & ~n552 ) | ( n551 & ~n552 ) ;
  assign n554 = ( n538 & n541 ) | ( n538 & n543 ) | ( n541 & n543 ) ;
  assign n555 = ( n514 & n519 ) | ( n514 & ~n554 ) | ( n519 & ~n554 ) ;
  assign n556 = ( n514 & n519 ) | ( n514 & n554 ) | ( n519 & n554 ) ;
  assign n557 = ( n554 & n555 ) | ( n554 & ~n556 ) | ( n555 & ~n556 ) ;
  assign n558 = x3 & x19 ;
  assign n559 = x4 & x18 ;
  assign n560 = x5 & x17 ;
  assign n561 = ( ~n558 & n559 ) | ( ~n558 & n560 ) | ( n559 & n560 ) ;
  assign n562 = ( n558 & n559 ) | ( n558 & n560 ) | ( n559 & n560 ) ;
  assign n563 = ( n558 & n561 ) | ( n558 & ~n562 ) | ( n561 & ~n562 ) ;
  assign n564 = x0 & x22 ;
  assign n565 = x8 & x14 ;
  assign n566 = x7 & x15 ;
  assign n567 = ( ~n564 & n565 ) | ( ~n564 & n566 ) | ( n565 & n566 ) ;
  assign n568 = ( n564 & n565 ) | ( n564 & n566 ) | ( n565 & n566 ) ;
  assign n569 = ( n564 & n567 ) | ( n564 & ~n568 ) | ( n567 & ~n568 ) ;
  assign n570 = x6 & x16 ;
  assign n571 = x9 & x13 ;
  assign n572 = x2 & x20 ;
  assign n573 = ( ~n570 & n571 ) | ( ~n570 & n572 ) | ( n571 & n572 ) ;
  assign n574 = ( n570 & n571 ) | ( n570 & n572 ) | ( n571 & n572 ) ;
  assign n575 = ( n570 & n573 ) | ( n570 & ~n574 ) | ( n573 & ~n574 ) ;
  assign n576 = ( ~n563 & n569 ) | ( ~n563 & n575 ) | ( n569 & n575 ) ;
  assign n577 = ( n563 & n569 ) | ( n563 & n575 ) | ( n569 & n575 ) ;
  assign n578 = ( n563 & n576 ) | ( n563 & ~n577 ) | ( n576 & ~n577 ) ;
  assign n579 = ( n546 & n557 ) | ( n546 & n578 ) | ( n557 & n578 ) ;
  assign n580 = ( ~n546 & n557 ) | ( ~n546 & n578 ) | ( n557 & n578 ) ;
  assign n581 = ( n546 & ~n579 ) | ( n546 & n580 ) | ( ~n579 & n580 ) ;
  assign n582 = x1 & x21 ;
  assign n583 = x10 & x12 ;
  assign n584 = n582 | n583 ;
  assign n585 = x10 & x21 ;
  assign n586 = n251 & n585 ;
  assign n587 = n584 & ~n586 ;
  assign n588 = ( n525 & n535 ) | ( n525 & n587 ) | ( n535 & n587 ) ;
  assign n589 = ( n525 & ~n535 ) | ( n525 & n587 ) | ( ~n535 & n587 ) ;
  assign n590 = ( n535 & ~n588 ) | ( n535 & n589 ) | ( ~n588 & n589 ) ;
  assign n591 = ( n508 & n528 ) | ( n508 & n590 ) | ( n528 & n590 ) ;
  assign n592 = ( ~n508 & n528 ) | ( ~n508 & n590 ) | ( n528 & n590 ) ;
  assign n593 = ( n508 & ~n591 ) | ( n508 & n592 ) | ( ~n591 & n592 ) ;
  assign n594 = ( n531 & n581 ) | ( n531 & n593 ) | ( n581 & n593 ) ;
  assign n595 = ( ~n531 & n581 ) | ( ~n531 & n593 ) | ( n581 & n593 ) ;
  assign n596 = ( n531 & ~n594 ) | ( n531 & n595 ) | ( ~n594 & n595 ) ;
  assign n597 = ( n548 & n552 ) | ( n548 & n596 ) | ( n552 & n596 ) ;
  assign n598 = ( n548 & ~n552 ) | ( n548 & n596 ) | ( ~n552 & n596 ) ;
  assign n599 = ( n552 & ~n597 ) | ( n552 & n598 ) | ( ~n597 & n598 ) ;
  assign n600 = x1 & x22 ;
  assign n601 = x12 | n600 ;
  assign n602 = x22 & n251 ;
  assign n603 = n601 & ~n602 ;
  assign n604 = ( n562 & ~n574 ) | ( n562 & n603 ) | ( ~n574 & n603 ) ;
  assign n605 = ( n562 & n574 ) | ( n562 & n603 ) | ( n574 & n603 ) ;
  assign n606 = ( n574 & n604 ) | ( n574 & ~n605 ) | ( n604 & ~n605 ) ;
  assign n607 = ( ~n556 & n577 ) | ( ~n556 & n606 ) | ( n577 & n606 ) ;
  assign n608 = ( n556 & n577 ) | ( n556 & n606 ) | ( n577 & n606 ) ;
  assign n609 = ( n556 & n607 ) | ( n556 & ~n608 ) | ( n607 & ~n608 ) ;
  assign n610 = x2 & x21 ;
  assign n611 = x0 & x23 ;
  assign n612 = ( ~n586 & n610 ) | ( ~n586 & n611 ) | ( n610 & n611 ) ;
  assign n613 = ( n586 & n610 ) | ( n586 & n611 ) | ( n610 & n611 ) ;
  assign n614 = ( n586 & n612 ) | ( n586 & ~n613 ) | ( n612 & ~n613 ) ;
  assign n615 = x7 & x16 ;
  assign n616 = x9 & x14 ;
  assign n617 = x8 & x15 ;
  assign n618 = ( ~n615 & n616 ) | ( ~n615 & n617 ) | ( n616 & n617 ) ;
  assign n619 = ( n615 & n616 ) | ( n615 & n617 ) | ( n616 & n617 ) ;
  assign n620 = ( n615 & n618 ) | ( n615 & ~n619 ) | ( n618 & ~n619 ) ;
  assign n621 = ( n568 & ~n614 ) | ( n568 & n620 ) | ( ~n614 & n620 ) ;
  assign n622 = ( n568 & n614 ) | ( n568 & n620 ) | ( n614 & n620 ) ;
  assign n623 = ( n614 & n621 ) | ( n614 & ~n622 ) | ( n621 & ~n622 ) ;
  assign n624 = x3 & x20 ;
  assign n625 = x6 & x17 ;
  assign n626 = x5 & x18 ;
  assign n627 = ( ~n624 & n625 ) | ( ~n624 & n626 ) | ( n625 & n626 ) ;
  assign n628 = ( n624 & n625 ) | ( n624 & n626 ) | ( n625 & n626 ) ;
  assign n629 = ( n624 & n627 ) | ( n624 & ~n628 ) | ( n627 & ~n628 ) ;
  assign n630 = x11 & x12 ;
  assign n631 = x4 & x19 ;
  assign n632 = x10 & x13 ;
  assign n633 = ( ~n630 & n631 ) | ( ~n630 & n632 ) | ( n631 & n632 ) ;
  assign n634 = ( n630 & n631 ) | ( n630 & n632 ) | ( n631 & n632 ) ;
  assign n635 = ( n630 & n633 ) | ( n630 & ~n634 ) | ( n633 & ~n634 ) ;
  assign n636 = ( ~n588 & n629 ) | ( ~n588 & n635 ) | ( n629 & n635 ) ;
  assign n637 = ( n588 & n629 ) | ( n588 & n635 ) | ( n629 & n635 ) ;
  assign n638 = ( n588 & n636 ) | ( n588 & ~n637 ) | ( n636 & ~n637 ) ;
  assign n639 = ( n591 & n623 ) | ( n591 & n638 ) | ( n623 & n638 ) ;
  assign n640 = ( ~n591 & n623 ) | ( ~n591 & n638 ) | ( n623 & n638 ) ;
  assign n641 = ( n591 & ~n639 ) | ( n591 & n640 ) | ( ~n639 & n640 ) ;
  assign n642 = ( n579 & ~n609 ) | ( n579 & n641 ) | ( ~n609 & n641 ) ;
  assign n643 = ( n579 & n609 ) | ( n579 & n641 ) | ( n609 & n641 ) ;
  assign n644 = ( n609 & n642 ) | ( n609 & ~n643 ) | ( n642 & ~n643 ) ;
  assign n645 = ( n594 & n597 ) | ( n594 & n644 ) | ( n597 & n644 ) ;
  assign n646 = ( n594 & ~n597 ) | ( n594 & n644 ) | ( ~n597 & n644 ) ;
  assign n647 = ( n597 & ~n645 ) | ( n597 & n646 ) | ( ~n645 & n646 ) ;
  assign n648 = x1 & x23 ;
  assign n649 = x11 & x13 ;
  assign n650 = n648 & n649 ;
  assign n651 = n648 | n649 ;
  assign n652 = ~n650 & n651 ;
  assign n653 = x0 & x24 ;
  assign n654 = ( n602 & n652 ) | ( n602 & n653 ) | ( n652 & n653 ) ;
  assign n655 = ( n602 & ~n652 ) | ( n602 & n653 ) | ( ~n652 & n653 ) ;
  assign n656 = ( n652 & ~n654 ) | ( n652 & n655 ) | ( ~n654 & n655 ) ;
  assign n657 = x6 & x18 ;
  assign n658 = x7 & x17 ;
  assign n659 = x2 & x22 ;
  assign n660 = ( ~n657 & n658 ) | ( ~n657 & n659 ) | ( n658 & n659 ) ;
  assign n661 = ( n657 & n658 ) | ( n657 & n659 ) | ( n658 & n659 ) ;
  assign n662 = ( n657 & n660 ) | ( n657 & ~n661 ) | ( n660 & ~n661 ) ;
  assign n663 = ( n605 & n656 ) | ( n605 & n662 ) | ( n656 & n662 ) ;
  assign n664 = ( n605 & ~n656 ) | ( n605 & n662 ) | ( ~n656 & n662 ) ;
  assign n665 = ( n656 & ~n663 ) | ( n656 & n664 ) | ( ~n663 & n664 ) ;
  assign n666 = x8 & x16 ;
  assign n667 = x10 & x14 ;
  assign n668 = ( ~n334 & n666 ) | ( ~n334 & n667 ) | ( n666 & n667 ) ;
  assign n669 = ( n334 & n666 ) | ( n334 & n667 ) | ( n666 & n667 ) ;
  assign n670 = ( n334 & n668 ) | ( n334 & ~n669 ) | ( n668 & ~n669 ) ;
  assign n671 = x4 & x20 ;
  assign n672 = x3 & x21 ;
  assign n673 = x5 & x19 ;
  assign n674 = ( ~n671 & n672 ) | ( ~n671 & n673 ) | ( n672 & n673 ) ;
  assign n675 = ( n671 & n672 ) | ( n671 & n673 ) | ( n672 & n673 ) ;
  assign n676 = ( n671 & n674 ) | ( n671 & ~n675 ) | ( n674 & ~n675 ) ;
  assign n677 = ( ~n613 & n670 ) | ( ~n613 & n676 ) | ( n670 & n676 ) ;
  assign n678 = ( n613 & n670 ) | ( n613 & n676 ) | ( n670 & n676 ) ;
  assign n679 = ( n613 & n677 ) | ( n613 & ~n678 ) | ( n677 & ~n678 ) ;
  assign n680 = ( n608 & n665 ) | ( n608 & n679 ) | ( n665 & n679 ) ;
  assign n681 = ( n608 & ~n665 ) | ( n608 & n679 ) | ( ~n665 & n679 ) ;
  assign n682 = ( n665 & ~n680 ) | ( n665 & n681 ) | ( ~n680 & n681 ) ;
  assign n683 = ( ~n619 & n628 ) | ( ~n619 & n634 ) | ( n628 & n634 ) ;
  assign n684 = ( n619 & n628 ) | ( n619 & n634 ) | ( n628 & n634 ) ;
  assign n685 = ( n619 & n683 ) | ( n619 & ~n684 ) | ( n683 & ~n684 ) ;
  assign n686 = ( n622 & n637 ) | ( n622 & n685 ) | ( n637 & n685 ) ;
  assign n687 = ( n622 & ~n637 ) | ( n622 & n685 ) | ( ~n637 & n685 ) ;
  assign n688 = ( n637 & ~n686 ) | ( n637 & n687 ) | ( ~n686 & n687 ) ;
  assign n689 = ( ~n639 & n682 ) | ( ~n639 & n688 ) | ( n682 & n688 ) ;
  assign n690 = ( n639 & n682 ) | ( n639 & n688 ) | ( n682 & n688 ) ;
  assign n691 = ( n639 & n689 ) | ( n639 & ~n690 ) | ( n689 & ~n690 ) ;
  assign n692 = ( n643 & n645 ) | ( n643 & n691 ) | ( n645 & n691 ) ;
  assign n693 = ( n643 & ~n645 ) | ( n643 & n691 ) | ( ~n645 & n691 ) ;
  assign n694 = ( n645 & ~n692 ) | ( n645 & n693 ) | ( ~n692 & n693 ) ;
  assign n695 = x1 & x24 ;
  assign n696 = ( x13 & ~n648 ) | ( x13 & n652 ) | ( ~n648 & n652 ) ;
  assign n697 = ( n675 & n695 ) | ( n675 & n696 ) | ( n695 & n696 ) ;
  assign n698 = ( ~n675 & n695 ) | ( ~n675 & n696 ) | ( n695 & n696 ) ;
  assign n699 = ( n675 & ~n697 ) | ( n675 & n698 ) | ( ~n697 & n698 ) ;
  assign n700 = x12 & x13 ;
  assign n701 = x11 & x14 ;
  assign n702 = x5 & x20 ;
  assign n703 = ( ~n700 & n701 ) | ( ~n700 & n702 ) | ( n701 & n702 ) ;
  assign n704 = ( n700 & n701 ) | ( n700 & n702 ) | ( n701 & n702 ) ;
  assign n705 = ( n700 & n703 ) | ( n700 & ~n704 ) | ( n703 & ~n704 ) ;
  assign n706 = ( n684 & ~n699 ) | ( n684 & n705 ) | ( ~n699 & n705 ) ;
  assign n707 = ( n684 & n699 ) | ( n684 & n705 ) | ( n699 & n705 ) ;
  assign n708 = ( n699 & n706 ) | ( n699 & ~n707 ) | ( n706 & ~n707 ) ;
  assign n709 = x10 & x15 ;
  assign n710 = x0 & x25 ;
  assign n711 = x2 & x23 ;
  assign n712 = ( ~n709 & n710 ) | ( ~n709 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( n709 & n710 ) | ( n709 & n711 ) | ( n710 & n711 ) ;
  assign n714 = ( n709 & n712 ) | ( n709 & ~n713 ) | ( n712 & ~n713 ) ;
  assign n715 = x9 & x16 ;
  assign n716 = x7 & x18 ;
  assign n717 = x8 & x17 ;
  assign n718 = ( ~n715 & n716 ) | ( ~n715 & n717 ) | ( n716 & n717 ) ;
  assign n719 = ( n715 & n716 ) | ( n715 & n717 ) | ( n716 & n717 ) ;
  assign n720 = ( n715 & n718 ) | ( n715 & ~n719 ) | ( n718 & ~n719 ) ;
  assign n721 = x4 & x21 ;
  assign n722 = x6 & x19 ;
  assign n723 = x3 & x22 ;
  assign n724 = ( ~n721 & n722 ) | ( ~n721 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ( n721 & n722 ) | ( n721 & n723 ) | ( n722 & n723 ) ;
  assign n726 = ( n721 & n724 ) | ( n721 & ~n725 ) | ( n724 & ~n725 ) ;
  assign n727 = ( ~n714 & n720 ) | ( ~n714 & n726 ) | ( n720 & n726 ) ;
  assign n728 = ( n714 & n720 ) | ( n714 & n726 ) | ( n720 & n726 ) ;
  assign n729 = ( n714 & n727 ) | ( n714 & ~n728 ) | ( n727 & ~n728 ) ;
  assign n730 = ( n686 & n708 ) | ( n686 & n729 ) | ( n708 & n729 ) ;
  assign n731 = ( ~n686 & n708 ) | ( ~n686 & n729 ) | ( n708 & n729 ) ;
  assign n732 = ( n686 & ~n730 ) | ( n686 & n731 ) | ( ~n730 & n731 ) ;
  assign n733 = ( ~n654 & n661 ) | ( ~n654 & n669 ) | ( n661 & n669 ) ;
  assign n734 = ( n654 & n661 ) | ( n654 & n669 ) | ( n661 & n669 ) ;
  assign n735 = ( n654 & n733 ) | ( n654 & ~n734 ) | ( n733 & ~n734 ) ;
  assign n736 = ( n663 & n678 ) | ( n663 & n735 ) | ( n678 & n735 ) ;
  assign n737 = ( n663 & n678 ) | ( n663 & ~n735 ) | ( n678 & ~n735 ) ;
  assign n738 = ( n735 & ~n736 ) | ( n735 & n737 ) | ( ~n736 & n737 ) ;
  assign n739 = ( n680 & n732 ) | ( n680 & n738 ) | ( n732 & n738 ) ;
  assign n740 = ( n680 & ~n732 ) | ( n680 & n738 ) | ( ~n732 & n738 ) ;
  assign n741 = ( n732 & ~n739 ) | ( n732 & n740 ) | ( ~n739 & n740 ) ;
  assign n742 = ( n690 & n692 ) | ( n690 & n741 ) | ( n692 & n741 ) ;
  assign n743 = ( n690 & ~n692 ) | ( n690 & n741 ) | ( ~n692 & n741 ) ;
  assign n744 = ( n692 & ~n742 ) | ( n692 & n743 ) | ( ~n742 & n743 ) ;
  assign n745 = x5 & x21 ;
  assign n746 = x4 & x22 ;
  assign n747 = x6 & x20 ;
  assign n748 = ( ~n745 & n746 ) | ( ~n745 & n747 ) | ( n746 & n747 ) ;
  assign n749 = ( n745 & n746 ) | ( n745 & n747 ) | ( n746 & n747 ) ;
  assign n750 = ( n745 & n748 ) | ( n745 & ~n749 ) | ( n748 & ~n749 ) ;
  assign n751 = x7 & x19 ;
  assign n752 = x2 & x24 ;
  assign n753 = x3 & x23 ;
  assign n754 = ( ~n751 & n752 ) | ( ~n751 & n753 ) | ( n752 & n753 ) ;
  assign n755 = ( n751 & n752 ) | ( n751 & n753 ) | ( n752 & n753 ) ;
  assign n756 = ( n751 & n754 ) | ( n751 & ~n755 ) | ( n754 & ~n755 ) ;
  assign n757 = x10 & x16 ;
  assign n758 = x9 & x17 ;
  assign n759 = x11 & x15 ;
  assign n760 = ( ~n757 & n758 ) | ( ~n757 & n759 ) | ( n758 & n759 ) ;
  assign n761 = ( n757 & n758 ) | ( n757 & n759 ) | ( n758 & n759 ) ;
  assign n762 = ( n757 & n760 ) | ( n757 & ~n761 ) | ( n760 & ~n761 ) ;
  assign n763 = ( ~n750 & n756 ) | ( ~n750 & n762 ) | ( n756 & n762 ) ;
  assign n764 = ( n750 & n756 ) | ( n750 & n762 ) | ( n756 & n762 ) ;
  assign n765 = ( n750 & n763 ) | ( n750 & ~n764 ) | ( n763 & ~n764 ) ;
  assign n766 = ( n650 & n675 ) | ( n650 & ~n699 ) | ( n675 & ~n699 ) ;
  assign n767 = x13 & n695 ;
  assign n768 = x0 & x26 ;
  assign n769 = x8 & x18 ;
  assign n770 = ( ~n767 & n768 ) | ( ~n767 & n769 ) | ( n768 & n769 ) ;
  assign n771 = ( n767 & n768 ) | ( n767 & n769 ) | ( n768 & n769 ) ;
  assign n772 = ( n767 & n770 ) | ( n767 & ~n771 ) | ( n770 & ~n771 ) ;
  assign n773 = ( n713 & n719 ) | ( n713 & ~n772 ) | ( n719 & ~n772 ) ;
  assign n774 = ( n713 & n719 ) | ( n713 & n772 ) | ( n719 & n772 ) ;
  assign n775 = ( n772 & n773 ) | ( n772 & ~n774 ) | ( n773 & ~n774 ) ;
  assign n776 = ( n734 & n766 ) | ( n734 & n775 ) | ( n766 & n775 ) ;
  assign n777 = ( n734 & ~n766 ) | ( n734 & n775 ) | ( ~n766 & n775 ) ;
  assign n778 = ( n766 & ~n776 ) | ( n766 & n777 ) | ( ~n776 & n777 ) ;
  assign n779 = ( n736 & n765 ) | ( n736 & n778 ) | ( n765 & n778 ) ;
  assign n780 = ( n736 & ~n765 ) | ( n736 & n778 ) | ( ~n765 & n778 ) ;
  assign n781 = ( n765 & ~n779 ) | ( n765 & n780 ) | ( ~n779 & n780 ) ;
  assign n782 = x1 & x25 ;
  assign n783 = x12 & x14 ;
  assign n784 = n782 | n783 ;
  assign n785 = x14 & x25 ;
  assign n786 = n251 & n785 ;
  assign n787 = n784 & ~n786 ;
  assign n788 = ( ~n704 & n725 ) | ( ~n704 & n787 ) | ( n725 & n787 ) ;
  assign n789 = ( n704 & n725 ) | ( n704 & n787 ) | ( n725 & n787 ) ;
  assign n790 = ( n704 & n788 ) | ( n704 & ~n789 ) | ( n788 & ~n789 ) ;
  assign n791 = ( ~n707 & n728 ) | ( ~n707 & n790 ) | ( n728 & n790 ) ;
  assign n792 = ( n707 & n728 ) | ( n707 & n790 ) | ( n728 & n790 ) ;
  assign n793 = ( n707 & n791 ) | ( n707 & ~n792 ) | ( n791 & ~n792 ) ;
  assign n794 = ( n730 & n781 ) | ( n730 & n793 ) | ( n781 & n793 ) ;
  assign n795 = ( n730 & ~n781 ) | ( n730 & n793 ) | ( ~n781 & n793 ) ;
  assign n796 = ( n781 & ~n794 ) | ( n781 & n795 ) | ( ~n794 & n795 ) ;
  assign n797 = ( n739 & n742 ) | ( n739 & n796 ) | ( n742 & n796 ) ;
  assign n798 = ( n739 & ~n742 ) | ( n739 & n796 ) | ( ~n742 & n796 ) ;
  assign n799 = ( n742 & ~n797 ) | ( n742 & n798 ) | ( ~n797 & n798 ) ;
  assign n800 = ( n764 & n774 ) | ( n764 & ~n789 ) | ( n774 & ~n789 ) ;
  assign n801 = ( n764 & n774 ) | ( n764 & n789 ) | ( n774 & n789 ) ;
  assign n802 = ( n789 & n800 ) | ( n789 & ~n801 ) | ( n800 & ~n801 ) ;
  assign n803 = x8 & x19 ;
  assign n804 = x9 & x18 ;
  assign n805 = ( ~n399 & n803 ) | ( ~n399 & n804 ) | ( n803 & n804 ) ;
  assign n806 = ( n399 & n803 ) | ( n399 & n804 ) | ( n803 & n804 ) ;
  assign n807 = ( n399 & n805 ) | ( n399 & ~n806 ) | ( n805 & ~n806 ) ;
  assign n808 = x2 & x25 ;
  assign n809 = x11 & x16 ;
  assign n810 = x7 & x20 ;
  assign n811 = ( ~n808 & n809 ) | ( ~n808 & n810 ) | ( n809 & n810 ) ;
  assign n812 = ( n808 & n809 ) | ( n808 & n810 ) | ( n809 & n810 ) ;
  assign n813 = ( n808 & n811 ) | ( n808 & ~n812 ) | ( n811 & ~n812 ) ;
  assign n814 = ( ~n771 & n807 ) | ( ~n771 & n813 ) | ( n807 & n813 ) ;
  assign n815 = ( n771 & n807 ) | ( n771 & n813 ) | ( n807 & n813 ) ;
  assign n816 = ( n771 & n814 ) | ( n771 & ~n815 ) | ( n814 & ~n815 ) ;
  assign n817 = ( n792 & n802 ) | ( n792 & n816 ) | ( n802 & n816 ) ;
  assign n818 = ( ~n792 & n802 ) | ( ~n792 & n816 ) | ( n802 & n816 ) ;
  assign n819 = ( n792 & ~n817 ) | ( n792 & n818 ) | ( ~n817 & n818 ) ;
  assign n820 = x1 & x26 ;
  assign n821 = x14 & ~n786 ;
  assign n822 = x0 & x27 ;
  assign n823 = ( ~n820 & n821 ) | ( ~n820 & n822 ) | ( n821 & n822 ) ;
  assign n824 = ( n820 & n821 ) | ( n820 & n822 ) | ( n821 & n822 ) ;
  assign n825 = ( n820 & n823 ) | ( n820 & ~n824 ) | ( n823 & ~n824 ) ;
  assign n826 = x3 & x24 ;
  assign n827 = x4 & x23 ;
  assign n828 = x6 & x21 ;
  assign n829 = ( ~n826 & n827 ) | ( ~n826 & n828 ) | ( n827 & n828 ) ;
  assign n830 = ( n826 & n827 ) | ( n826 & n828 ) | ( n827 & n828 ) ;
  assign n831 = ( n826 & n829 ) | ( n826 & ~n830 ) | ( n829 & ~n830 ) ;
  assign n832 = x13 & x14 ;
  assign n833 = x5 & x22 ;
  assign n834 = x12 & x15 ;
  assign n835 = ( ~n832 & n833 ) | ( ~n832 & n834 ) | ( n833 & n834 ) ;
  assign n836 = ( n832 & n833 ) | ( n832 & n834 ) | ( n833 & n834 ) ;
  assign n837 = ( n832 & n835 ) | ( n832 & ~n836 ) | ( n835 & ~n836 ) ;
  assign n838 = ( n825 & n831 ) | ( n825 & n837 ) | ( n831 & n837 ) ;
  assign n839 = ( ~n825 & n831 ) | ( ~n825 & n837 ) | ( n831 & n837 ) ;
  assign n840 = ( n825 & ~n838 ) | ( n825 & n839 ) | ( ~n838 & n839 ) ;
  assign n841 = ( ~n749 & n755 ) | ( ~n749 & n761 ) | ( n755 & n761 ) ;
  assign n842 = ( n749 & n755 ) | ( n749 & n761 ) | ( n755 & n761 ) ;
  assign n843 = ( n749 & n841 ) | ( n749 & ~n842 ) | ( n841 & ~n842 ) ;
  assign n844 = ( n776 & n840 ) | ( n776 & n843 ) | ( n840 & n843 ) ;
  assign n845 = ( ~n776 & n840 ) | ( ~n776 & n843 ) | ( n840 & n843 ) ;
  assign n846 = ( n776 & ~n844 ) | ( n776 & n845 ) | ( ~n844 & n845 ) ;
  assign n847 = ( ~n779 & n819 ) | ( ~n779 & n846 ) | ( n819 & n846 ) ;
  assign n848 = ( n779 & n819 ) | ( n779 & n846 ) | ( n819 & n846 ) ;
  assign n849 = ( n779 & n847 ) | ( n779 & ~n848 ) | ( n847 & ~n848 ) ;
  assign n850 = ( n794 & ~n797 ) | ( n794 & n849 ) | ( ~n797 & n849 ) ;
  assign n851 = ( n794 & n797 ) | ( n794 & n849 ) | ( n797 & n849 ) ;
  assign n852 = ( n797 & n850 ) | ( n797 & ~n851 ) | ( n850 & ~n851 ) ;
  assign n853 = ( n806 & n812 ) | ( n806 & ~n830 ) | ( n812 & ~n830 ) ;
  assign n854 = ( n806 & n812 ) | ( n806 & n830 ) | ( n812 & n830 ) ;
  assign n855 = ( n830 & n853 ) | ( n830 & ~n854 ) | ( n853 & ~n854 ) ;
  assign n856 = x2 & x26 ;
  assign n857 = ( ~n437 & n533 ) | ( ~n437 & n856 ) | ( n533 & n856 ) ;
  assign n858 = ( n437 & n533 ) | ( n437 & n856 ) | ( n533 & n856 ) ;
  assign n859 = ( n437 & n857 ) | ( n437 & ~n858 ) | ( n857 & ~n858 ) ;
  assign n860 = x11 & x17 ;
  assign n861 = x0 & x28 ;
  assign n862 = x12 & x16 ;
  assign n863 = ( ~n860 & n861 ) | ( ~n860 & n862 ) | ( n861 & n862 ) ;
  assign n864 = ( n860 & n861 ) | ( n860 & n862 ) | ( n861 & n862 ) ;
  assign n865 = ( n860 & n863 ) | ( n860 & ~n864 ) | ( n863 & ~n864 ) ;
  assign n866 = ( ~n842 & n859 ) | ( ~n842 & n865 ) | ( n859 & n865 ) ;
  assign n867 = ( n842 & n859 ) | ( n842 & n865 ) | ( n859 & n865 ) ;
  assign n868 = ( n842 & n866 ) | ( n842 & ~n867 ) | ( n866 & ~n867 ) ;
  assign n869 = ( n801 & n855 ) | ( n801 & n868 ) | ( n855 & n868 ) ;
  assign n870 = ( ~n801 & n855 ) | ( ~n801 & n868 ) | ( n855 & n868 ) ;
  assign n871 = ( n801 & ~n869 ) | ( n801 & n870 ) | ( ~n869 & n870 ) ;
  assign n872 = ( n817 & ~n848 ) | ( n817 & n871 ) | ( ~n848 & n871 ) ;
  assign n873 = ( n817 & n848 ) | ( n817 & n871 ) | ( n848 & n871 ) ;
  assign n874 = ( n848 & n872 ) | ( n848 & ~n873 ) | ( n872 & ~n873 ) ;
  assign n875 = x14 & n820 ;
  assign n876 = ( n786 & n824 ) | ( n786 & ~n875 ) | ( n824 & ~n875 ) ;
  assign n877 = x3 & x25 ;
  assign n878 = x8 & x20 ;
  assign n879 = x4 & x24 ;
  assign n880 = ( ~n877 & n878 ) | ( ~n877 & n879 ) | ( n878 & n879 ) ;
  assign n881 = ( n877 & n878 ) | ( n877 & n879 ) | ( n878 & n879 ) ;
  assign n882 = ( n877 & n880 ) | ( n877 & ~n881 ) | ( n880 & ~n881 ) ;
  assign n883 = x5 & x23 ;
  assign n884 = x6 & x22 ;
  assign n885 = x7 & x21 ;
  assign n886 = ( ~n883 & n884 ) | ( ~n883 & n885 ) | ( n884 & n885 ) ;
  assign n887 = ( n883 & n884 ) | ( n883 & n885 ) | ( n884 & n885 ) ;
  assign n888 = ( n883 & n886 ) | ( n883 & ~n887 ) | ( n886 & ~n887 ) ;
  assign n889 = ( ~n876 & n882 ) | ( ~n876 & n888 ) | ( n882 & n888 ) ;
  assign n890 = ( n876 & n882 ) | ( n876 & n888 ) | ( n882 & n888 ) ;
  assign n891 = ( n876 & n889 ) | ( n876 & ~n890 ) | ( n889 & ~n890 ) ;
  assign n892 = x1 & x27 ;
  assign n893 = x13 & x15 ;
  assign n894 = n892 | n893 ;
  assign n895 = x15 & x27 ;
  assign n896 = n278 & n895 ;
  assign n897 = n894 & ~n896 ;
  assign n898 = ( ~n836 & n875 ) | ( ~n836 & n897 ) | ( n875 & n897 ) ;
  assign n899 = ( n836 & n875 ) | ( n836 & n897 ) | ( n875 & n897 ) ;
  assign n900 = ( n836 & n898 ) | ( n836 & ~n899 ) | ( n898 & ~n899 ) ;
  assign n901 = ( n815 & n838 ) | ( n815 & n900 ) | ( n838 & n900 ) ;
  assign n902 = ( n815 & ~n838 ) | ( n815 & n900 ) | ( ~n838 & n900 ) ;
  assign n903 = ( n838 & ~n901 ) | ( n838 & n902 ) | ( ~n901 & n902 ) ;
  assign n904 = ( n844 & n891 ) | ( n844 & n903 ) | ( n891 & n903 ) ;
  assign n905 = ( ~n844 & n891 ) | ( ~n844 & n903 ) | ( n891 & n903 ) ;
  assign n906 = ( n844 & ~n904 ) | ( n844 & n905 ) | ( ~n904 & n905 ) ;
  assign n907 = ( n851 & n874 ) | ( n851 & n906 ) | ( n874 & n906 ) ;
  assign n908 = ( ~n851 & n874 ) | ( ~n851 & n906 ) | ( n874 & n906 ) ;
  assign n909 = ( n851 & ~n907 ) | ( n851 & n908 ) | ( ~n907 & n908 ) ;
  assign n910 = x2 & x27 ;
  assign n911 = x0 & x29 ;
  assign n912 = ( ~n896 & n910 ) | ( ~n896 & n911 ) | ( n910 & n911 ) ;
  assign n913 = ( n896 & n910 ) | ( n896 & n911 ) | ( n910 & n911 ) ;
  assign n914 = ( n896 & n912 ) | ( n896 & ~n913 ) | ( n912 & ~n913 ) ;
  assign n915 = ( n858 & n864 ) | ( n858 & ~n914 ) | ( n864 & ~n914 ) ;
  assign n916 = ( n858 & n864 ) | ( n858 & n914 ) | ( n864 & n914 ) ;
  assign n917 = ( n914 & n915 ) | ( n914 & ~n916 ) | ( n915 & ~n916 ) ;
  assign n918 = ( n867 & n890 ) | ( n867 & n917 ) | ( n890 & n917 ) ;
  assign n919 = ( n867 & n890 ) | ( n867 & ~n917 ) | ( n890 & ~n917 ) ;
  assign n920 = ( n917 & ~n918 ) | ( n917 & n919 ) | ( ~n918 & n919 ) ;
  assign n921 = ( n869 & n901 ) | ( n869 & ~n920 ) | ( n901 & ~n920 ) ;
  assign n922 = ( n869 & n901 ) | ( n869 & n920 ) | ( n901 & n920 ) ;
  assign n923 = ( n920 & n921 ) | ( n920 & ~n922 ) | ( n921 & ~n922 ) ;
  assign n924 = x14 & x15 ;
  assign n925 = x6 & x23 ;
  assign n926 = x13 & x16 ;
  assign n927 = ( ~n924 & n925 ) | ( ~n924 & n926 ) | ( n925 & n926 ) ;
  assign n928 = ( n924 & n925 ) | ( n924 & n926 ) | ( n925 & n926 ) ;
  assign n929 = ( n924 & n927 ) | ( n924 & ~n928 ) | ( n927 & ~n928 ) ;
  assign n930 = ( n854 & n899 ) | ( n854 & ~n929 ) | ( n899 & ~n929 ) ;
  assign n931 = ( n854 & n899 ) | ( n854 & n929 ) | ( n899 & n929 ) ;
  assign n932 = ( n929 & n930 ) | ( n929 & ~n931 ) | ( n930 & ~n931 ) ;
  assign n933 = x1 & x28 ;
  assign n934 = x15 | n933 ;
  assign n935 = x28 & n331 ;
  assign n936 = n934 & ~n935 ;
  assign n937 = ( n881 & n887 ) | ( n881 & ~n936 ) | ( n887 & ~n936 ) ;
  assign n938 = ( n881 & n887 ) | ( n881 & n936 ) | ( n887 & n936 ) ;
  assign n939 = ( n936 & n937 ) | ( n936 & ~n938 ) | ( n937 & ~n938 ) ;
  assign n940 = x3 & x26 ;
  assign n941 = x8 & x21 ;
  assign n942 = x12 & x17 ;
  assign n943 = ( ~n940 & n941 ) | ( ~n940 & n942 ) | ( n941 & n942 ) ;
  assign n944 = ( n940 & n941 ) | ( n940 & n942 ) | ( n941 & n942 ) ;
  assign n945 = ( n940 & n943 ) | ( n940 & ~n944 ) | ( n943 & ~n944 ) ;
  assign n946 = x11 & x18 ;
  assign n947 = x9 & x20 ;
  assign n948 = x10 & x19 ;
  assign n949 = ( ~n946 & n947 ) | ( ~n946 & n948 ) | ( n947 & n948 ) ;
  assign n950 = ( n946 & n947 ) | ( n946 & n948 ) | ( n947 & n948 ) ;
  assign n951 = ( n946 & n949 ) | ( n946 & ~n950 ) | ( n949 & ~n950 ) ;
  assign n952 = x4 & x25 ;
  assign n953 = x5 & x24 ;
  assign n954 = x7 & x22 ;
  assign n955 = ( ~n952 & n953 ) | ( ~n952 & n954 ) | ( n953 & n954 ) ;
  assign n956 = ( n952 & n953 ) | ( n952 & n954 ) | ( n953 & n954 ) ;
  assign n957 = ( n952 & n955 ) | ( n952 & ~n956 ) | ( n955 & ~n956 ) ;
  assign n958 = ( ~n945 & n951 ) | ( ~n945 & n957 ) | ( n951 & n957 ) ;
  assign n959 = ( n945 & n951 ) | ( n945 & n957 ) | ( n951 & n957 ) ;
  assign n960 = ( n945 & n958 ) | ( n945 & ~n959 ) | ( n958 & ~n959 ) ;
  assign n961 = ( n932 & n939 ) | ( n932 & n960 ) | ( n939 & n960 ) ;
  assign n962 = ( ~n932 & n939 ) | ( ~n932 & n960 ) | ( n939 & n960 ) ;
  assign n963 = ( n932 & ~n961 ) | ( n932 & n962 ) | ( ~n961 & n962 ) ;
  assign n964 = ( n904 & n923 ) | ( n904 & n963 ) | ( n923 & n963 ) ;
  assign n965 = ( ~n904 & n923 ) | ( ~n904 & n963 ) | ( n923 & n963 ) ;
  assign n966 = ( n904 & ~n964 ) | ( n904 & n965 ) | ( ~n964 & n965 ) ;
  assign n967 = ( n873 & ~n907 ) | ( n873 & n966 ) | ( ~n907 & n966 ) ;
  assign n968 = ( n873 & n907 ) | ( n873 & n966 ) | ( n907 & n966 ) ;
  assign n969 = ( n907 & n967 ) | ( n907 & ~n968 ) | ( n967 & ~n968 ) ;
  assign n970 = x1 & x29 ;
  assign n971 = x14 & x16 ;
  assign n972 = n970 | n971 ;
  assign n973 = x16 & x29 ;
  assign n974 = n294 & n973 ;
  assign n975 = n972 & ~n974 ;
  assign n976 = x0 & x30 ;
  assign n977 = ( n935 & n975 ) | ( n935 & n976 ) | ( n975 & n976 ) ;
  assign n978 = ( n935 & ~n975 ) | ( n935 & n976 ) | ( ~n975 & n976 ) ;
  assign n979 = ( n975 & ~n977 ) | ( n975 & n978 ) | ( ~n977 & n978 ) ;
  assign n980 = ( n916 & n938 ) | ( n916 & n979 ) | ( n938 & n979 ) ;
  assign n981 = ( ~n916 & n938 ) | ( ~n916 & n979 ) | ( n938 & n979 ) ;
  assign n982 = ( n916 & ~n980 ) | ( n916 & n981 ) | ( ~n980 & n981 ) ;
  assign n983 = ( ~n913 & n944 ) | ( ~n913 & n950 ) | ( n944 & n950 ) ;
  assign n984 = ( n913 & n944 ) | ( n913 & n950 ) | ( n944 & n950 ) ;
  assign n985 = ( n913 & n983 ) | ( n913 & ~n984 ) | ( n983 & ~n984 ) ;
  assign n986 = x13 & x17 ;
  assign n987 = x2 & x28 ;
  assign n988 = x9 & x21 ;
  assign n989 = ( ~n986 & n987 ) | ( ~n986 & n988 ) | ( n987 & n988 ) ;
  assign n990 = ( n986 & n987 ) | ( n986 & n988 ) | ( n987 & n988 ) ;
  assign n991 = ( n986 & n989 ) | ( n986 & ~n990 ) | ( n989 & ~n990 ) ;
  assign n992 = ( n928 & n956 ) | ( n928 & ~n991 ) | ( n956 & ~n991 ) ;
  assign n993 = ( n928 & n956 ) | ( n928 & n991 ) | ( n956 & n991 ) ;
  assign n994 = ( n991 & n992 ) | ( n991 & ~n993 ) | ( n992 & ~n993 ) ;
  assign n995 = ( n959 & n985 ) | ( n959 & n994 ) | ( n985 & n994 ) ;
  assign n996 = ( n959 & ~n985 ) | ( n959 & n994 ) | ( ~n985 & n994 ) ;
  assign n997 = ( n985 & ~n995 ) | ( n985 & n996 ) | ( ~n995 & n996 ) ;
  assign n998 = ( n961 & n982 ) | ( n961 & n997 ) | ( n982 & n997 ) ;
  assign n999 = ( ~n961 & n982 ) | ( ~n961 & n997 ) | ( n982 & n997 ) ;
  assign n1000 = ( n961 & ~n998 ) | ( n961 & n999 ) | ( ~n998 & n999 ) ;
  assign n1001 = x3 & x27 ;
  assign n1002 = x4 & x26 ;
  assign n1003 = x8 & x22 ;
  assign n1004 = ( ~n1001 & n1002 ) | ( ~n1001 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1005 = ( n1001 & n1002 ) | ( n1001 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1006 = ( n1001 & n1004 ) | ( n1001 & ~n1005 ) | ( n1004 & ~n1005 ) ;
  assign n1007 = x11 & x19 ;
  assign n1008 = x10 & x20 ;
  assign n1009 = x12 & x18 ;
  assign n1010 = ( ~n1007 & n1008 ) | ( ~n1007 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1011 = ( n1007 & n1008 ) | ( n1007 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1012 = ( n1007 & n1010 ) | ( n1007 & ~n1011 ) | ( n1010 & ~n1011 ) ;
  assign n1013 = x7 & x23 ;
  assign n1014 = x6 & x24 ;
  assign n1015 = x5 & x25 ;
  assign n1016 = ( ~n1013 & n1014 ) | ( ~n1013 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = ( n1013 & n1014 ) | ( n1013 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1018 = ( n1013 & n1016 ) | ( n1013 & ~n1017 ) | ( n1016 & ~n1017 ) ;
  assign n1019 = ( ~n1006 & n1012 ) | ( ~n1006 & n1018 ) | ( n1012 & n1018 ) ;
  assign n1020 = ( n1006 & n1012 ) | ( n1006 & n1018 ) | ( n1012 & n1018 ) ;
  assign n1021 = ( n1006 & n1019 ) | ( n1006 & ~n1020 ) | ( n1019 & ~n1020 ) ;
  assign n1022 = ( n918 & n931 ) | ( n918 & ~n1021 ) | ( n931 & ~n1021 ) ;
  assign n1023 = ( n918 & n931 ) | ( n918 & n1021 ) | ( n931 & n1021 ) ;
  assign n1024 = ( n1021 & n1022 ) | ( n1021 & ~n1023 ) | ( n1022 & ~n1023 ) ;
  assign n1025 = ( ~n922 & n1000 ) | ( ~n922 & n1024 ) | ( n1000 & n1024 ) ;
  assign n1026 = ( n922 & n1000 ) | ( n922 & n1024 ) | ( n1000 & n1024 ) ;
  assign n1027 = ( n922 & n1025 ) | ( n922 & ~n1026 ) | ( n1025 & ~n1026 ) ;
  assign n1028 = ( n964 & ~n968 ) | ( n964 & n1027 ) | ( ~n968 & n1027 ) ;
  assign n1029 = ( n964 & n968 ) | ( n964 & n1027 ) | ( n968 & n1027 ) ;
  assign n1030 = ( n968 & n1028 ) | ( n968 & ~n1029 ) | ( n1028 & ~n1029 ) ;
  assign n1031 = ( ~n990 & n1005 ) | ( ~n990 & n1011 ) | ( n1005 & n1011 ) ;
  assign n1032 = ( n990 & n1005 ) | ( n990 & n1011 ) | ( n1005 & n1011 ) ;
  assign n1033 = ( n990 & n1031 ) | ( n990 & ~n1032 ) | ( n1031 & ~n1032 ) ;
  assign n1034 = ( n980 & n1020 ) | ( n980 & ~n1033 ) | ( n1020 & ~n1033 ) ;
  assign n1035 = ( n980 & n1020 ) | ( n980 & n1033 ) | ( n1020 & n1033 ) ;
  assign n1036 = ( n1033 & n1034 ) | ( n1033 & ~n1035 ) | ( n1034 & ~n1035 ) ;
  assign n1037 = x1 & x30 ;
  assign n1038 = x16 & ~n974 ;
  assign n1039 = ( n1017 & n1037 ) | ( n1017 & ~n1038 ) | ( n1037 & ~n1038 ) ;
  assign n1040 = ( ~n1017 & n1037 ) | ( ~n1017 & n1038 ) | ( n1037 & n1038 ) ;
  assign n1041 = ( ~n1037 & n1039 ) | ( ~n1037 & n1040 ) | ( n1039 & n1040 ) ;
  assign n1042 = ( n984 & n993 ) | ( n984 & n1041 ) | ( n993 & n1041 ) ;
  assign n1043 = ( ~n984 & n993 ) | ( ~n984 & n1041 ) | ( n993 & n1041 ) ;
  assign n1044 = ( n984 & ~n1042 ) | ( n984 & n1043 ) | ( ~n1042 & n1043 ) ;
  assign n1045 = ( n1023 & n1036 ) | ( n1023 & n1044 ) | ( n1036 & n1044 ) ;
  assign n1046 = ( ~n1023 & n1036 ) | ( ~n1023 & n1044 ) | ( n1036 & n1044 ) ;
  assign n1047 = ( n1023 & ~n1045 ) | ( n1023 & n1046 ) | ( ~n1045 & n1046 ) ;
  assign n1048 = x9 & x22 ;
  assign n1049 = x0 & x31 ;
  assign n1050 = ( ~n585 & n1048 ) | ( ~n585 & n1049 ) | ( n1048 & n1049 ) ;
  assign n1051 = ( n585 & n1048 ) | ( n585 & n1049 ) | ( n1048 & n1049 ) ;
  assign n1052 = ( n585 & n1050 ) | ( n585 & ~n1051 ) | ( n1050 & ~n1051 ) ;
  assign n1053 = x12 & x19 ;
  assign n1054 = x11 & x20 ;
  assign n1055 = x13 & x18 ;
  assign n1056 = ( ~n1053 & n1054 ) | ( ~n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( n1053 & n1054 ) | ( n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1058 = ( n1053 & n1056 ) | ( n1053 & ~n1057 ) | ( n1056 & ~n1057 ) ;
  assign n1059 = ( ~n977 & n1052 ) | ( ~n977 & n1058 ) | ( n1052 & n1058 ) ;
  assign n1060 = ( n977 & n1052 ) | ( n977 & n1058 ) | ( n1052 & n1058 ) ;
  assign n1061 = ( n977 & n1059 ) | ( n977 & ~n1060 ) | ( n1059 & ~n1060 ) ;
  assign n1062 = x3 & x28 ;
  assign n1063 = x2 & x29 ;
  assign n1064 = x4 & x27 ;
  assign n1065 = ( ~n1062 & n1063 ) | ( ~n1062 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1066 = ( n1062 & n1063 ) | ( n1062 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1067 = ( n1062 & n1065 ) | ( n1062 & ~n1066 ) | ( n1065 & ~n1066 ) ;
  assign n1068 = x7 & x24 ;
  assign n1069 = x8 & x23 ;
  assign n1070 = x5 & x26 ;
  assign n1071 = ( ~n1068 & n1069 ) | ( ~n1068 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1072 = ( n1068 & n1069 ) | ( n1068 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1073 = ( n1068 & n1071 ) | ( n1068 & ~n1072 ) | ( n1071 & ~n1072 ) ;
  assign n1074 = x15 & x16 ;
  assign n1075 = x14 & x17 ;
  assign n1076 = x6 & x25 ;
  assign n1077 = ( ~n1074 & n1075 ) | ( ~n1074 & n1076 ) | ( n1075 & n1076 ) ;
  assign n1078 = ( n1074 & n1075 ) | ( n1074 & n1076 ) | ( n1075 & n1076 ) ;
  assign n1079 = ( n1074 & n1077 ) | ( n1074 & ~n1078 ) | ( n1077 & ~n1078 ) ;
  assign n1080 = ( ~n1067 & n1073 ) | ( ~n1067 & n1079 ) | ( n1073 & n1079 ) ;
  assign n1081 = ( n1067 & n1073 ) | ( n1067 & n1079 ) | ( n1073 & n1079 ) ;
  assign n1082 = ( n1067 & n1080 ) | ( n1067 & ~n1081 ) | ( n1080 & ~n1081 ) ;
  assign n1083 = ( n995 & n1061 ) | ( n995 & n1082 ) | ( n1061 & n1082 ) ;
  assign n1084 = ( ~n995 & n1061 ) | ( ~n995 & n1082 ) | ( n1061 & n1082 ) ;
  assign n1085 = ( n995 & ~n1083 ) | ( n995 & n1084 ) | ( ~n1083 & n1084 ) ;
  assign n1086 = ( n998 & n1047 ) | ( n998 & n1085 ) | ( n1047 & n1085 ) ;
  assign n1087 = ( n998 & ~n1047 ) | ( n998 & n1085 ) | ( ~n1047 & n1085 ) ;
  assign n1088 = ( n1047 & ~n1086 ) | ( n1047 & n1087 ) | ( ~n1086 & n1087 ) ;
  assign n1089 = ( n1026 & ~n1029 ) | ( n1026 & n1088 ) | ( ~n1029 & n1088 ) ;
  assign n1090 = ( n1026 & n1029 ) | ( n1026 & n1088 ) | ( n1029 & n1088 ) ;
  assign n1091 = ( n1029 & n1089 ) | ( n1029 & ~n1090 ) | ( n1089 & ~n1090 ) ;
  assign n1092 = ( ~n1032 & n1060 ) | ( ~n1032 & n1081 ) | ( n1060 & n1081 ) ;
  assign n1093 = ( n1032 & n1060 ) | ( n1032 & n1081 ) | ( n1060 & n1081 ) ;
  assign n1094 = ( n1032 & n1092 ) | ( n1032 & ~n1093 ) | ( n1092 & ~n1093 ) ;
  assign n1095 = ( n1051 & n1057 ) | ( n1051 & ~n1066 ) | ( n1057 & ~n1066 ) ;
  assign n1096 = ( n1051 & n1057 ) | ( n1051 & n1066 ) | ( n1057 & n1066 ) ;
  assign n1097 = ( n1066 & n1095 ) | ( n1066 & ~n1096 ) | ( n1095 & ~n1096 ) ;
  assign n1098 = x1 & x31 ;
  assign n1099 = x15 & x17 ;
  assign n1100 = n1098 & n1099 ;
  assign n1101 = n1098 | n1099 ;
  assign n1102 = ~n1100 & n1101 ;
  assign n1103 = ( n1072 & ~n1078 ) | ( n1072 & n1102 ) | ( ~n1078 & n1102 ) ;
  assign n1104 = ( n1072 & n1078 ) | ( n1072 & n1102 ) | ( n1078 & n1102 ) ;
  assign n1105 = ( n1078 & n1103 ) | ( n1078 & ~n1104 ) | ( n1103 & ~n1104 ) ;
  assign n1106 = ( n1042 & n1097 ) | ( n1042 & n1105 ) | ( n1097 & n1105 ) ;
  assign n1107 = ( ~n1042 & n1097 ) | ( ~n1042 & n1105 ) | ( n1097 & n1105 ) ;
  assign n1108 = ( n1042 & ~n1106 ) | ( n1042 & n1107 ) | ( ~n1106 & n1107 ) ;
  assign n1109 = ( n1083 & n1094 ) | ( n1083 & n1108 ) | ( n1094 & n1108 ) ;
  assign n1110 = ( ~n1083 & n1094 ) | ( ~n1083 & n1108 ) | ( n1094 & n1108 ) ;
  assign n1111 = ( n1083 & ~n1109 ) | ( n1083 & n1110 ) | ( ~n1109 & n1110 ) ;
  assign n1112 = ( n974 & n1017 ) | ( n974 & ~n1041 ) | ( n1017 & ~n1041 ) ;
  assign n1113 = x4 & x28 ;
  assign n1114 = x5 & x27 ;
  assign n1115 = x9 & x23 ;
  assign n1116 = ( ~n1113 & n1114 ) | ( ~n1113 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1117 = ( n1113 & n1114 ) | ( n1113 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1118 = ( n1113 & n1116 ) | ( n1113 & ~n1117 ) | ( n1116 & ~n1117 ) ;
  assign n1119 = x7 & x25 ;
  assign n1120 = x8 & x24 ;
  assign n1121 = x6 & x26 ;
  assign n1122 = ( ~n1119 & n1120 ) | ( ~n1119 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = ( n1119 & n1120 ) | ( n1119 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1124 = ( n1119 & n1122 ) | ( n1119 & ~n1123 ) | ( n1122 & ~n1123 ) ;
  assign n1125 = ( ~n1112 & n1118 ) | ( ~n1112 & n1124 ) | ( n1118 & n1124 ) ;
  assign n1126 = ( n1112 & n1118 ) | ( n1112 & n1124 ) | ( n1118 & n1124 ) ;
  assign n1127 = ( n1112 & n1125 ) | ( n1112 & ~n1126 ) | ( n1125 & ~n1126 ) ;
  assign n1128 = ( x2 & ~x30 ) | ( x2 & n355 ) | ( ~x30 & n355 ) ;
  assign n1129 = x0 & x32 ;
  assign n1130 = x2 | n355 ;
  assign n1131 = ( ~n1128 & n1129 ) | ( ~n1128 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1132 = ( n1128 & n1129 ) | ( n1128 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1133 = ( n1128 & n1131 ) | ( n1128 & ~n1132 ) | ( n1131 & ~n1132 ) ;
  assign n1134 = x11 & x21 ;
  assign n1135 = x13 & x19 ;
  assign n1136 = x12 & x20 ;
  assign n1137 = ( ~n1134 & n1135 ) | ( ~n1134 & n1136 ) | ( n1135 & n1136 ) ;
  assign n1138 = ( n1134 & n1135 ) | ( n1134 & n1136 ) | ( n1135 & n1136 ) ;
  assign n1139 = ( n1134 & n1137 ) | ( n1134 & ~n1138 ) | ( n1137 & ~n1138 ) ;
  assign n1140 = x3 & x29 ;
  assign n1141 = x14 & x18 ;
  assign n1142 = x10 & x22 ;
  assign n1143 = ( ~n1140 & n1141 ) | ( ~n1140 & n1142 ) | ( n1141 & n1142 ) ;
  assign n1144 = ( n1140 & n1141 ) | ( n1140 & n1142 ) | ( n1141 & n1142 ) ;
  assign n1145 = ( n1140 & n1143 ) | ( n1140 & ~n1144 ) | ( n1143 & ~n1144 ) ;
  assign n1146 = ( ~n1133 & n1139 ) | ( ~n1133 & n1145 ) | ( n1139 & n1145 ) ;
  assign n1147 = ( n1133 & n1139 ) | ( n1133 & n1145 ) | ( n1139 & n1145 ) ;
  assign n1148 = ( n1133 & n1146 ) | ( n1133 & ~n1147 ) | ( n1146 & ~n1147 ) ;
  assign n1149 = ( n1035 & n1127 ) | ( n1035 & n1148 ) | ( n1127 & n1148 ) ;
  assign n1150 = ( ~n1035 & n1127 ) | ( ~n1035 & n1148 ) | ( n1127 & n1148 ) ;
  assign n1151 = ( n1035 & ~n1149 ) | ( n1035 & n1150 ) | ( ~n1149 & n1150 ) ;
  assign n1152 = ( n1045 & ~n1111 ) | ( n1045 & n1151 ) | ( ~n1111 & n1151 ) ;
  assign n1153 = ( n1045 & n1111 ) | ( n1045 & n1151 ) | ( n1111 & n1151 ) ;
  assign n1154 = ( n1111 & n1152 ) | ( n1111 & ~n1153 ) | ( n1152 & ~n1153 ) ;
  assign n1155 = ( n1086 & n1090 ) | ( n1086 & n1154 ) | ( n1090 & n1154 ) ;
  assign n1156 = ( n1086 & ~n1090 ) | ( n1086 & n1154 ) | ( ~n1090 & n1154 ) ;
  assign n1157 = ( n1090 & ~n1155 ) | ( n1090 & n1156 ) | ( ~n1155 & n1156 ) ;
  assign n1158 = ( ~n1096 & n1126 ) | ( ~n1096 & n1147 ) | ( n1126 & n1147 ) ;
  assign n1159 = ( n1096 & n1126 ) | ( n1096 & n1147 ) | ( n1126 & n1147 ) ;
  assign n1160 = ( n1096 & n1158 ) | ( n1096 & ~n1159 ) | ( n1158 & ~n1159 ) ;
  assign n1161 = x5 & x28 ;
  assign n1162 = x8 & x25 ;
  assign n1163 = x6 & x27 ;
  assign n1164 = ( ~n1161 & n1162 ) | ( ~n1161 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1165 = ( n1161 & n1162 ) | ( n1161 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1166 = ( n1161 & n1164 ) | ( n1161 & ~n1165 ) | ( n1164 & ~n1165 ) ;
  assign n1167 = x16 & x17 ;
  assign n1168 = x7 & x26 ;
  assign n1169 = x15 & x18 ;
  assign n1170 = ( ~n1167 & n1168 ) | ( ~n1167 & n1169 ) | ( n1168 & n1169 ) ;
  assign n1171 = ( n1167 & n1168 ) | ( n1167 & n1169 ) | ( n1168 & n1169 ) ;
  assign n1172 = ( n1167 & n1170 ) | ( n1167 & ~n1171 ) | ( n1170 & ~n1171 ) ;
  assign n1173 = x4 & x29 ;
  assign n1174 = x3 & x30 ;
  assign n1175 = x9 & x24 ;
  assign n1176 = ( ~n1173 & n1174 ) | ( ~n1173 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1177 = ( n1173 & n1174 ) | ( n1173 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1178 = ( n1173 & n1176 ) | ( n1173 & ~n1177 ) | ( n1176 & ~n1177 ) ;
  assign n1179 = ( ~n1166 & n1172 ) | ( ~n1166 & n1178 ) | ( n1172 & n1178 ) ;
  assign n1180 = ( n1166 & n1172 ) | ( n1166 & n1178 ) | ( n1172 & n1178 ) ;
  assign n1181 = ( n1166 & n1179 ) | ( n1166 & ~n1180 ) | ( n1179 & ~n1180 ) ;
  assign n1182 = ( x2 & n355 ) | ( x2 & n1129 ) | ( n355 & n1129 ) ;
  assign n1183 = x30 & n1182 ;
  assign n1184 = ( n1138 & n1144 ) | ( n1138 & n1183 ) | ( n1144 & n1183 ) ;
  assign n1185 = ( n1138 & n1144 ) | ( n1138 & ~n1183 ) | ( n1144 & ~n1183 ) ;
  assign n1186 = ( n1183 & ~n1184 ) | ( n1183 & n1185 ) | ( ~n1184 & n1185 ) ;
  assign n1187 = x0 & x33 ;
  assign n1188 = x2 & x31 ;
  assign n1189 = x11 & x22 ;
  assign n1190 = ( ~n1187 & n1188 ) | ( ~n1187 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1191 = ( n1187 & n1188 ) | ( n1187 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1192 = ( n1187 & n1190 ) | ( n1187 & ~n1191 ) | ( n1190 & ~n1191 ) ;
  assign n1193 = ( n1117 & n1123 ) | ( n1117 & ~n1192 ) | ( n1123 & ~n1192 ) ;
  assign n1194 = ( n1117 & n1123 ) | ( n1117 & n1192 ) | ( n1123 & n1192 ) ;
  assign n1195 = ( n1192 & n1193 ) | ( n1192 & ~n1194 ) | ( n1193 & ~n1194 ) ;
  assign n1196 = ( n1181 & n1186 ) | ( n1181 & n1195 ) | ( n1186 & n1195 ) ;
  assign n1197 = ( ~n1181 & n1186 ) | ( ~n1181 & n1195 ) | ( n1186 & n1195 ) ;
  assign n1198 = ( n1181 & ~n1196 ) | ( n1181 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = ( n1149 & n1160 ) | ( n1149 & n1198 ) | ( n1160 & n1198 ) ;
  assign n1200 = ( ~n1149 & n1160 ) | ( ~n1149 & n1198 ) | ( n1160 & n1198 ) ;
  assign n1201 = ( n1149 & ~n1199 ) | ( n1149 & n1200 ) | ( ~n1199 & n1200 ) ;
  assign n1202 = ~x32 & n1100 ;
  assign n1203 = x10 & x23 ;
  assign n1204 = x15 & x31 ;
  assign n1205 = x1 & x32 ;
  assign n1206 = x17 & n1205 ;
  assign n1207 = ~n1204 & n1206 ;
  assign n1208 = x17 | n1205 ;
  assign n1209 = ~n1207 & n1208 ;
  assign n1210 = ( ~n1202 & n1203 ) | ( ~n1202 & n1209 ) | ( n1203 & n1209 ) ;
  assign n1211 = ( n1202 & n1203 ) | ( n1202 & n1209 ) | ( n1203 & n1209 ) ;
  assign n1212 = ( n1202 & n1210 ) | ( n1202 & ~n1211 ) | ( n1210 & ~n1211 ) ;
  assign n1213 = x12 & x21 ;
  assign n1214 = x13 & x20 ;
  assign n1215 = x14 & x19 ;
  assign n1216 = ( ~n1213 & n1214 ) | ( ~n1213 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1217 = ( n1213 & n1214 ) | ( n1213 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1218 = ( n1213 & n1216 ) | ( n1213 & ~n1217 ) | ( n1216 & ~n1217 ) ;
  assign n1219 = ( n1104 & ~n1212 ) | ( n1104 & n1218 ) | ( ~n1212 & n1218 ) ;
  assign n1220 = ( n1104 & n1212 ) | ( n1104 & n1218 ) | ( n1212 & n1218 ) ;
  assign n1221 = ( n1212 & n1219 ) | ( n1212 & ~n1220 ) | ( n1219 & ~n1220 ) ;
  assign n1222 = ( n1093 & ~n1106 ) | ( n1093 & n1221 ) | ( ~n1106 & n1221 ) ;
  assign n1223 = ( n1093 & n1106 ) | ( n1093 & n1221 ) | ( n1106 & n1221 ) ;
  assign n1224 = ( n1106 & n1222 ) | ( n1106 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1225 = ( n1109 & n1201 ) | ( n1109 & n1224 ) | ( n1201 & n1224 ) ;
  assign n1226 = ( n1109 & ~n1201 ) | ( n1109 & n1224 ) | ( ~n1201 & n1224 ) ;
  assign n1227 = ( n1201 & ~n1225 ) | ( n1201 & n1226 ) | ( ~n1225 & n1226 ) ;
  assign n1228 = ( n1153 & ~n1155 ) | ( n1153 & n1227 ) | ( ~n1155 & n1227 ) ;
  assign n1229 = ( n1153 & n1155 ) | ( n1153 & n1227 ) | ( n1155 & n1227 ) ;
  assign n1230 = ( n1155 & n1228 ) | ( n1155 & ~n1229 ) | ( n1228 & ~n1229 ) ;
  assign n1231 = x4 & x30 ;
  assign n1232 = x0 & x34 ;
  assign n1233 = x3 & x31 ;
  assign n1234 = ( ~n1231 & n1232 ) | ( ~n1231 & n1233 ) | ( n1232 & n1233 ) ;
  assign n1235 = ( n1231 & n1232 ) | ( n1231 & n1233 ) | ( n1232 & n1233 ) ;
  assign n1236 = ( n1231 & n1234 ) | ( n1231 & ~n1235 ) | ( n1234 & ~n1235 ) ;
  assign n1237 = ( n1184 & n1194 ) | ( n1184 & n1236 ) | ( n1194 & n1236 ) ;
  assign n1238 = ( ~n1184 & n1194 ) | ( ~n1184 & n1236 ) | ( n1194 & n1236 ) ;
  assign n1239 = ( n1184 & ~n1237 ) | ( n1184 & n1238 ) | ( ~n1237 & n1238 ) ;
  assign n1240 = ( n1159 & n1196 ) | ( n1159 & n1239 ) | ( n1196 & n1239 ) ;
  assign n1241 = ( n1159 & n1196 ) | ( n1159 & ~n1239 ) | ( n1196 & ~n1239 ) ;
  assign n1242 = ( n1239 & ~n1240 ) | ( n1239 & n1241 ) | ( ~n1240 & n1241 ) ;
  assign n1243 = x11 & x23 ;
  assign n1244 = x2 & x32 ;
  assign n1245 = x12 & x22 ;
  assign n1246 = ( ~n1243 & n1244 ) | ( ~n1243 & n1245 ) | ( n1244 & n1245 ) ;
  assign n1247 = ( n1243 & n1244 ) | ( n1243 & n1245 ) | ( n1244 & n1245 ) ;
  assign n1248 = ( n1243 & n1246 ) | ( n1243 & ~n1247 ) | ( n1246 & ~n1247 ) ;
  assign n1249 = ( n1211 & n1217 ) | ( n1211 & n1248 ) | ( n1217 & n1248 ) ;
  assign n1250 = ( ~n1211 & n1217 ) | ( ~n1211 & n1248 ) | ( n1217 & n1248 ) ;
  assign n1251 = ( n1211 & ~n1249 ) | ( n1211 & n1250 ) | ( ~n1249 & n1250 ) ;
  assign n1252 = x5 & x29 ;
  assign n1253 = x10 & x24 ;
  assign n1254 = x9 & x25 ;
  assign n1255 = ( ~n1252 & n1253 ) | ( ~n1252 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1256 = ( n1252 & n1253 ) | ( n1252 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1257 = ( n1252 & n1255 ) | ( n1252 & ~n1256 ) | ( n1255 & ~n1256 ) ;
  assign n1258 = x14 & x20 ;
  assign n1259 = x13 & x21 ;
  assign n1260 = x15 & x19 ;
  assign n1261 = ( ~n1258 & n1259 ) | ( ~n1258 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1262 = ( n1258 & n1259 ) | ( n1258 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1263 = ( n1258 & n1261 ) | ( n1258 & ~n1262 ) | ( n1261 & ~n1262 ) ;
  assign n1264 = x7 & x27 ;
  assign n1265 = x6 & x28 ;
  assign n1266 = x8 & x26 ;
  assign n1267 = ( ~n1264 & n1265 ) | ( ~n1264 & n1266 ) | ( n1265 & n1266 ) ;
  assign n1268 = ( n1264 & n1265 ) | ( n1264 & n1266 ) | ( n1265 & n1266 ) ;
  assign n1269 = ( n1264 & n1267 ) | ( n1264 & ~n1268 ) | ( n1267 & ~n1268 ) ;
  assign n1270 = ( ~n1257 & n1263 ) | ( ~n1257 & n1269 ) | ( n1263 & n1269 ) ;
  assign n1271 = ( n1257 & n1263 ) | ( n1257 & n1269 ) | ( n1263 & n1269 ) ;
  assign n1272 = ( n1257 & n1270 ) | ( n1257 & ~n1271 ) | ( n1270 & ~n1271 ) ;
  assign n1273 = ( n1220 & n1251 ) | ( n1220 & n1272 ) | ( n1251 & n1272 ) ;
  assign n1274 = ( ~n1220 & n1251 ) | ( ~n1220 & n1272 ) | ( n1251 & n1272 ) ;
  assign n1275 = ( n1220 & ~n1273 ) | ( n1220 & n1274 ) | ( ~n1273 & n1274 ) ;
  assign n1276 = x16 & x18 ;
  assign n1277 = x1 & x33 ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = x18 & x33 ;
  assign n1280 = n355 & n1279 ;
  assign n1281 = n1278 & ~n1280 ;
  assign n1282 = ( n1171 & n1206 ) | ( n1171 & n1281 ) | ( n1206 & n1281 ) ;
  assign n1283 = ( n1171 & ~n1206 ) | ( n1171 & n1281 ) | ( ~n1206 & n1281 ) ;
  assign n1284 = ( n1206 & ~n1282 ) | ( n1206 & n1283 ) | ( ~n1282 & n1283 ) ;
  assign n1285 = ( ~n1165 & n1177 ) | ( ~n1165 & n1191 ) | ( n1177 & n1191 ) ;
  assign n1286 = ( n1165 & n1177 ) | ( n1165 & n1191 ) | ( n1177 & n1191 ) ;
  assign n1287 = ( n1165 & n1285 ) | ( n1165 & ~n1286 ) | ( n1285 & ~n1286 ) ;
  assign n1288 = ( n1180 & n1284 ) | ( n1180 & n1287 ) | ( n1284 & n1287 ) ;
  assign n1289 = ( ~n1180 & n1284 ) | ( ~n1180 & n1287 ) | ( n1284 & n1287 ) ;
  assign n1290 = ( n1180 & ~n1288 ) | ( n1180 & n1289 ) | ( ~n1288 & n1289 ) ;
  assign n1291 = ( n1223 & ~n1275 ) | ( n1223 & n1290 ) | ( ~n1275 & n1290 ) ;
  assign n1292 = ( n1223 & n1275 ) | ( n1223 & n1290 ) | ( n1275 & n1290 ) ;
  assign n1293 = ( n1275 & n1291 ) | ( n1275 & ~n1292 ) | ( n1291 & ~n1292 ) ;
  assign n1294 = ( n1199 & n1242 ) | ( n1199 & n1293 ) | ( n1242 & n1293 ) ;
  assign n1295 = ( n1199 & ~n1242 ) | ( n1199 & n1293 ) | ( ~n1242 & n1293 ) ;
  assign n1296 = ( n1242 & ~n1294 ) | ( n1242 & n1295 ) | ( ~n1294 & n1295 ) ;
  assign n1297 = ( n1225 & n1229 ) | ( n1225 & n1296 ) | ( n1229 & n1296 ) ;
  assign n1298 = ( n1225 & ~n1229 ) | ( n1225 & n1296 ) | ( ~n1229 & n1296 ) ;
  assign n1299 = ( n1229 & ~n1297 ) | ( n1229 & n1298 ) | ( ~n1297 & n1298 ) ;
  assign n1300 = x2 & x33 ;
  assign n1301 = x0 & x35 ;
  assign n1302 = ( ~n1280 & n1300 ) | ( ~n1280 & n1301 ) | ( n1300 & n1301 ) ;
  assign n1303 = ( n1280 & n1300 ) | ( n1280 & n1301 ) | ( n1300 & n1301 ) ;
  assign n1304 = ( n1280 & n1302 ) | ( n1280 & ~n1303 ) | ( n1302 & ~n1303 ) ;
  assign n1305 = x12 & x23 ;
  assign n1306 = x3 & x32 ;
  assign n1307 = x11 & x24 ;
  assign n1308 = ( ~n1305 & n1306 ) | ( ~n1305 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1309 = ( n1305 & n1306 ) | ( n1305 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1310 = ( n1305 & n1308 ) | ( n1305 & ~n1309 ) | ( n1308 & ~n1309 ) ;
  assign n1311 = x13 & x22 ;
  assign n1312 = x14 & x21 ;
  assign n1313 = x15 & x20 ;
  assign n1314 = ( ~n1311 & n1312 ) | ( ~n1311 & n1313 ) | ( n1312 & n1313 ) ;
  assign n1315 = ( n1311 & n1312 ) | ( n1311 & n1313 ) | ( n1312 & n1313 ) ;
  assign n1316 = ( n1311 & n1314 ) | ( n1311 & ~n1315 ) | ( n1314 & ~n1315 ) ;
  assign n1317 = ( ~n1304 & n1310 ) | ( ~n1304 & n1316 ) | ( n1310 & n1316 ) ;
  assign n1318 = ( n1304 & n1310 ) | ( n1304 & n1316 ) | ( n1310 & n1316 ) ;
  assign n1319 = ( n1304 & n1317 ) | ( n1304 & ~n1318 ) | ( n1317 & ~n1318 ) ;
  assign n1320 = x8 & x27 ;
  assign n1321 = x6 & x29 ;
  assign n1322 = x5 & x30 ;
  assign n1323 = ( ~n1320 & n1321 ) | ( ~n1320 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1324 = ( n1320 & n1321 ) | ( n1320 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1325 = ( n1320 & n1323 ) | ( n1320 & ~n1324 ) | ( n1323 & ~n1324 ) ;
  assign n1326 = x9 & x26 ;
  assign n1327 = x10 & x25 ;
  assign n1328 = x4 & x31 ;
  assign n1329 = ( ~n1326 & n1327 ) | ( ~n1326 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = ( n1326 & n1327 ) | ( n1326 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1331 = ( n1326 & n1329 ) | ( n1326 & ~n1330 ) | ( n1329 & ~n1330 ) ;
  assign n1332 = x16 & x19 ;
  assign n1333 = x17 & x18 ;
  assign n1334 = x7 & x28 ;
  assign n1335 = ( ~n1332 & n1333 ) | ( ~n1332 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1336 = ( n1332 & n1333 ) | ( n1332 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1337 = ( n1332 & n1335 ) | ( n1332 & ~n1336 ) | ( n1335 & ~n1336 ) ;
  assign n1338 = ( ~n1325 & n1331 ) | ( ~n1325 & n1337 ) | ( n1331 & n1337 ) ;
  assign n1339 = ( n1325 & n1331 ) | ( n1325 & n1337 ) | ( n1331 & n1337 ) ;
  assign n1340 = ( n1325 & n1338 ) | ( n1325 & ~n1339 ) | ( n1338 & ~n1339 ) ;
  assign n1341 = ( n1237 & n1319 ) | ( n1237 & n1340 ) | ( n1319 & n1340 ) ;
  assign n1342 = ( ~n1237 & n1319 ) | ( ~n1237 & n1340 ) | ( n1319 & n1340 ) ;
  assign n1343 = ( n1237 & ~n1341 ) | ( n1237 & n1342 ) | ( ~n1341 & n1342 ) ;
  assign n1344 = ( ~n1235 & n1247 ) | ( ~n1235 & n1262 ) | ( n1247 & n1262 ) ;
  assign n1345 = ( n1235 & n1247 ) | ( n1235 & n1262 ) | ( n1247 & n1262 ) ;
  assign n1346 = ( n1235 & n1344 ) | ( n1235 & ~n1345 ) | ( n1344 & ~n1345 ) ;
  assign n1347 = ~x1 & x18 ;
  assign n1348 = ( x1 & x18 ) | ( x1 & x34 ) | ( x18 & x34 ) ;
  assign n1349 = x18 & x34 ;
  assign n1350 = ( n1347 & n1348 ) | ( n1347 & ~n1349 ) | ( n1348 & ~n1349 ) ;
  assign n1351 = ( n1256 & n1268 ) | ( n1256 & n1350 ) | ( n1268 & n1350 ) ;
  assign n1352 = ( ~n1256 & n1268 ) | ( ~n1256 & n1350 ) | ( n1268 & n1350 ) ;
  assign n1353 = ( n1256 & ~n1351 ) | ( n1256 & n1352 ) | ( ~n1351 & n1352 ) ;
  assign n1354 = ( n1271 & n1346 ) | ( n1271 & n1353 ) | ( n1346 & n1353 ) ;
  assign n1355 = ( ~n1271 & n1346 ) | ( ~n1271 & n1353 ) | ( n1346 & n1353 ) ;
  assign n1356 = ( n1271 & ~n1354 ) | ( n1271 & n1355 ) | ( ~n1354 & n1355 ) ;
  assign n1357 = ( n1240 & n1343 ) | ( n1240 & n1356 ) | ( n1343 & n1356 ) ;
  assign n1358 = ( ~n1240 & n1343 ) | ( ~n1240 & n1356 ) | ( n1343 & n1356 ) ;
  assign n1359 = ( n1240 & ~n1357 ) | ( n1240 & n1358 ) | ( ~n1357 & n1358 ) ;
  assign n1360 = ( n1249 & ~n1282 ) | ( n1249 & n1286 ) | ( ~n1282 & n1286 ) ;
  assign n1361 = ( n1249 & n1282 ) | ( n1249 & n1286 ) | ( n1282 & n1286 ) ;
  assign n1362 = ( n1282 & n1360 ) | ( n1282 & ~n1361 ) | ( n1360 & ~n1361 ) ;
  assign n1363 = ( n1273 & n1288 ) | ( n1273 & n1362 ) | ( n1288 & n1362 ) ;
  assign n1364 = ( n1273 & n1288 ) | ( n1273 & ~n1362 ) | ( n1288 & ~n1362 ) ;
  assign n1365 = ( n1362 & ~n1363 ) | ( n1362 & n1364 ) | ( ~n1363 & n1364 ) ;
  assign n1366 = ( n1292 & n1359 ) | ( n1292 & n1365 ) | ( n1359 & n1365 ) ;
  assign n1367 = ( n1292 & ~n1359 ) | ( n1292 & n1365 ) | ( ~n1359 & n1365 ) ;
  assign n1368 = ( n1359 & ~n1366 ) | ( n1359 & n1367 ) | ( ~n1366 & n1367 ) ;
  assign n1369 = ( n1294 & n1297 ) | ( n1294 & n1368 ) | ( n1297 & n1368 ) ;
  assign n1370 = ( n1294 & ~n1297 ) | ( n1294 & n1368 ) | ( ~n1297 & n1368 ) ;
  assign n1371 = ( n1297 & ~n1369 ) | ( n1297 & n1370 ) | ( ~n1369 & n1370 ) ;
  assign n1372 = x17 & x35 ;
  assign n1373 = n481 & n1372 ;
  assign n1374 = ( ~x1 & x35 ) | ( ~x1 & n1373 ) | ( x35 & n1373 ) ;
  assign n1375 = x19 & ~n1373 ;
  assign n1376 = x17 & n1375 ;
  assign n1377 = ( x35 & ~n1374 ) | ( x35 & n1376 ) | ( ~n1374 & n1376 ) ;
  assign n1378 = x1 & n1349 ;
  assign n1379 = x0 & x36 ;
  assign n1380 = ( n1377 & n1378 ) | ( n1377 & n1379 ) | ( n1378 & n1379 ) ;
  assign n1381 = ( ~n1377 & n1378 ) | ( ~n1377 & n1379 ) | ( n1378 & n1379 ) ;
  assign n1382 = ( n1377 & ~n1380 ) | ( n1377 & n1381 ) | ( ~n1380 & n1381 ) ;
  assign n1383 = x16 & x20 ;
  assign n1384 = x15 & x21 ;
  assign n1385 = x14 & x22 ;
  assign n1386 = ( ~n1383 & n1384 ) | ( ~n1383 & n1385 ) | ( n1384 & n1385 ) ;
  assign n1387 = ( n1383 & n1384 ) | ( n1383 & n1385 ) | ( n1384 & n1385 ) ;
  assign n1388 = ( n1383 & n1386 ) | ( n1383 & ~n1387 ) | ( n1386 & ~n1387 ) ;
  assign n1389 = x4 & x32 ;
  assign n1390 = x3 & x33 ;
  assign n1391 = x11 & x25 ;
  assign n1392 = ( ~n1389 & n1390 ) | ( ~n1389 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = ( n1389 & n1390 ) | ( n1389 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1394 = ( n1389 & n1392 ) | ( n1389 & ~n1393 ) | ( n1392 & ~n1393 ) ;
  assign n1395 = ( n1382 & n1388 ) | ( n1382 & n1394 ) | ( n1388 & n1394 ) ;
  assign n1396 = ( ~n1382 & n1388 ) | ( ~n1382 & n1394 ) | ( n1388 & n1394 ) ;
  assign n1397 = ( n1382 & ~n1395 ) | ( n1382 & n1396 ) | ( ~n1395 & n1396 ) ;
  assign n1398 = x7 & x29 ;
  assign n1399 = x8 & x28 ;
  assign n1400 = x6 & x30 ;
  assign n1401 = ( ~n1398 & n1399 ) | ( ~n1398 & n1400 ) | ( n1399 & n1400 ) ;
  assign n1402 = ( n1398 & n1399 ) | ( n1398 & n1400 ) | ( n1399 & n1400 ) ;
  assign n1403 = ( n1398 & n1401 ) | ( n1398 & ~n1402 ) | ( n1401 & ~n1402 ) ;
  assign n1404 = x2 & x34 ;
  assign n1405 = x12 & x24 ;
  assign n1406 = x13 & x23 ;
  assign n1407 = ( ~n1404 & n1405 ) | ( ~n1404 & n1406 ) | ( n1405 & n1406 ) ;
  assign n1408 = ( n1404 & n1405 ) | ( n1404 & n1406 ) | ( n1405 & n1406 ) ;
  assign n1409 = ( n1404 & n1407 ) | ( n1404 & ~n1408 ) | ( n1407 & ~n1408 ) ;
  assign n1410 = x9 & x27 ;
  assign n1411 = x10 & x26 ;
  assign n1412 = x5 & x31 ;
  assign n1413 = ( ~n1410 & n1411 ) | ( ~n1410 & n1412 ) | ( n1411 & n1412 ) ;
  assign n1414 = ( n1410 & n1411 ) | ( n1410 & n1412 ) | ( n1411 & n1412 ) ;
  assign n1415 = ( n1410 & n1413 ) | ( n1410 & ~n1414 ) | ( n1413 & ~n1414 ) ;
  assign n1416 = ( ~n1403 & n1409 ) | ( ~n1403 & n1415 ) | ( n1409 & n1415 ) ;
  assign n1417 = ( n1403 & n1409 ) | ( n1403 & n1415 ) | ( n1409 & n1415 ) ;
  assign n1418 = ( n1403 & n1416 ) | ( n1403 & ~n1417 ) | ( n1416 & ~n1417 ) ;
  assign n1419 = ( n1361 & n1397 ) | ( n1361 & n1418 ) | ( n1397 & n1418 ) ;
  assign n1420 = ( n1361 & ~n1397 ) | ( n1361 & n1418 ) | ( ~n1397 & n1418 ) ;
  assign n1421 = ( n1397 & ~n1419 ) | ( n1397 & n1420 ) | ( ~n1419 & n1420 ) ;
  assign n1422 = ( ~n1303 & n1309 ) | ( ~n1303 & n1315 ) | ( n1309 & n1315 ) ;
  assign n1423 = ( n1303 & n1309 ) | ( n1303 & n1315 ) | ( n1309 & n1315 ) ;
  assign n1424 = ( n1303 & n1422 ) | ( n1303 & ~n1423 ) | ( n1422 & ~n1423 ) ;
  assign n1425 = ( n1324 & ~n1330 ) | ( n1324 & n1336 ) | ( ~n1330 & n1336 ) ;
  assign n1426 = ( n1324 & n1330 ) | ( n1324 & n1336 ) | ( n1330 & n1336 ) ;
  assign n1427 = ( n1330 & n1425 ) | ( n1330 & ~n1426 ) | ( n1425 & ~n1426 ) ;
  assign n1428 = ( n1339 & n1424 ) | ( n1339 & n1427 ) | ( n1424 & n1427 ) ;
  assign n1429 = ( n1339 & ~n1424 ) | ( n1339 & n1427 ) | ( ~n1424 & n1427 ) ;
  assign n1430 = ( n1424 & ~n1428 ) | ( n1424 & n1429 ) | ( ~n1428 & n1429 ) ;
  assign n1431 = ( n1363 & n1421 ) | ( n1363 & n1430 ) | ( n1421 & n1430 ) ;
  assign n1432 = ( n1363 & ~n1421 ) | ( n1363 & n1430 ) | ( ~n1421 & n1430 ) ;
  assign n1433 = ( n1421 & ~n1431 ) | ( n1421 & n1432 ) | ( ~n1431 & n1432 ) ;
  assign n1434 = ( n1318 & n1345 ) | ( n1318 & ~n1351 ) | ( n1345 & ~n1351 ) ;
  assign n1435 = ( n1318 & n1345 ) | ( n1318 & n1351 ) | ( n1345 & n1351 ) ;
  assign n1436 = ( n1351 & n1434 ) | ( n1351 & ~n1435 ) | ( n1434 & ~n1435 ) ;
  assign n1437 = ( n1341 & n1354 ) | ( n1341 & n1436 ) | ( n1354 & n1436 ) ;
  assign n1438 = ( ~n1341 & n1354 ) | ( ~n1341 & n1436 ) | ( n1354 & n1436 ) ;
  assign n1439 = ( n1341 & ~n1437 ) | ( n1341 & n1438 ) | ( ~n1437 & n1438 ) ;
  assign n1440 = ( n1357 & n1433 ) | ( n1357 & n1439 ) | ( n1433 & n1439 ) ;
  assign n1441 = ( ~n1357 & n1433 ) | ( ~n1357 & n1439 ) | ( n1433 & n1439 ) ;
  assign n1442 = ( n1357 & ~n1440 ) | ( n1357 & n1441 ) | ( ~n1440 & n1441 ) ;
  assign n1443 = ( n1366 & ~n1369 ) | ( n1366 & n1442 ) | ( ~n1369 & n1442 ) ;
  assign n1444 = ( n1366 & n1369 ) | ( n1366 & n1442 ) | ( n1369 & n1442 ) ;
  assign n1445 = ( n1369 & n1443 ) | ( n1369 & ~n1444 ) | ( n1443 & ~n1444 ) ;
  assign n1446 = x10 & x27 ;
  assign n1447 = x11 & x26 ;
  assign n1448 = x5 & x32 ;
  assign n1449 = ( ~n1446 & n1447 ) | ( ~n1446 & n1448 ) | ( n1447 & n1448 ) ;
  assign n1450 = ( n1446 & n1447 ) | ( n1446 & n1448 ) | ( n1447 & n1448 ) ;
  assign n1451 = ( n1446 & n1449 ) | ( n1446 & ~n1450 ) | ( n1449 & ~n1450 ) ;
  assign n1452 = x18 & x19 ;
  assign n1453 = x17 & x20 ;
  assign n1454 = x8 & x29 ;
  assign n1455 = ( ~n1452 & n1453 ) | ( ~n1452 & n1454 ) | ( n1453 & n1454 ) ;
  assign n1456 = ( n1452 & n1453 ) | ( n1452 & n1454 ) | ( n1453 & n1454 ) ;
  assign n1457 = ( n1452 & n1455 ) | ( n1452 & ~n1456 ) | ( n1455 & ~n1456 ) ;
  assign n1458 = ( ~n1423 & n1451 ) | ( ~n1423 & n1457 ) | ( n1451 & n1457 ) ;
  assign n1459 = ( n1423 & n1451 ) | ( n1423 & n1457 ) | ( n1451 & n1457 ) ;
  assign n1460 = ( n1423 & n1458 ) | ( n1423 & ~n1459 ) | ( n1458 & ~n1459 ) ;
  assign n1461 = x4 & x33 ;
  assign n1462 = x0 & x37 ;
  assign n1463 = x12 & x25 ;
  assign n1464 = ( ~n1461 & n1462 ) | ( ~n1461 & n1463 ) | ( n1462 & n1463 ) ;
  assign n1465 = ( n1461 & n1462 ) | ( n1461 & n1463 ) | ( n1462 & n1463 ) ;
  assign n1466 = ( n1461 & n1464 ) | ( n1461 & ~n1465 ) | ( n1464 & ~n1465 ) ;
  assign n1467 = x9 & x28 ;
  assign n1468 = x6 & x31 ;
  assign n1469 = x7 & x30 ;
  assign n1470 = ( ~n1467 & n1468 ) | ( ~n1467 & n1469 ) | ( n1468 & n1469 ) ;
  assign n1471 = ( n1467 & n1468 ) | ( n1467 & n1469 ) | ( n1468 & n1469 ) ;
  assign n1472 = ( n1467 & n1470 ) | ( n1467 & ~n1471 ) | ( n1470 & ~n1471 ) ;
  assign n1473 = x16 & x21 ;
  assign n1474 = x3 & x34 ;
  assign n1475 = x2 & x35 ;
  assign n1476 = ( ~n1473 & n1474 ) | ( ~n1473 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1477 = ( n1473 & n1474 ) | ( n1473 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1478 = ( n1473 & n1476 ) | ( n1473 & ~n1477 ) | ( n1476 & ~n1477 ) ;
  assign n1479 = ( ~n1466 & n1472 ) | ( ~n1466 & n1478 ) | ( n1472 & n1478 ) ;
  assign n1480 = ( n1466 & n1472 ) | ( n1466 & n1478 ) | ( n1472 & n1478 ) ;
  assign n1481 = ( n1466 & n1479 ) | ( n1466 & ~n1480 ) | ( n1479 & ~n1480 ) ;
  assign n1482 = ( n1435 & n1460 ) | ( n1435 & n1481 ) | ( n1460 & n1481 ) ;
  assign n1483 = ( ~n1435 & n1460 ) | ( ~n1435 & n1481 ) | ( n1460 & n1481 ) ;
  assign n1484 = ( n1435 & ~n1482 ) | ( n1435 & n1483 ) | ( ~n1482 & n1483 ) ;
  assign n1485 = x13 & x24 ;
  assign n1486 = x15 & x22 ;
  assign n1487 = x14 & x23 ;
  assign n1488 = ( ~n1485 & n1486 ) | ( ~n1485 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1489 = ( n1485 & n1486 ) | ( n1485 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1490 = ( n1485 & n1488 ) | ( n1485 & ~n1489 ) | ( n1488 & ~n1489 ) ;
  assign n1491 = ( ~n1380 & n1414 ) | ( ~n1380 & n1490 ) | ( n1414 & n1490 ) ;
  assign n1492 = ( n1380 & n1414 ) | ( n1380 & n1490 ) | ( n1414 & n1490 ) ;
  assign n1493 = ( n1380 & n1491 ) | ( n1380 & ~n1492 ) | ( n1491 & ~n1492 ) ;
  assign n1494 = ( n1387 & n1393 ) | ( n1387 & ~n1408 ) | ( n1393 & ~n1408 ) ;
  assign n1495 = ( n1387 & n1393 ) | ( n1387 & n1408 ) | ( n1393 & n1408 ) ;
  assign n1496 = ( n1408 & n1494 ) | ( n1408 & ~n1495 ) | ( n1494 & ~n1495 ) ;
  assign n1497 = ( n1395 & n1493 ) | ( n1395 & n1496 ) | ( n1493 & n1496 ) ;
  assign n1498 = ( ~n1395 & n1493 ) | ( ~n1395 & n1496 ) | ( n1493 & n1496 ) ;
  assign n1499 = ( n1395 & ~n1497 ) | ( n1395 & n1498 ) | ( ~n1497 & n1498 ) ;
  assign n1500 = ( n1437 & n1484 ) | ( n1437 & n1499 ) | ( n1484 & n1499 ) ;
  assign n1501 = ( ~n1437 & n1484 ) | ( ~n1437 & n1499 ) | ( n1484 & n1499 ) ;
  assign n1502 = ( n1437 & ~n1500 ) | ( n1437 & n1501 ) | ( ~n1500 & n1501 ) ;
  assign n1503 = x1 & x36 ;
  assign n1504 = ( n1375 & n1402 ) | ( n1375 & ~n1503 ) | ( n1402 & ~n1503 ) ;
  assign n1505 = ( n1375 & ~n1402 ) | ( n1375 & n1503 ) | ( ~n1402 & n1503 ) ;
  assign n1506 = ( ~n1375 & n1504 ) | ( ~n1375 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1507 = ( n1417 & n1426 ) | ( n1417 & ~n1506 ) | ( n1426 & ~n1506 ) ;
  assign n1508 = ( n1417 & n1426 ) | ( n1417 & n1506 ) | ( n1426 & n1506 ) ;
  assign n1509 = ( n1506 & n1507 ) | ( n1506 & ~n1508 ) | ( n1507 & ~n1508 ) ;
  assign n1510 = ( n1419 & n1428 ) | ( n1419 & n1509 ) | ( n1428 & n1509 ) ;
  assign n1511 = ( ~n1419 & n1428 ) | ( ~n1419 & n1509 ) | ( n1428 & n1509 ) ;
  assign n1512 = ( n1419 & ~n1510 ) | ( n1419 & n1511 ) | ( ~n1510 & n1511 ) ;
  assign n1513 = ( n1431 & n1502 ) | ( n1431 & n1512 ) | ( n1502 & n1512 ) ;
  assign n1514 = ( n1431 & ~n1502 ) | ( n1431 & n1512 ) | ( ~n1502 & n1512 ) ;
  assign n1515 = ( n1502 & ~n1513 ) | ( n1502 & n1514 ) | ( ~n1513 & n1514 ) ;
  assign n1516 = ( n1440 & ~n1444 ) | ( n1440 & n1515 ) | ( ~n1444 & n1515 ) ;
  assign n1517 = ( n1440 & n1444 ) | ( n1440 & n1515 ) | ( n1444 & n1515 ) ;
  assign n1518 = ( n1444 & n1516 ) | ( n1444 & ~n1517 ) | ( n1516 & ~n1517 ) ;
  assign n1519 = ( n1465 & n1477 ) | ( n1465 & ~n1489 ) | ( n1477 & ~n1489 ) ;
  assign n1520 = ( n1465 & n1477 ) | ( n1465 & n1489 ) | ( n1477 & n1489 ) ;
  assign n1521 = ( n1489 & n1519 ) | ( n1489 & ~n1520 ) | ( n1519 & ~n1520 ) ;
  assign n1522 = x17 & x21 ;
  assign n1523 = x16 & x22 ;
  assign n1524 = x15 & x23 ;
  assign n1525 = ( ~n1522 & n1523 ) | ( ~n1522 & n1524 ) | ( n1523 & n1524 ) ;
  assign n1526 = ( n1522 & n1523 ) | ( n1522 & n1524 ) | ( n1523 & n1524 ) ;
  assign n1527 = ( n1522 & n1525 ) | ( n1522 & ~n1526 ) | ( n1525 & ~n1526 ) ;
  assign n1528 = x7 & x31 ;
  assign n1529 = x8 & x30 ;
  assign n1530 = x9 & x29 ;
  assign n1531 = ( ~n1528 & n1529 ) | ( ~n1528 & n1530 ) | ( n1529 & n1530 ) ;
  assign n1532 = ( n1528 & n1529 ) | ( n1528 & n1530 ) | ( n1529 & n1530 ) ;
  assign n1533 = ( n1528 & n1531 ) | ( n1528 & ~n1532 ) | ( n1531 & ~n1532 ) ;
  assign n1534 = x10 & x28 ;
  assign n1535 = x5 & x33 ;
  assign n1536 = x6 & x32 ;
  assign n1537 = ( ~n1534 & n1535 ) | ( ~n1534 & n1536 ) | ( n1535 & n1536 ) ;
  assign n1538 = ( n1534 & n1535 ) | ( n1534 & n1536 ) | ( n1535 & n1536 ) ;
  assign n1539 = ( n1534 & n1537 ) | ( n1534 & ~n1538 ) | ( n1537 & ~n1538 ) ;
  assign n1540 = ( ~n1527 & n1533 ) | ( ~n1527 & n1539 ) | ( n1533 & n1539 ) ;
  assign n1541 = ( n1527 & n1533 ) | ( n1527 & n1539 ) | ( n1533 & n1539 ) ;
  assign n1542 = ( n1527 & n1540 ) | ( n1527 & ~n1541 ) | ( n1540 & ~n1541 ) ;
  assign n1543 = ( n1459 & n1521 ) | ( n1459 & n1542 ) | ( n1521 & n1542 ) ;
  assign n1544 = ( ~n1459 & n1521 ) | ( ~n1459 & n1542 ) | ( n1521 & n1542 ) ;
  assign n1545 = ( n1459 & ~n1543 ) | ( n1459 & n1544 ) | ( ~n1543 & n1544 ) ;
  assign n1546 = ( ~n1482 & n1497 ) | ( ~n1482 & n1545 ) | ( n1497 & n1545 ) ;
  assign n1547 = ( n1482 & n1497 ) | ( n1482 & n1545 ) | ( n1497 & n1545 ) ;
  assign n1548 = ( n1482 & n1546 ) | ( n1482 & ~n1547 ) | ( n1546 & ~n1547 ) ;
  assign n1549 = ( n1373 & n1402 ) | ( n1373 & ~n1506 ) | ( n1402 & ~n1506 ) ;
  assign n1550 = x4 & x34 ;
  assign n1551 = x12 & x26 ;
  assign n1552 = x11 & x27 ;
  assign n1553 = ( ~n1550 & n1551 ) | ( ~n1550 & n1552 ) | ( n1551 & n1552 ) ;
  assign n1554 = ( n1550 & n1551 ) | ( n1550 & n1552 ) | ( n1551 & n1552 ) ;
  assign n1555 = ( n1550 & n1553 ) | ( n1550 & ~n1554 ) | ( n1553 & ~n1554 ) ;
  assign n1556 = ( n1495 & ~n1549 ) | ( n1495 & n1555 ) | ( ~n1549 & n1555 ) ;
  assign n1557 = ( n1495 & n1549 ) | ( n1495 & n1555 ) | ( n1549 & n1555 ) ;
  assign n1558 = ( n1549 & n1556 ) | ( n1549 & ~n1557 ) | ( n1556 & ~n1557 ) ;
  assign n1559 = ( x2 & ~x36 ) | ( x2 & n481 ) | ( ~x36 & n481 ) ;
  assign n1560 = x0 & x38 ;
  assign n1561 = x2 | n481 ;
  assign n1562 = ( ~n1559 & n1560 ) | ( ~n1559 & n1561 ) | ( n1560 & n1561 ) ;
  assign n1563 = ( n1559 & n1560 ) | ( n1559 & n1561 ) | ( n1560 & n1561 ) ;
  assign n1564 = ( n1559 & n1562 ) | ( n1559 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n1565 = x3 & x35 ;
  assign n1566 = x13 & x25 ;
  assign n1567 = x14 & x24 ;
  assign n1568 = ( ~n1565 & n1566 ) | ( ~n1565 & n1567 ) | ( n1566 & n1567 ) ;
  assign n1569 = ( n1565 & n1566 ) | ( n1565 & n1567 ) | ( n1566 & n1567 ) ;
  assign n1570 = ( n1565 & n1568 ) | ( n1565 & ~n1569 ) | ( n1568 & ~n1569 ) ;
  assign n1571 = ( n1450 & ~n1564 ) | ( n1450 & n1570 ) | ( ~n1564 & n1570 ) ;
  assign n1572 = ( n1450 & n1564 ) | ( n1450 & n1570 ) | ( n1564 & n1570 ) ;
  assign n1573 = ( n1564 & n1571 ) | ( n1564 & ~n1572 ) | ( n1571 & ~n1572 ) ;
  assign n1574 = ( n1508 & n1558 ) | ( n1508 & n1573 ) | ( n1558 & n1573 ) ;
  assign n1575 = ( n1508 & ~n1558 ) | ( n1508 & n1573 ) | ( ~n1558 & n1573 ) ;
  assign n1576 = ( n1558 & ~n1574 ) | ( n1558 & n1575 ) | ( ~n1574 & n1575 ) ;
  assign n1577 = x18 & x20 ;
  assign n1578 = x1 & x37 ;
  assign n1579 = n1577 | n1578 ;
  assign n1580 = x18 & x37 ;
  assign n1581 = n534 & n1580 ;
  assign n1582 = n1579 & ~n1581 ;
  assign n1583 = ( n1456 & n1471 ) | ( n1456 & ~n1582 ) | ( n1471 & ~n1582 ) ;
  assign n1584 = ( n1456 & n1471 ) | ( n1456 & n1582 ) | ( n1471 & n1582 ) ;
  assign n1585 = ( n1582 & n1583 ) | ( n1582 & ~n1584 ) | ( n1583 & ~n1584 ) ;
  assign n1586 = ( n1480 & n1492 ) | ( n1480 & ~n1585 ) | ( n1492 & ~n1585 ) ;
  assign n1587 = ( n1480 & n1492 ) | ( n1480 & n1585 ) | ( n1492 & n1585 ) ;
  assign n1588 = ( n1585 & n1586 ) | ( n1585 & ~n1587 ) | ( n1586 & ~n1587 ) ;
  assign n1589 = ( n1510 & n1576 ) | ( n1510 & n1588 ) | ( n1576 & n1588 ) ;
  assign n1590 = ( n1510 & ~n1576 ) | ( n1510 & n1588 ) | ( ~n1576 & n1588 ) ;
  assign n1591 = ( n1576 & ~n1589 ) | ( n1576 & n1590 ) | ( ~n1589 & n1590 ) ;
  assign n1592 = ( ~n1500 & n1548 ) | ( ~n1500 & n1591 ) | ( n1548 & n1591 ) ;
  assign n1593 = ( n1500 & n1548 ) | ( n1500 & n1591 ) | ( n1548 & n1591 ) ;
  assign n1594 = ( n1500 & n1592 ) | ( n1500 & ~n1593 ) | ( n1592 & ~n1593 ) ;
  assign n1595 = ( n1513 & n1517 ) | ( n1513 & n1594 ) | ( n1517 & n1594 ) ;
  assign n1596 = ( n1513 & n1517 ) | ( n1513 & ~n1594 ) | ( n1517 & ~n1594 ) ;
  assign n1597 = ( n1594 & ~n1595 ) | ( n1594 & n1596 ) | ( ~n1595 & n1596 ) ;
  assign n1598 = ( x2 & n481 ) | ( x2 & n1560 ) | ( n481 & n1560 ) ;
  assign n1599 = x36 & n1598 ;
  assign n1600 = ( n1526 & n1569 ) | ( n1526 & n1599 ) | ( n1569 & n1599 ) ;
  assign n1601 = ( n1526 & n1569 ) | ( n1526 & ~n1599 ) | ( n1569 & ~n1599 ) ;
  assign n1602 = ( n1599 & ~n1600 ) | ( n1599 & n1601 ) | ( ~n1600 & n1601 ) ;
  assign n1603 = ( n1541 & ~n1572 ) | ( n1541 & n1602 ) | ( ~n1572 & n1602 ) ;
  assign n1604 = ( n1541 & n1572 ) | ( n1541 & n1602 ) | ( n1572 & n1602 ) ;
  assign n1605 = ( n1572 & n1603 ) | ( n1572 & ~n1604 ) | ( n1603 & ~n1604 ) ;
  assign n1606 = x20 & ~n1581 ;
  assign n1607 = x0 & x39 ;
  assign n1608 = x1 & x38 ;
  assign n1609 = ( ~n1606 & n1607 ) | ( ~n1606 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1610 = ( n1606 & n1607 ) | ( n1606 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1611 = ( n1606 & n1609 ) | ( n1606 & ~n1610 ) | ( n1609 & ~n1610 ) ;
  assign n1612 = ( ~n1520 & n1584 ) | ( ~n1520 & n1611 ) | ( n1584 & n1611 ) ;
  assign n1613 = ( n1520 & n1584 ) | ( n1520 & n1611 ) | ( n1584 & n1611 ) ;
  assign n1614 = ( n1520 & n1612 ) | ( n1520 & ~n1613 ) | ( n1612 & ~n1613 ) ;
  assign n1615 = ( n1574 & ~n1605 ) | ( n1574 & n1614 ) | ( ~n1605 & n1614 ) ;
  assign n1616 = ( n1574 & n1605 ) | ( n1574 & n1614 ) | ( n1605 & n1614 ) ;
  assign n1617 = ( n1605 & n1615 ) | ( n1605 & ~n1616 ) | ( n1615 & ~n1616 ) ;
  assign n1618 = x17 & x22 ;
  assign n1619 = x4 & x35 ;
  assign n1620 = x12 & x27 ;
  assign n1621 = ( ~n1618 & n1619 ) | ( ~n1618 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1622 = ( n1618 & n1619 ) | ( n1618 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1623 = ( n1618 & n1621 ) | ( n1618 & ~n1622 ) | ( n1621 & ~n1622 ) ;
  assign n1624 = x19 & x20 ;
  assign n1625 = x18 & x21 ;
  assign n1626 = x8 & x31 ;
  assign n1627 = ( ~n1624 & n1625 ) | ( ~n1624 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1628 = ( n1624 & n1625 ) | ( n1624 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1629 = ( n1624 & n1627 ) | ( n1624 & ~n1628 ) | ( n1627 & ~n1628 ) ;
  assign n1630 = x10 & x29 ;
  assign n1631 = x5 & x34 ;
  assign n1632 = x11 & x28 ;
  assign n1633 = ( ~n1630 & n1631 ) | ( ~n1630 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1634 = ( n1630 & n1631 ) | ( n1630 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1635 = ( n1630 & n1633 ) | ( n1630 & ~n1634 ) | ( n1633 & ~n1634 ) ;
  assign n1636 = ( ~n1623 & n1629 ) | ( ~n1623 & n1635 ) | ( n1629 & n1635 ) ;
  assign n1637 = ( n1623 & n1629 ) | ( n1623 & n1635 ) | ( n1629 & n1635 ) ;
  assign n1638 = ( n1623 & n1636 ) | ( n1623 & ~n1637 ) | ( n1636 & ~n1637 ) ;
  assign n1639 = ( ~n1532 & n1538 ) | ( ~n1532 & n1554 ) | ( n1538 & n1554 ) ;
  assign n1640 = ( n1532 & n1538 ) | ( n1532 & n1554 ) | ( n1538 & n1554 ) ;
  assign n1641 = ( n1532 & n1639 ) | ( n1532 & ~n1640 ) | ( n1639 & ~n1640 ) ;
  assign n1642 = ( n1557 & n1638 ) | ( n1557 & n1641 ) | ( n1638 & n1641 ) ;
  assign n1643 = ( ~n1557 & n1638 ) | ( ~n1557 & n1641 ) | ( n1638 & n1641 ) ;
  assign n1644 = ( n1557 & ~n1642 ) | ( n1557 & n1643 ) | ( ~n1642 & n1643 ) ;
  assign n1645 = x13 & x26 ;
  assign n1646 = x3 & x36 ;
  assign n1647 = x2 & x37 ;
  assign n1648 = ( ~n1645 & n1646 ) | ( ~n1645 & n1647 ) | ( n1646 & n1647 ) ;
  assign n1649 = ( n1645 & n1646 ) | ( n1645 & n1647 ) | ( n1646 & n1647 ) ;
  assign n1650 = ( n1645 & n1648 ) | ( n1645 & ~n1649 ) | ( n1648 & ~n1649 ) ;
  assign n1651 = x15 & x24 ;
  assign n1652 = x16 & x23 ;
  assign n1653 = ( ~n785 & n1651 ) | ( ~n785 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1654 = ( n785 & n1651 ) | ( n785 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1655 = ( n785 & n1653 ) | ( n785 & ~n1654 ) | ( n1653 & ~n1654 ) ;
  assign n1656 = x7 & x32 ;
  assign n1657 = x9 & x30 ;
  assign n1658 = x6 & x33 ;
  assign n1659 = ( ~n1656 & n1657 ) | ( ~n1656 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = ( n1656 & n1657 ) | ( n1656 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1661 = ( n1656 & n1659 ) | ( n1656 & ~n1660 ) | ( n1659 & ~n1660 ) ;
  assign n1662 = ( ~n1650 & n1655 ) | ( ~n1650 & n1661 ) | ( n1655 & n1661 ) ;
  assign n1663 = ( n1650 & n1655 ) | ( n1650 & n1661 ) | ( n1655 & n1661 ) ;
  assign n1664 = ( n1650 & n1662 ) | ( n1650 & ~n1663 ) | ( n1662 & ~n1663 ) ;
  assign n1665 = ( n1543 & n1587 ) | ( n1543 & n1664 ) | ( n1587 & n1664 ) ;
  assign n1666 = ( ~n1543 & n1587 ) | ( ~n1543 & n1664 ) | ( n1587 & n1664 ) ;
  assign n1667 = ( n1543 & ~n1665 ) | ( n1543 & n1666 ) | ( ~n1665 & n1666 ) ;
  assign n1668 = ( n1547 & n1644 ) | ( n1547 & n1667 ) | ( n1644 & n1667 ) ;
  assign n1669 = ( ~n1547 & n1644 ) | ( ~n1547 & n1667 ) | ( n1644 & n1667 ) ;
  assign n1670 = ( n1547 & ~n1668 ) | ( n1547 & n1669 ) | ( ~n1668 & n1669 ) ;
  assign n1671 = ( n1589 & n1617 ) | ( n1589 & n1670 ) | ( n1617 & n1670 ) ;
  assign n1672 = ( ~n1589 & n1617 ) | ( ~n1589 & n1670 ) | ( n1617 & n1670 ) ;
  assign n1673 = ( n1589 & ~n1671 ) | ( n1589 & n1672 ) | ( ~n1671 & n1672 ) ;
  assign n1674 = ( n1593 & n1595 ) | ( n1593 & n1673 ) | ( n1595 & n1673 ) ;
  assign n1675 = ( n1593 & ~n1595 ) | ( n1593 & n1673 ) | ( ~n1595 & n1673 ) ;
  assign n1676 = ( n1595 & ~n1674 ) | ( n1595 & n1675 ) | ( ~n1674 & n1675 ) ;
  assign n1677 = x20 & x38 ;
  assign n1678 = ( ~x1 & x39 ) | ( ~x1 & n1677 ) | ( x39 & n1677 ) ;
  assign n1679 = ( x1 & x39 ) | ( x1 & n1677 ) | ( x39 & n1677 ) ;
  assign n1680 = ~n1678 & n1679 ;
  assign n1681 = x19 & x21 ;
  assign n1682 = ( n1628 & n1680 ) | ( n1628 & n1681 ) | ( n1680 & n1681 ) ;
  assign n1683 = ( ~n1628 & n1680 ) | ( ~n1628 & n1681 ) | ( n1680 & n1681 ) ;
  assign n1684 = ( n1628 & ~n1682 ) | ( n1628 & n1683 ) | ( ~n1682 & n1683 ) ;
  assign n1685 = ( n1600 & n1640 ) | ( n1600 & ~n1684 ) | ( n1640 & ~n1684 ) ;
  assign n1686 = ( n1600 & n1640 ) | ( n1600 & n1684 ) | ( n1640 & n1684 ) ;
  assign n1687 = ( n1684 & n1685 ) | ( n1684 & ~n1686 ) | ( n1685 & ~n1686 ) ;
  assign n1688 = x10 & x30 ;
  assign n1689 = x11 & x29 ;
  assign n1690 = x6 & x34 ;
  assign n1691 = ( ~n1688 & n1689 ) | ( ~n1688 & n1690 ) | ( n1689 & n1690 ) ;
  assign n1692 = ( n1688 & n1689 ) | ( n1688 & n1690 ) | ( n1689 & n1690 ) ;
  assign n1693 = ( n1688 & n1691 ) | ( n1688 & ~n1692 ) | ( n1691 & ~n1692 ) ;
  assign n1694 = x16 & x24 ;
  assign n1695 = x17 & x23 ;
  assign n1696 = x15 & x25 ;
  assign n1697 = ( ~n1694 & n1695 ) | ( ~n1694 & n1696 ) | ( n1695 & n1696 ) ;
  assign n1698 = ( n1694 & n1695 ) | ( n1694 & n1696 ) | ( n1695 & n1696 ) ;
  assign n1699 = ( n1694 & n1697 ) | ( n1694 & ~n1698 ) | ( n1697 & ~n1698 ) ;
  assign n1700 = x14 & x26 ;
  assign n1701 = x3 & x37 ;
  assign n1702 = x13 & x27 ;
  assign n1703 = ( ~n1700 & n1701 ) | ( ~n1700 & n1702 ) | ( n1701 & n1702 ) ;
  assign n1704 = ( n1700 & n1701 ) | ( n1700 & n1702 ) | ( n1701 & n1702 ) ;
  assign n1705 = ( n1700 & n1703 ) | ( n1700 & ~n1704 ) | ( n1703 & ~n1704 ) ;
  assign n1706 = ( ~n1693 & n1699 ) | ( ~n1693 & n1705 ) | ( n1699 & n1705 ) ;
  assign n1707 = ( n1693 & n1699 ) | ( n1693 & n1705 ) | ( n1699 & n1705 ) ;
  assign n1708 = ( n1693 & n1706 ) | ( n1693 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1709 = ( n1604 & n1687 ) | ( n1604 & n1708 ) | ( n1687 & n1708 ) ;
  assign n1710 = ( n1604 & ~n1687 ) | ( n1604 & n1708 ) | ( ~n1687 & n1708 ) ;
  assign n1711 = ( n1687 & ~n1709 ) | ( n1687 & n1710 ) | ( ~n1709 & n1710 ) ;
  assign n1712 = x38 & n534 ;
  assign n1713 = ( n1581 & n1610 ) | ( n1581 & ~n1712 ) | ( n1610 & ~n1712 ) ;
  assign n1714 = ( n1654 & n1660 ) | ( n1654 & ~n1713 ) | ( n1660 & ~n1713 ) ;
  assign n1715 = ( n1654 & n1660 ) | ( n1654 & n1713 ) | ( n1660 & n1713 ) ;
  assign n1716 = ( n1713 & n1714 ) | ( n1713 & ~n1715 ) | ( n1714 & ~n1715 ) ;
  assign n1717 = x7 & x33 ;
  assign n1718 = x8 & x32 ;
  assign n1719 = x9 & x31 ;
  assign n1720 = ( ~n1717 & n1718 ) | ( ~n1717 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1721 = ( n1717 & n1718 ) | ( n1717 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1722 = ( n1717 & n1720 ) | ( n1717 & ~n1721 ) | ( n1720 & ~n1721 ) ;
  assign n1723 = x18 & x22 ;
  assign n1724 = x0 & x40 ;
  assign n1725 = x2 & x38 ;
  assign n1726 = ( ~n1723 & n1724 ) | ( ~n1723 & n1725 ) | ( n1724 & n1725 ) ;
  assign n1727 = ( n1723 & n1724 ) | ( n1723 & n1725 ) | ( n1724 & n1725 ) ;
  assign n1728 = ( n1723 & n1726 ) | ( n1723 & ~n1727 ) | ( n1726 & ~n1727 ) ;
  assign n1729 = x12 & x28 ;
  assign n1730 = x4 & x36 ;
  assign n1731 = x5 & x35 ;
  assign n1732 = ( ~n1729 & n1730 ) | ( ~n1729 & n1731 ) | ( n1730 & n1731 ) ;
  assign n1733 = ( n1729 & n1730 ) | ( n1729 & n1731 ) | ( n1730 & n1731 ) ;
  assign n1734 = ( n1729 & n1732 ) | ( n1729 & ~n1733 ) | ( n1732 & ~n1733 ) ;
  assign n1735 = ( ~n1722 & n1728 ) | ( ~n1722 & n1734 ) | ( n1728 & n1734 ) ;
  assign n1736 = ( n1722 & n1728 ) | ( n1722 & n1734 ) | ( n1728 & n1734 ) ;
  assign n1737 = ( n1722 & n1735 ) | ( n1722 & ~n1736 ) | ( n1735 & ~n1736 ) ;
  assign n1738 = ( n1613 & n1716 ) | ( n1613 & n1737 ) | ( n1716 & n1737 ) ;
  assign n1739 = ( n1613 & ~n1716 ) | ( n1613 & n1737 ) | ( ~n1716 & n1737 ) ;
  assign n1740 = ( n1716 & ~n1738 ) | ( n1716 & n1739 ) | ( ~n1738 & n1739 ) ;
  assign n1741 = ( ~n1616 & n1711 ) | ( ~n1616 & n1740 ) | ( n1711 & n1740 ) ;
  assign n1742 = ( n1616 & n1711 ) | ( n1616 & n1740 ) | ( n1711 & n1740 ) ;
  assign n1743 = ( n1616 & n1741 ) | ( n1616 & ~n1742 ) | ( n1741 & ~n1742 ) ;
  assign n1744 = ( n1622 & n1634 ) | ( n1622 & ~n1649 ) | ( n1634 & ~n1649 ) ;
  assign n1745 = ( n1622 & n1634 ) | ( n1622 & n1649 ) | ( n1634 & n1649 ) ;
  assign n1746 = ( n1649 & n1744 ) | ( n1649 & ~n1745 ) | ( n1744 & ~n1745 ) ;
  assign n1747 = ( n1637 & n1663 ) | ( n1637 & n1746 ) | ( n1663 & n1746 ) ;
  assign n1748 = ( n1637 & n1663 ) | ( n1637 & ~n1746 ) | ( n1663 & ~n1746 ) ;
  assign n1749 = ( n1746 & ~n1747 ) | ( n1746 & n1748 ) | ( ~n1747 & n1748 ) ;
  assign n1750 = ( ~n1642 & n1665 ) | ( ~n1642 & n1749 ) | ( n1665 & n1749 ) ;
  assign n1751 = ( n1642 & n1665 ) | ( n1642 & n1749 ) | ( n1665 & n1749 ) ;
  assign n1752 = ( n1642 & n1750 ) | ( n1642 & ~n1751 ) | ( n1750 & ~n1751 ) ;
  assign n1753 = ( n1668 & n1743 ) | ( n1668 & n1752 ) | ( n1743 & n1752 ) ;
  assign n1754 = ( n1668 & ~n1743 ) | ( n1668 & n1752 ) | ( ~n1743 & n1752 ) ;
  assign n1755 = ( n1743 & ~n1753 ) | ( n1743 & n1754 ) | ( ~n1753 & n1754 ) ;
  assign n1756 = ( n1671 & ~n1674 ) | ( n1671 & n1755 ) | ( ~n1674 & n1755 ) ;
  assign n1757 = ( n1671 & n1674 ) | ( n1671 & n1755 ) | ( n1674 & n1755 ) ;
  assign n1758 = ( n1674 & n1756 ) | ( n1674 & ~n1757 ) | ( n1756 & ~n1757 ) ;
  assign n1759 = ( n1707 & ~n1715 ) | ( n1707 & n1745 ) | ( ~n1715 & n1745 ) ;
  assign n1760 = ( n1707 & n1715 ) | ( n1707 & n1745 ) | ( n1715 & n1745 ) ;
  assign n1761 = ( n1715 & n1759 ) | ( n1715 & ~n1760 ) | ( n1759 & ~n1760 ) ;
  assign n1762 = x0 & x41 ;
  assign n1763 = ( x2 & n66 ) | ( x2 & ~n1681 ) | ( n66 & ~n1681 ) ;
  assign n1764 = n67 & n1681 ;
  assign n1765 = ( x39 & n1763 ) | ( x39 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1766 = n1762 & n1765 ;
  assign n1767 = n1762 | n1765 ;
  assign n1768 = ~n1766 & n1767 ;
  assign n1769 = x13 & x28 ;
  assign n1770 = x3 & x38 ;
  assign n1771 = x15 & x26 ;
  assign n1772 = ( ~n1769 & n1770 ) | ( ~n1769 & n1771 ) | ( n1770 & n1771 ) ;
  assign n1773 = ( n1769 & n1770 ) | ( n1769 & n1771 ) | ( n1770 & n1771 ) ;
  assign n1774 = ( n1769 & n1772 ) | ( n1769 & ~n1773 ) | ( n1772 & ~n1773 ) ;
  assign n1775 = ( n1733 & n1768 ) | ( n1733 & n1774 ) | ( n1768 & n1774 ) ;
  assign n1776 = ( n1733 & ~n1768 ) | ( n1733 & n1774 ) | ( ~n1768 & n1774 ) ;
  assign n1777 = ( n1768 & ~n1775 ) | ( n1768 & n1776 ) | ( ~n1775 & n1776 ) ;
  assign n1778 = ( n1747 & n1761 ) | ( n1747 & n1777 ) | ( n1761 & n1777 ) ;
  assign n1779 = ( n1747 & ~n1761 ) | ( n1747 & n1777 ) | ( ~n1761 & n1777 ) ;
  assign n1780 = ( n1761 & ~n1778 ) | ( n1761 & n1779 ) | ( ~n1778 & n1779 ) ;
  assign n1781 = ( n1628 & ~n1684 ) | ( n1628 & n1712 ) | ( ~n1684 & n1712 ) ;
  assign n1782 = x19 & x22 ;
  assign n1783 = x20 & x21 ;
  assign n1784 = x8 & x33 ;
  assign n1785 = ( ~n1782 & n1783 ) | ( ~n1782 & n1784 ) | ( n1783 & n1784 ) ;
  assign n1786 = ( n1782 & n1783 ) | ( n1782 & n1784 ) | ( n1783 & n1784 ) ;
  assign n1787 = ( n1782 & n1785 ) | ( n1782 & ~n1786 ) | ( n1785 & ~n1786 ) ;
  assign n1788 = x6 & x35 ;
  assign n1789 = x5 & x36 ;
  assign n1790 = x11 & x30 ;
  assign n1791 = ( ~n1788 & n1789 ) | ( ~n1788 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1792 = ( n1788 & n1789 ) | ( n1788 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1793 = ( n1788 & n1791 ) | ( n1788 & ~n1792 ) | ( n1791 & ~n1792 ) ;
  assign n1794 = ( ~n1781 & n1787 ) | ( ~n1781 & n1793 ) | ( n1787 & n1793 ) ;
  assign n1795 = ( n1781 & n1787 ) | ( n1781 & n1793 ) | ( n1787 & n1793 ) ;
  assign n1796 = ( n1781 & n1794 ) | ( n1781 & ~n1795 ) | ( n1794 & ~n1795 ) ;
  assign n1797 = x16 & x25 ;
  assign n1798 = x18 & x23 ;
  assign n1799 = x17 & x24 ;
  assign n1800 = ( ~n1797 & n1798 ) | ( ~n1797 & n1799 ) | ( n1798 & n1799 ) ;
  assign n1801 = ( n1797 & n1798 ) | ( n1797 & n1799 ) | ( n1798 & n1799 ) ;
  assign n1802 = ( n1797 & n1800 ) | ( n1797 & ~n1801 ) | ( n1800 & ~n1801 ) ;
  assign n1803 = x14 & x27 ;
  assign n1804 = x12 & x29 ;
  assign n1805 = x4 & x37 ;
  assign n1806 = ( ~n1803 & n1804 ) | ( ~n1803 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1807 = ( n1803 & n1804 ) | ( n1803 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1808 = ( n1803 & n1806 ) | ( n1803 & ~n1807 ) | ( n1806 & ~n1807 ) ;
  assign n1809 = x10 & x31 ;
  assign n1810 = x9 & x32 ;
  assign n1811 = x7 & x34 ;
  assign n1812 = ( ~n1809 & n1810 ) | ( ~n1809 & n1811 ) | ( n1810 & n1811 ) ;
  assign n1813 = ( n1809 & n1810 ) | ( n1809 & n1811 ) | ( n1810 & n1811 ) ;
  assign n1814 = ( n1809 & n1812 ) | ( n1809 & ~n1813 ) | ( n1812 & ~n1813 ) ;
  assign n1815 = ( ~n1802 & n1808 ) | ( ~n1802 & n1814 ) | ( n1808 & n1814 ) ;
  assign n1816 = ( n1802 & n1808 ) | ( n1802 & n1814 ) | ( n1808 & n1814 ) ;
  assign n1817 = ( n1802 & n1815 ) | ( n1802 & ~n1816 ) | ( n1815 & ~n1816 ) ;
  assign n1818 = ( n1686 & n1796 ) | ( n1686 & n1817 ) | ( n1796 & n1817 ) ;
  assign n1819 = ( n1686 & ~n1796 ) | ( n1686 & n1817 ) | ( ~n1796 & n1817 ) ;
  assign n1820 = ( n1796 & ~n1818 ) | ( n1796 & n1819 ) | ( ~n1818 & n1819 ) ;
  assign n1821 = ( n1751 & ~n1780 ) | ( n1751 & n1820 ) | ( ~n1780 & n1820 ) ;
  assign n1822 = ( n1751 & n1780 ) | ( n1751 & n1820 ) | ( n1780 & n1820 ) ;
  assign n1823 = ( n1780 & n1821 ) | ( n1780 & ~n1822 ) | ( n1821 & ~n1822 ) ;
  assign n1824 = ~x1 & x21 ;
  assign n1825 = ( x1 & x21 ) | ( x1 & x40 ) | ( x21 & x40 ) ;
  assign n1826 = x21 & x40 ;
  assign n1827 = ( n1824 & n1825 ) | ( n1824 & ~n1826 ) | ( n1825 & ~n1826 ) ;
  assign n1828 = ( ~n1692 & n1721 ) | ( ~n1692 & n1827 ) | ( n1721 & n1827 ) ;
  assign n1829 = ( n1692 & n1721 ) | ( n1692 & n1827 ) | ( n1721 & n1827 ) ;
  assign n1830 = ( n1692 & n1828 ) | ( n1692 & ~n1829 ) | ( n1828 & ~n1829 ) ;
  assign n1831 = ( ~n1698 & n1704 ) | ( ~n1698 & n1727 ) | ( n1704 & n1727 ) ;
  assign n1832 = ( n1698 & n1704 ) | ( n1698 & n1727 ) | ( n1704 & n1727 ) ;
  assign n1833 = ( n1698 & n1831 ) | ( n1698 & ~n1832 ) | ( n1831 & ~n1832 ) ;
  assign n1834 = ( n1736 & n1830 ) | ( n1736 & n1833 ) | ( n1830 & n1833 ) ;
  assign n1835 = ( ~n1736 & n1830 ) | ( ~n1736 & n1833 ) | ( n1830 & n1833 ) ;
  assign n1836 = ( n1736 & ~n1834 ) | ( n1736 & n1835 ) | ( ~n1834 & n1835 ) ;
  assign n1837 = ( n1709 & n1738 ) | ( n1709 & n1836 ) | ( n1738 & n1836 ) ;
  assign n1838 = ( ~n1709 & n1738 ) | ( ~n1709 & n1836 ) | ( n1738 & n1836 ) ;
  assign n1839 = ( n1709 & ~n1837 ) | ( n1709 & n1838 ) | ( ~n1837 & n1838 ) ;
  assign n1840 = ( n1742 & n1823 ) | ( n1742 & n1839 ) | ( n1823 & n1839 ) ;
  assign n1841 = ( ~n1742 & n1823 ) | ( ~n1742 & n1839 ) | ( n1823 & n1839 ) ;
  assign n1842 = ( n1742 & ~n1840 ) | ( n1742 & n1841 ) | ( ~n1840 & n1841 ) ;
  assign n1843 = ( n1753 & n1757 ) | ( n1753 & n1842 ) | ( n1757 & n1842 ) ;
  assign n1844 = ( n1753 & ~n1757 ) | ( n1753 & n1842 ) | ( ~n1757 & n1842 ) ;
  assign n1845 = ( n1757 & ~n1843 ) | ( n1757 & n1844 ) | ( ~n1843 & n1844 ) ;
  assign n1846 = ( n1775 & n1816 ) | ( n1775 & ~n1832 ) | ( n1816 & ~n1832 ) ;
  assign n1847 = ( n1775 & n1816 ) | ( n1775 & n1832 ) | ( n1816 & n1832 ) ;
  assign n1848 = ( n1832 & n1846 ) | ( n1832 & ~n1847 ) | ( n1846 & ~n1847 ) ;
  assign n1849 = ( n1778 & n1818 ) | ( n1778 & n1848 ) | ( n1818 & n1848 ) ;
  assign n1850 = ( ~n1778 & n1818 ) | ( ~n1778 & n1848 ) | ( n1818 & n1848 ) ;
  assign n1851 = ( n1778 & ~n1849 ) | ( n1778 & n1850 ) | ( ~n1849 & n1850 ) ;
  assign n1852 = x17 & x25 ;
  assign n1853 = x19 & x23 ;
  assign n1854 = x18 & x24 ;
  assign n1855 = ( ~n1852 & n1853 ) | ( ~n1852 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1856 = ( n1852 & n1853 ) | ( n1852 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1857 = ( n1852 & n1855 ) | ( n1852 & ~n1856 ) | ( n1855 & ~n1856 ) ;
  assign n1858 = x14 & x28 ;
  assign n1859 = x4 & x38 ;
  assign n1860 = ( ~n895 & n1858 ) | ( ~n895 & n1859 ) | ( n1858 & n1859 ) ;
  assign n1861 = ( n895 & n1858 ) | ( n895 & n1859 ) | ( n1858 & n1859 ) ;
  assign n1862 = ( n895 & n1860 ) | ( n895 & ~n1861 ) | ( n1860 & ~n1861 ) ;
  assign n1863 = x3 & x39 ;
  assign n1864 = x16 & x26 ;
  assign n1865 = x2 & x40 ;
  assign n1866 = ( ~n1863 & n1864 ) | ( ~n1863 & n1865 ) | ( n1864 & n1865 ) ;
  assign n1867 = ( n1863 & n1864 ) | ( n1863 & n1865 ) | ( n1864 & n1865 ) ;
  assign n1868 = ( n1863 & n1866 ) | ( n1863 & ~n1867 ) | ( n1866 & ~n1867 ) ;
  assign n1869 = ( ~n1857 & n1862 ) | ( ~n1857 & n1868 ) | ( n1862 & n1868 ) ;
  assign n1870 = ( n1857 & n1862 ) | ( n1857 & n1868 ) | ( n1862 & n1868 ) ;
  assign n1871 = ( n1857 & n1869 ) | ( n1857 & ~n1870 ) | ( n1869 & ~n1870 ) ;
  assign n1872 = x6 & x36 ;
  assign n1873 = x11 & x31 ;
  assign n1874 = x7 & x35 ;
  assign n1875 = ( ~n1872 & n1873 ) | ( ~n1872 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1876 = ( n1872 & n1873 ) | ( n1872 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1877 = ( n1872 & n1875 ) | ( n1872 & ~n1876 ) | ( n1875 & ~n1876 ) ;
  assign n1878 = x9 & x33 ;
  assign n1879 = x8 & x34 ;
  assign n1880 = x10 & x32 ;
  assign n1881 = ( ~n1878 & n1879 ) | ( ~n1878 & n1880 ) | ( n1879 & n1880 ) ;
  assign n1882 = ( n1878 & n1879 ) | ( n1878 & n1880 ) | ( n1879 & n1880 ) ;
  assign n1883 = ( n1878 & n1881 ) | ( n1878 & ~n1882 ) | ( n1881 & ~n1882 ) ;
  assign n1884 = ( ~n1813 & n1877 ) | ( ~n1813 & n1883 ) | ( n1877 & n1883 ) ;
  assign n1885 = ( n1813 & n1877 ) | ( n1813 & n1883 ) | ( n1877 & n1883 ) ;
  assign n1886 = ( n1813 & n1884 ) | ( n1813 & ~n1885 ) | ( n1884 & ~n1885 ) ;
  assign n1887 = ( n1760 & n1871 ) | ( n1760 & n1886 ) | ( n1871 & n1886 ) ;
  assign n1888 = ( ~n1760 & n1871 ) | ( ~n1760 & n1886 ) | ( n1871 & n1886 ) ;
  assign n1889 = ( n1760 & ~n1887 ) | ( n1760 & n1888 ) | ( ~n1887 & n1888 ) ;
  assign n1890 = x20 & x22 ;
  assign n1891 = x1 & x41 ;
  assign n1892 = n1890 | n1891 ;
  assign n1893 = x22 & x41 ;
  assign n1894 = n534 & n1893 ;
  assign n1895 = n1892 & ~n1894 ;
  assign n1896 = x40 & n582 ;
  assign n1897 = x0 & x42 ;
  assign n1898 = ( n1895 & n1896 ) | ( n1895 & n1897 ) | ( n1896 & n1897 ) ;
  assign n1899 = ( ~n1895 & n1896 ) | ( ~n1895 & n1897 ) | ( n1896 & n1897 ) ;
  assign n1900 = ( n1895 & ~n1898 ) | ( n1895 & n1899 ) | ( ~n1898 & n1899 ) ;
  assign n1901 = x5 & x37 ;
  assign n1902 = x12 & x30 ;
  assign n1903 = x13 & x29 ;
  assign n1904 = ( ~n1901 & n1902 ) | ( ~n1901 & n1903 ) | ( n1902 & n1903 ) ;
  assign n1905 = ( n1901 & n1902 ) | ( n1901 & n1903 ) | ( n1902 & n1903 ) ;
  assign n1906 = ( n1901 & n1904 ) | ( n1901 & ~n1905 ) | ( n1904 & ~n1905 ) ;
  assign n1907 = ( n1829 & n1900 ) | ( n1829 & n1906 ) | ( n1900 & n1906 ) ;
  assign n1908 = ( n1829 & ~n1900 ) | ( n1829 & n1906 ) | ( ~n1900 & n1906 ) ;
  assign n1909 = ( n1900 & ~n1907 ) | ( n1900 & n1908 ) | ( ~n1907 & n1908 ) ;
  assign n1910 = x2 & n481 ;
  assign n1911 = x21 & x39 ;
  assign n1912 = n1910 & n1911 ;
  assign n1913 = n1766 | n1912 ;
  assign n1914 = ( n1773 & n1801 ) | ( n1773 & ~n1913 ) | ( n1801 & ~n1913 ) ;
  assign n1915 = ( n1773 & n1801 ) | ( n1773 & n1913 ) | ( n1801 & n1913 ) ;
  assign n1916 = ( n1913 & n1914 ) | ( n1913 & ~n1915 ) | ( n1914 & ~n1915 ) ;
  assign n1917 = ( n1786 & n1792 ) | ( n1786 & ~n1807 ) | ( n1792 & ~n1807 ) ;
  assign n1918 = ( n1786 & n1792 ) | ( n1786 & n1807 ) | ( n1792 & n1807 ) ;
  assign n1919 = ( n1807 & n1917 ) | ( n1807 & ~n1918 ) | ( n1917 & ~n1918 ) ;
  assign n1920 = ( n1795 & n1916 ) | ( n1795 & n1919 ) | ( n1916 & n1919 ) ;
  assign n1921 = ( ~n1795 & n1916 ) | ( ~n1795 & n1919 ) | ( n1916 & n1919 ) ;
  assign n1922 = ( n1795 & ~n1920 ) | ( n1795 & n1921 ) | ( ~n1920 & n1921 ) ;
  assign n1923 = ( n1834 & ~n1909 ) | ( n1834 & n1922 ) | ( ~n1909 & n1922 ) ;
  assign n1924 = ( n1834 & n1909 ) | ( n1834 & n1922 ) | ( n1909 & n1922 ) ;
  assign n1925 = ( n1909 & n1923 ) | ( n1909 & ~n1924 ) | ( n1923 & ~n1924 ) ;
  assign n1926 = ( n1837 & ~n1889 ) | ( n1837 & n1925 ) | ( ~n1889 & n1925 ) ;
  assign n1927 = ( n1837 & n1889 ) | ( n1837 & n1925 ) | ( n1889 & n1925 ) ;
  assign n1928 = ( n1889 & n1926 ) | ( n1889 & ~n1927 ) | ( n1926 & ~n1927 ) ;
  assign n1929 = ( n1822 & ~n1851 ) | ( n1822 & n1928 ) | ( ~n1851 & n1928 ) ;
  assign n1930 = ( n1822 & n1851 ) | ( n1822 & n1928 ) | ( n1851 & n1928 ) ;
  assign n1931 = ( n1851 & n1929 ) | ( n1851 & ~n1930 ) | ( n1929 & ~n1930 ) ;
  assign n1932 = ( n1840 & ~n1843 ) | ( n1840 & n1931 ) | ( ~n1843 & n1931 ) ;
  assign n1933 = ( n1840 & n1843 ) | ( n1840 & n1931 ) | ( n1843 & n1931 ) ;
  assign n1934 = ( n1843 & n1932 ) | ( n1843 & ~n1933 ) | ( n1932 & ~n1933 ) ;
  assign n1935 = x42 & n600 ;
  assign n1936 = x1 & x42 ;
  assign n1937 = x22 | n1936 ;
  assign n1938 = ~n1935 & n1937 ;
  assign n1939 = ( n1882 & n1894 ) | ( n1882 & n1938 ) | ( n1894 & n1938 ) ;
  assign n1940 = ( ~n1882 & n1894 ) | ( ~n1882 & n1938 ) | ( n1894 & n1938 ) ;
  assign n1941 = ( n1882 & ~n1939 ) | ( n1882 & n1940 ) | ( ~n1939 & n1940 ) ;
  assign n1942 = ( n1870 & n1885 ) | ( n1870 & ~n1941 ) | ( n1885 & ~n1941 ) ;
  assign n1943 = ( n1870 & n1885 ) | ( n1870 & n1941 ) | ( n1885 & n1941 ) ;
  assign n1944 = ( n1941 & n1942 ) | ( n1941 & ~n1943 ) | ( n1942 & ~n1943 ) ;
  assign n1945 = ( n1887 & n1924 ) | ( n1887 & n1944 ) | ( n1924 & n1944 ) ;
  assign n1946 = ( n1887 & n1924 ) | ( n1887 & ~n1944 ) | ( n1924 & ~n1944 ) ;
  assign n1947 = ( n1944 & ~n1945 ) | ( n1944 & n1946 ) | ( ~n1945 & n1946 ) ;
  assign n1948 = x19 & x24 ;
  assign n1949 = x17 & x26 ;
  assign n1950 = x18 & x25 ;
  assign n1951 = ( ~n1948 & n1949 ) | ( ~n1948 & n1950 ) | ( n1949 & n1950 ) ;
  assign n1952 = ( n1948 & n1949 ) | ( n1948 & n1950 ) | ( n1949 & n1950 ) ;
  assign n1953 = ( n1948 & n1951 ) | ( n1948 & ~n1952 ) | ( n1951 & ~n1952 ) ;
  assign n1954 = x4 & x39 ;
  assign n1955 = x0 & x43 ;
  assign n1956 = x3 & x40 ;
  assign n1957 = ( ~n1954 & n1955 ) | ( ~n1954 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1958 = ( n1954 & n1955 ) | ( n1954 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1959 = ( n1954 & n1957 ) | ( n1954 & ~n1958 ) | ( n1957 & ~n1958 ) ;
  assign n1960 = x16 & x27 ;
  assign n1961 = x15 & x28 ;
  assign n1962 = x14 & x29 ;
  assign n1963 = ( ~n1960 & n1961 ) | ( ~n1960 & n1962 ) | ( n1961 & n1962 ) ;
  assign n1964 = ( n1960 & n1961 ) | ( n1960 & n1962 ) | ( n1961 & n1962 ) ;
  assign n1965 = ( n1960 & n1963 ) | ( n1960 & ~n1964 ) | ( n1963 & ~n1964 ) ;
  assign n1966 = ( ~n1953 & n1959 ) | ( ~n1953 & n1965 ) | ( n1959 & n1965 ) ;
  assign n1967 = ( n1953 & n1959 ) | ( n1953 & n1965 ) | ( n1959 & n1965 ) ;
  assign n1968 = ( n1953 & n1966 ) | ( n1953 & ~n1967 ) | ( n1966 & ~n1967 ) ;
  assign n1969 = x21 & x22 ;
  assign n1970 = x9 & x34 ;
  assign n1971 = x20 & x23 ;
  assign n1972 = ( ~n1969 & n1970 ) | ( ~n1969 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1973 = ( n1969 & n1970 ) | ( n1969 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1974 = ( n1969 & n1972 ) | ( n1969 & ~n1973 ) | ( n1972 & ~n1973 ) ;
  assign n1975 = x8 & x35 ;
  assign n1976 = x7 & x36 ;
  assign n1977 = x10 & x33 ;
  assign n1978 = ( ~n1975 & n1976 ) | ( ~n1975 & n1977 ) | ( n1976 & n1977 ) ;
  assign n1979 = ( n1975 & n1976 ) | ( n1975 & n1977 ) | ( n1976 & n1977 ) ;
  assign n1980 = ( n1975 & n1978 ) | ( n1975 & ~n1979 ) | ( n1978 & ~n1979 ) ;
  assign n1981 = x13 & x30 ;
  assign n1982 = x5 & x38 ;
  assign n1983 = x2 & x41 ;
  assign n1984 = ( ~n1981 & n1982 ) | ( ~n1981 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1985 = ( n1981 & n1982 ) | ( n1981 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1986 = ( n1981 & n1984 ) | ( n1981 & ~n1985 ) | ( n1984 & ~n1985 ) ;
  assign n1987 = ( ~n1974 & n1980 ) | ( ~n1974 & n1986 ) | ( n1980 & n1986 ) ;
  assign n1988 = ( n1974 & n1980 ) | ( n1974 & n1986 ) | ( n1980 & n1986 ) ;
  assign n1989 = ( n1974 & n1987 ) | ( n1974 & ~n1988 ) | ( n1987 & ~n1988 ) ;
  assign n1990 = ( n1847 & n1968 ) | ( n1847 & n1989 ) | ( n1968 & n1989 ) ;
  assign n1991 = ( ~n1847 & n1968 ) | ( ~n1847 & n1989 ) | ( n1968 & n1989 ) ;
  assign n1992 = ( n1847 & ~n1990 ) | ( n1847 & n1991 ) | ( ~n1990 & n1991 ) ;
  assign n1993 = x6 & x37 ;
  assign n1994 = x11 & x32 ;
  assign n1995 = x12 & x31 ;
  assign n1996 = ( ~n1993 & n1994 ) | ( ~n1993 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1997 = ( n1993 & n1994 ) | ( n1993 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1998 = ( n1993 & n1996 ) | ( n1993 & ~n1997 ) | ( n1996 & ~n1997 ) ;
  assign n1999 = ( n1915 & n1918 ) | ( n1915 & ~n1998 ) | ( n1918 & ~n1998 ) ;
  assign n2000 = ( n1915 & n1918 ) | ( n1915 & n1998 ) | ( n1918 & n1998 ) ;
  assign n2001 = ( n1998 & n1999 ) | ( n1998 & ~n2000 ) | ( n1999 & ~n2000 ) ;
  assign n2002 = ( n1867 & ~n1898 ) | ( n1867 & n1905 ) | ( ~n1898 & n1905 ) ;
  assign n2003 = ( n1867 & n1898 ) | ( n1867 & n1905 ) | ( n1898 & n1905 ) ;
  assign n2004 = ( n1898 & n2002 ) | ( n1898 & ~n2003 ) | ( n2002 & ~n2003 ) ;
  assign n2005 = ( ~n1856 & n1861 ) | ( ~n1856 & n1876 ) | ( n1861 & n1876 ) ;
  assign n2006 = ( n1856 & n1861 ) | ( n1856 & n1876 ) | ( n1861 & n1876 ) ;
  assign n2007 = ( n1856 & n2005 ) | ( n1856 & ~n2006 ) | ( n2005 & ~n2006 ) ;
  assign n2008 = ( n1907 & n2004 ) | ( n1907 & n2007 ) | ( n2004 & n2007 ) ;
  assign n2009 = ( ~n1907 & n2004 ) | ( ~n1907 & n2007 ) | ( n2004 & n2007 ) ;
  assign n2010 = ( n1907 & ~n2008 ) | ( n1907 & n2009 ) | ( ~n2008 & n2009 ) ;
  assign n2011 = ( n1920 & n2001 ) | ( n1920 & n2010 ) | ( n2001 & n2010 ) ;
  assign n2012 = ( ~n1920 & n2001 ) | ( ~n1920 & n2010 ) | ( n2001 & n2010 ) ;
  assign n2013 = ( n1920 & ~n2011 ) | ( n1920 & n2012 ) | ( ~n2011 & n2012 ) ;
  assign n2014 = ( n1849 & n1992 ) | ( n1849 & n2013 ) | ( n1992 & n2013 ) ;
  assign n2015 = ( n1849 & ~n1992 ) | ( n1849 & n2013 ) | ( ~n1992 & n2013 ) ;
  assign n2016 = ( n1992 & ~n2014 ) | ( n1992 & n2015 ) | ( ~n2014 & n2015 ) ;
  assign n2017 = ( n1927 & ~n1947 ) | ( n1927 & n2016 ) | ( ~n1947 & n2016 ) ;
  assign n2018 = ( n1927 & n1947 ) | ( n1927 & n2016 ) | ( n1947 & n2016 ) ;
  assign n2019 = ( n1947 & n2017 ) | ( n1947 & ~n2018 ) | ( n2017 & ~n2018 ) ;
  assign n2020 = ( n1930 & ~n1933 ) | ( n1930 & n2019 ) | ( ~n1933 & n2019 ) ;
  assign n2021 = ( n1930 & n1933 ) | ( n1930 & n2019 ) | ( n1933 & n2019 ) ;
  assign n2022 = ( n1933 & n2020 ) | ( n1933 & ~n2021 ) | ( n2020 & ~n2021 ) ;
  assign n2023 = x8 & x36 ;
  assign n2024 = x9 & x35 ;
  assign n2025 = x10 & x34 ;
  assign n2026 = ( ~n2023 & n2024 ) | ( ~n2023 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2027 = ( n2023 & n2024 ) | ( n2023 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2028 = ( n2023 & n2026 ) | ( n2023 & ~n2027 ) | ( n2026 & ~n2027 ) ;
  assign n2029 = x16 & x28 ;
  assign n2030 = x4 & x40 ;
  assign n2031 = x14 & x30 ;
  assign n2032 = ( ~n2029 & n2030 ) | ( ~n2029 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = ( n2029 & n2030 ) | ( n2029 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2034 = ( n2029 & n2032 ) | ( n2029 & ~n2033 ) | ( n2032 & ~n2033 ) ;
  assign n2035 = x12 & x32 ;
  assign n2036 = x5 & x39 ;
  assign n2037 = x13 & x31 ;
  assign n2038 = ( ~n2035 & n2036 ) | ( ~n2035 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2039 = ( n2035 & n2036 ) | ( n2035 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2040 = ( n2035 & n2038 ) | ( n2035 & ~n2039 ) | ( n2038 & ~n2039 ) ;
  assign n2041 = ( ~n2028 & n2034 ) | ( ~n2028 & n2040 ) | ( n2034 & n2040 ) ;
  assign n2042 = ( n2028 & n2034 ) | ( n2028 & n2040 ) | ( n2034 & n2040 ) ;
  assign n2043 = ( n2028 & n2041 ) | ( n2028 & ~n2042 ) | ( n2041 & ~n2042 ) ;
  assign n2044 = x7 & x37 ;
  assign n2045 = x11 & x33 ;
  assign n2046 = x6 & x38 ;
  assign n2047 = ( ~n2044 & n2045 ) | ( ~n2044 & n2046 ) | ( n2045 & n2046 ) ;
  assign n2048 = ( n2044 & n2045 ) | ( n2044 & n2046 ) | ( n2045 & n2046 ) ;
  assign n2049 = ( n2044 & n2047 ) | ( n2044 & ~n2048 ) | ( n2047 & ~n2048 ) ;
  assign n2050 = x20 & x24 ;
  assign n2051 = x19 & x25 ;
  assign n2052 = x18 & x26 ;
  assign n2053 = ( ~n2050 & n2051 ) | ( ~n2050 & n2052 ) | ( n2051 & n2052 ) ;
  assign n2054 = ( n2050 & n2051 ) | ( n2050 & n2052 ) | ( n2051 & n2052 ) ;
  assign n2055 = ( n2050 & n2053 ) | ( n2050 & ~n2054 ) | ( n2053 & ~n2054 ) ;
  assign n2056 = x17 & x27 ;
  assign n2057 = x15 & x29 ;
  assign n2058 = x3 & x41 ;
  assign n2059 = ( ~n2056 & n2057 ) | ( ~n2056 & n2058 ) | ( n2057 & n2058 ) ;
  assign n2060 = ( n2056 & n2057 ) | ( n2056 & n2058 ) | ( n2057 & n2058 ) ;
  assign n2061 = ( n2056 & n2059 ) | ( n2056 & ~n2060 ) | ( n2059 & ~n2060 ) ;
  assign n2062 = ( ~n2049 & n2055 ) | ( ~n2049 & n2061 ) | ( n2055 & n2061 ) ;
  assign n2063 = ( n2049 & n2055 ) | ( n2049 & n2061 ) | ( n2055 & n2061 ) ;
  assign n2064 = ( n2049 & n2062 ) | ( n2049 & ~n2063 ) | ( n2062 & ~n2063 ) ;
  assign n2065 = ( n1943 & n2043 ) | ( n1943 & n2064 ) | ( n2043 & n2064 ) ;
  assign n2066 = ( ~n1943 & n2043 ) | ( ~n1943 & n2064 ) | ( n2043 & n2064 ) ;
  assign n2067 = ( n1943 & ~n2065 ) | ( n1943 & n2066 ) | ( ~n2065 & n2066 ) ;
  assign n2068 = ( n1939 & ~n2003 ) | ( n1939 & n2006 ) | ( ~n2003 & n2006 ) ;
  assign n2069 = ( n1939 & n2003 ) | ( n1939 & n2006 ) | ( n2003 & n2006 ) ;
  assign n2070 = ( n2003 & n2068 ) | ( n2003 & ~n2069 ) | ( n2068 & ~n2069 ) ;
  assign n2071 = x21 & x23 ;
  assign n2072 = x1 & x43 ;
  assign n2073 = n2071 | n2072 ;
  assign n2074 = x23 & x43 ;
  assign n2075 = n582 & n2074 ;
  assign n2076 = n2073 & ~n2075 ;
  assign n2077 = ( ~n1973 & n1979 ) | ( ~n1973 & n2076 ) | ( n1979 & n2076 ) ;
  assign n2078 = ( n1973 & n1979 ) | ( n1973 & n2076 ) | ( n1979 & n2076 ) ;
  assign n2079 = ( n1973 & n2077 ) | ( n1973 & ~n2078 ) | ( n2077 & ~n2078 ) ;
  assign n2080 = x2 & x42 ;
  assign n2081 = x0 & x44 ;
  assign n2082 = ( ~n1935 & n2080 ) | ( ~n1935 & n2081 ) | ( n2080 & n2081 ) ;
  assign n2083 = ( n1935 & n2080 ) | ( n1935 & n2081 ) | ( n2080 & n2081 ) ;
  assign n2084 = ( n1935 & n2082 ) | ( n1935 & ~n2083 ) | ( n2082 & ~n2083 ) ;
  assign n2085 = ( n1964 & n1997 ) | ( n1964 & ~n2084 ) | ( n1997 & ~n2084 ) ;
  assign n2086 = ( n1964 & n1997 ) | ( n1964 & n2084 ) | ( n1997 & n2084 ) ;
  assign n2087 = ( n2084 & n2085 ) | ( n2084 & ~n2086 ) | ( n2085 & ~n2086 ) ;
  assign n2088 = ( n2000 & ~n2079 ) | ( n2000 & n2087 ) | ( ~n2079 & n2087 ) ;
  assign n2089 = ( n2000 & n2079 ) | ( n2000 & n2087 ) | ( n2079 & n2087 ) ;
  assign n2090 = ( n2079 & n2088 ) | ( n2079 & ~n2089 ) | ( n2088 & ~n2089 ) ;
  assign n2091 = ( n2008 & ~n2070 ) | ( n2008 & n2090 ) | ( ~n2070 & n2090 ) ;
  assign n2092 = ( n2008 & n2070 ) | ( n2008 & n2090 ) | ( n2070 & n2090 ) ;
  assign n2093 = ( n2070 & n2091 ) | ( n2070 & ~n2092 ) | ( n2091 & ~n2092 ) ;
  assign n2094 = ( n1945 & n2067 ) | ( n1945 & n2093 ) | ( n2067 & n2093 ) ;
  assign n2095 = ( ~n1945 & n2067 ) | ( ~n1945 & n2093 ) | ( n2067 & n2093 ) ;
  assign n2096 = ( n1945 & ~n2094 ) | ( n1945 & n2095 ) | ( ~n2094 & n2095 ) ;
  assign n2097 = ( ~n1952 & n1958 ) | ( ~n1952 & n1985 ) | ( n1958 & n1985 ) ;
  assign n2098 = ( n1952 & n1958 ) | ( n1952 & n1985 ) | ( n1958 & n1985 ) ;
  assign n2099 = ( n1952 & n2097 ) | ( n1952 & ~n2098 ) | ( n2097 & ~n2098 ) ;
  assign n2100 = ( n1967 & n1988 ) | ( n1967 & n2099 ) | ( n1988 & n2099 ) ;
  assign n2101 = ( ~n1967 & n1988 ) | ( ~n1967 & n2099 ) | ( n1988 & n2099 ) ;
  assign n2102 = ( n1967 & ~n2100 ) | ( n1967 & n2101 ) | ( ~n2100 & n2101 ) ;
  assign n2103 = ( n1990 & n2011 ) | ( n1990 & n2102 ) | ( n2011 & n2102 ) ;
  assign n2104 = ( n1990 & ~n2011 ) | ( n1990 & n2102 ) | ( ~n2011 & n2102 ) ;
  assign n2105 = ( n2011 & ~n2103 ) | ( n2011 & n2104 ) | ( ~n2103 & n2104 ) ;
  assign n2106 = ( ~n2014 & n2096 ) | ( ~n2014 & n2105 ) | ( n2096 & n2105 ) ;
  assign n2107 = ( n2014 & n2096 ) | ( n2014 & n2105 ) | ( n2096 & n2105 ) ;
  assign n2108 = ( n2014 & n2106 ) | ( n2014 & ~n2107 ) | ( n2106 & ~n2107 ) ;
  assign n2109 = ( n2018 & ~n2021 ) | ( n2018 & n2108 ) | ( ~n2021 & n2108 ) ;
  assign n2110 = ( n2018 & n2021 ) | ( n2018 & n2108 ) | ( n2021 & n2108 ) ;
  assign n2111 = ( n2021 & n2109 ) | ( n2021 & ~n2110 ) | ( n2109 & ~n2110 ) ;
  assign n2112 = x1 & x44 ;
  assign n2113 = x23 & ~n2075 ;
  assign n2114 = x3 & x42 ;
  assign n2115 = ( ~n2112 & n2113 ) | ( ~n2112 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2116 = ( n2112 & n2113 ) | ( n2112 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2117 = ( n2112 & n2115 ) | ( n2112 & ~n2116 ) | ( n2115 & ~n2116 ) ;
  assign n2118 = x12 & x33 ;
  assign n2119 = x11 & x34 ;
  assign n2120 = x6 & x39 ;
  assign n2121 = ( ~n2118 & n2119 ) | ( ~n2118 & n2120 ) | ( n2119 & n2120 ) ;
  assign n2122 = ( n2118 & n2119 ) | ( n2118 & n2120 ) | ( n2119 & n2120 ) ;
  assign n2123 = ( n2118 & n2121 ) | ( n2118 & ~n2122 ) | ( n2121 & ~n2122 ) ;
  assign n2124 = x15 & x30 ;
  assign n2125 = x17 & x28 ;
  assign n2126 = ( ~n973 & n2124 ) | ( ~n973 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( n973 & n2124 ) | ( n973 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2128 = ( n973 & n2126 ) | ( n973 & ~n2127 ) | ( n2126 & ~n2127 ) ;
  assign n2129 = ( n2117 & n2123 ) | ( n2117 & n2128 ) | ( n2123 & n2128 ) ;
  assign n2130 = ( ~n2117 & n2123 ) | ( ~n2117 & n2128 ) | ( n2123 & n2128 ) ;
  assign n2131 = ( n2117 & ~n2129 ) | ( n2117 & n2130 ) | ( ~n2129 & n2130 ) ;
  assign n2132 = ( n2054 & n2060 ) | ( n2054 & ~n2083 ) | ( n2060 & ~n2083 ) ;
  assign n2133 = ( n2054 & n2060 ) | ( n2054 & n2083 ) | ( n2060 & n2083 ) ;
  assign n2134 = ( n2083 & n2132 ) | ( n2083 & ~n2133 ) | ( n2132 & ~n2133 ) ;
  assign n2135 = ( n2069 & n2131 ) | ( n2069 & n2134 ) | ( n2131 & n2134 ) ;
  assign n2136 = ( ~n2069 & n2131 ) | ( ~n2069 & n2134 ) | ( n2131 & n2134 ) ;
  assign n2137 = ( n2069 & ~n2135 ) | ( n2069 & n2136 ) | ( ~n2135 & n2136 ) ;
  assign n2138 = ( n2065 & n2092 ) | ( n2065 & n2137 ) | ( n2092 & n2137 ) ;
  assign n2139 = ( n2065 & n2092 ) | ( n2065 & ~n2137 ) | ( n2092 & ~n2137 ) ;
  assign n2140 = ( n2137 & ~n2138 ) | ( n2137 & n2139 ) | ( ~n2138 & n2139 ) ;
  assign n2141 = x5 & x40 ;
  assign n2142 = x14 & x31 ;
  assign n2143 = x13 & x32 ;
  assign n2144 = ( ~n2141 & n2142 ) | ( ~n2141 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2145 = ( n2141 & n2142 ) | ( n2141 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2146 = ( n2141 & n2144 ) | ( n2141 & ~n2145 ) | ( n2144 & ~n2145 ) ;
  assign n2147 = x18 & x27 ;
  assign n2148 = x20 & x25 ;
  assign n2149 = x19 & x26 ;
  assign n2150 = ( ~n2147 & n2148 ) | ( ~n2147 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = ( n2147 & n2148 ) | ( n2147 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2152 = ( n2147 & n2150 ) | ( n2147 & ~n2151 ) | ( n2150 & ~n2151 ) ;
  assign n2153 = ( ~n2027 & n2146 ) | ( ~n2027 & n2152 ) | ( n2146 & n2152 ) ;
  assign n2154 = ( n2027 & n2146 ) | ( n2027 & n2152 ) | ( n2146 & n2152 ) ;
  assign n2155 = ( n2027 & n2153 ) | ( n2027 & ~n2154 ) | ( n2153 & ~n2154 ) ;
  assign n2156 = x22 & x23 ;
  assign n2157 = x10 & x35 ;
  assign n2158 = x21 & x24 ;
  assign n2159 = ( ~n2156 & n2157 ) | ( ~n2156 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = ( n2156 & n2157 ) | ( n2156 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2161 = ( n2156 & n2159 ) | ( n2156 & ~n2160 ) | ( n2159 & ~n2160 ) ;
  assign n2162 = x8 & x37 ;
  assign n2163 = x7 & x38 ;
  assign n2164 = x9 & x36 ;
  assign n2165 = ( ~n2162 & n2163 ) | ( ~n2162 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2166 = ( n2162 & n2163 ) | ( n2162 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2167 = ( n2162 & n2165 ) | ( n2162 & ~n2166 ) | ( n2165 & ~n2166 ) ;
  assign n2168 = x4 & x41 ;
  assign n2169 = x0 & x45 ;
  assign n2170 = x2 & x43 ;
  assign n2171 = ( ~n2168 & n2169 ) | ( ~n2168 & n2170 ) | ( n2169 & n2170 ) ;
  assign n2172 = ( n2168 & n2169 ) | ( n2168 & n2170 ) | ( n2169 & n2170 ) ;
  assign n2173 = ( n2168 & n2171 ) | ( n2168 & ~n2172 ) | ( n2171 & ~n2172 ) ;
  assign n2174 = ( ~n2161 & n2167 ) | ( ~n2161 & n2173 ) | ( n2167 & n2173 ) ;
  assign n2175 = ( n2161 & n2167 ) | ( n2161 & n2173 ) | ( n2167 & n2173 ) ;
  assign n2176 = ( n2161 & n2174 ) | ( n2161 & ~n2175 ) | ( n2174 & ~n2175 ) ;
  assign n2177 = ( n2100 & n2155 ) | ( n2100 & n2176 ) | ( n2155 & n2176 ) ;
  assign n2178 = ( ~n2100 & n2155 ) | ( ~n2100 & n2176 ) | ( n2155 & n2176 ) ;
  assign n2179 = ( n2100 & ~n2177 ) | ( n2100 & n2178 ) | ( ~n2177 & n2178 ) ;
  assign n2180 = ( n2033 & ~n2039 ) | ( n2033 & n2048 ) | ( ~n2039 & n2048 ) ;
  assign n2181 = ( n2033 & n2039 ) | ( n2033 & n2048 ) | ( n2039 & n2048 ) ;
  assign n2182 = ( n2039 & n2180 ) | ( n2039 & ~n2181 ) | ( n2180 & ~n2181 ) ;
  assign n2183 = ( n2042 & n2063 ) | ( n2042 & n2182 ) | ( n2063 & n2182 ) ;
  assign n2184 = ( ~n2042 & n2063 ) | ( ~n2042 & n2182 ) | ( n2063 & n2182 ) ;
  assign n2185 = ( n2042 & ~n2183 ) | ( n2042 & n2184 ) | ( ~n2183 & n2184 ) ;
  assign n2186 = ( ~n2078 & n2086 ) | ( ~n2078 & n2098 ) | ( n2086 & n2098 ) ;
  assign n2187 = ( n2078 & n2086 ) | ( n2078 & n2098 ) | ( n2086 & n2098 ) ;
  assign n2188 = ( n2078 & n2186 ) | ( n2078 & ~n2187 ) | ( n2186 & ~n2187 ) ;
  assign n2189 = ( n2089 & ~n2185 ) | ( n2089 & n2188 ) | ( ~n2185 & n2188 ) ;
  assign n2190 = ( n2089 & n2185 ) | ( n2089 & n2188 ) | ( n2185 & n2188 ) ;
  assign n2191 = ( n2185 & n2189 ) | ( n2185 & ~n2190 ) | ( n2189 & ~n2190 ) ;
  assign n2192 = ( n2103 & n2179 ) | ( n2103 & n2191 ) | ( n2179 & n2191 ) ;
  assign n2193 = ( ~n2103 & n2179 ) | ( ~n2103 & n2191 ) | ( n2179 & n2191 ) ;
  assign n2194 = ( n2103 & ~n2192 ) | ( n2103 & n2193 ) | ( ~n2192 & n2193 ) ;
  assign n2195 = ( n2094 & n2140 ) | ( n2094 & n2194 ) | ( n2140 & n2194 ) ;
  assign n2196 = ( ~n2094 & n2140 ) | ( ~n2094 & n2194 ) | ( n2140 & n2194 ) ;
  assign n2197 = ( n2094 & ~n2195 ) | ( n2094 & n2196 ) | ( ~n2195 & n2196 ) ;
  assign n2198 = ( n2107 & n2110 ) | ( n2107 & n2197 ) | ( n2110 & n2197 ) ;
  assign n2199 = ( n2107 & ~n2110 ) | ( n2107 & n2197 ) | ( ~n2110 & n2197 ) ;
  assign n2200 = ( n2110 & ~n2198 ) | ( n2110 & n2199 ) | ( ~n2198 & n2199 ) ;
  assign n2201 = ( ~n2129 & n2154 ) | ( ~n2129 & n2175 ) | ( n2154 & n2175 ) ;
  assign n2202 = ( n2129 & n2154 ) | ( n2129 & n2175 ) | ( n2154 & n2175 ) ;
  assign n2203 = ( n2129 & n2201 ) | ( n2129 & ~n2202 ) | ( n2201 & ~n2202 ) ;
  assign n2204 = ( ~n2145 & n2166 ) | ( ~n2145 & n2172 ) | ( n2166 & n2172 ) ;
  assign n2205 = ( n2145 & n2166 ) | ( n2145 & n2172 ) | ( n2166 & n2172 ) ;
  assign n2206 = ( n2145 & n2204 ) | ( n2145 & ~n2205 ) | ( n2204 & ~n2205 ) ;
  assign n2207 = x22 & x24 ;
  assign n2208 = x1 & x45 ;
  assign n2209 = n2207 & n2208 ;
  assign n2210 = n2207 | n2208 ;
  assign n2211 = ~n2209 & n2210 ;
  assign n2212 = x23 & n2112 ;
  assign n2213 = ( n2160 & ~n2211 ) | ( n2160 & n2212 ) | ( ~n2211 & n2212 ) ;
  assign n2214 = ( n2160 & n2211 ) | ( n2160 & n2212 ) | ( n2211 & n2212 ) ;
  assign n2215 = ( n2211 & n2213 ) | ( n2211 & ~n2214 ) | ( n2213 & ~n2214 ) ;
  assign n2216 = ( n2133 & n2206 ) | ( n2133 & n2215 ) | ( n2206 & n2215 ) ;
  assign n2217 = ( ~n2133 & n2206 ) | ( ~n2133 & n2215 ) | ( n2206 & n2215 ) ;
  assign n2218 = ( n2133 & ~n2216 ) | ( n2133 & n2217 ) | ( ~n2216 & n2217 ) ;
  assign n2219 = ( n2135 & n2203 ) | ( n2135 & n2218 ) | ( n2203 & n2218 ) ;
  assign n2220 = ( ~n2135 & n2203 ) | ( ~n2135 & n2218 ) | ( n2203 & n2218 ) ;
  assign n2221 = ( n2135 & ~n2219 ) | ( n2135 & n2220 ) | ( ~n2219 & n2220 ) ;
  assign n2222 = ( n2075 & n2116 ) | ( n2075 & ~n2212 ) | ( n2116 & ~n2212 ) ;
  assign n2223 = x12 & x34 ;
  assign n2224 = x7 & x39 ;
  assign n2225 = x8 & x38 ;
  assign n2226 = ( ~n2223 & n2224 ) | ( ~n2223 & n2225 ) | ( n2224 & n2225 ) ;
  assign n2227 = ( n2223 & n2224 ) | ( n2223 & n2225 ) | ( n2224 & n2225 ) ;
  assign n2228 = ( n2223 & n2226 ) | ( n2223 & ~n2227 ) | ( n2226 & ~n2227 ) ;
  assign n2229 = x16 & x30 ;
  assign n2230 = x18 & x28 ;
  assign n2231 = x17 & x29 ;
  assign n2232 = ( ~n2229 & n2230 ) | ( ~n2229 & n2231 ) | ( n2230 & n2231 ) ;
  assign n2233 = ( n2229 & n2230 ) | ( n2229 & n2231 ) | ( n2230 & n2231 ) ;
  assign n2234 = ( n2229 & n2232 ) | ( n2229 & ~n2233 ) | ( n2232 & ~n2233 ) ;
  assign n2235 = ( ~n2222 & n2228 ) | ( ~n2222 & n2234 ) | ( n2228 & n2234 ) ;
  assign n2236 = ( n2222 & n2228 ) | ( n2222 & n2234 ) | ( n2228 & n2234 ) ;
  assign n2237 = ( n2222 & n2235 ) | ( n2222 & ~n2236 ) | ( n2235 & ~n2236 ) ;
  assign n2238 = x19 & x27 ;
  assign n2239 = x21 & x25 ;
  assign n2240 = x20 & x26 ;
  assign n2241 = ( ~n2238 & n2239 ) | ( ~n2238 & n2240 ) | ( n2239 & n2240 ) ;
  assign n2242 = ( n2238 & n2239 ) | ( n2238 & n2240 ) | ( n2239 & n2240 ) ;
  assign n2243 = ( n2238 & n2241 ) | ( n2238 & ~n2242 ) | ( n2241 & ~n2242 ) ;
  assign n2244 = x10 & x36 ;
  assign n2245 = x11 & x35 ;
  assign n2246 = x9 & x37 ;
  assign n2247 = ( ~n2244 & n2245 ) | ( ~n2244 & n2246 ) | ( n2245 & n2246 ) ;
  assign n2248 = ( n2244 & n2245 ) | ( n2244 & n2246 ) | ( n2245 & n2246 ) ;
  assign n2249 = ( n2244 & n2247 ) | ( n2244 & ~n2248 ) | ( n2247 & ~n2248 ) ;
  assign n2250 = x4 & x42 ;
  assign n2251 = x3 & x43 ;
  assign n2252 = x0 & x46 ;
  assign n2253 = ( ~n2250 & n2251 ) | ( ~n2250 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2254 = ( n2250 & n2251 ) | ( n2250 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2255 = ( n2250 & n2253 ) | ( n2250 & ~n2254 ) | ( n2253 & ~n2254 ) ;
  assign n2256 = ( ~n2243 & n2249 ) | ( ~n2243 & n2255 ) | ( n2249 & n2255 ) ;
  assign n2257 = ( n2243 & n2249 ) | ( n2243 & n2255 ) | ( n2249 & n2255 ) ;
  assign n2258 = ( n2243 & n2256 ) | ( n2243 & ~n2257 ) | ( n2256 & ~n2257 ) ;
  assign n2259 = ( n2183 & n2237 ) | ( n2183 & n2258 ) | ( n2237 & n2258 ) ;
  assign n2260 = ( n2183 & ~n2237 ) | ( n2183 & n2258 ) | ( ~n2237 & n2258 ) ;
  assign n2261 = ( n2237 & ~n2259 ) | ( n2237 & n2260 ) | ( ~n2259 & n2260 ) ;
  assign n2262 = ( ~n2138 & n2221 ) | ( ~n2138 & n2261 ) | ( n2221 & n2261 ) ;
  assign n2263 = ( n2138 & n2221 ) | ( n2138 & n2261 ) | ( n2221 & n2261 ) ;
  assign n2264 = ( n2138 & n2262 ) | ( n2138 & ~n2263 ) | ( n2262 & ~n2263 ) ;
  assign n2265 = x2 & x44 ;
  assign n2266 = x5 & x41 ;
  assign n2267 = ( ~n1204 & n2265 ) | ( ~n1204 & n2266 ) | ( n2265 & n2266 ) ;
  assign n2268 = ( n1204 & n2265 ) | ( n1204 & n2266 ) | ( n2265 & n2266 ) ;
  assign n2269 = ( n1204 & n2267 ) | ( n1204 & ~n2268 ) | ( n2267 & ~n2268 ) ;
  assign n2270 = x13 & x33 ;
  assign n2271 = x14 & x32 ;
  assign n2272 = x6 & x40 ;
  assign n2273 = ( ~n2270 & n2271 ) | ( ~n2270 & n2272 ) | ( n2271 & n2272 ) ;
  assign n2274 = ( n2270 & n2271 ) | ( n2270 & n2272 ) | ( n2271 & n2272 ) ;
  assign n2275 = ( n2270 & n2273 ) | ( n2270 & ~n2274 ) | ( n2273 & ~n2274 ) ;
  assign n2276 = ( ~n2181 & n2269 ) | ( ~n2181 & n2275 ) | ( n2269 & n2275 ) ;
  assign n2277 = ( n2181 & n2269 ) | ( n2181 & n2275 ) | ( n2269 & n2275 ) ;
  assign n2278 = ( n2181 & n2276 ) | ( n2181 & ~n2277 ) | ( n2276 & ~n2277 ) ;
  assign n2279 = ( n2122 & n2127 ) | ( n2122 & ~n2151 ) | ( n2127 & ~n2151 ) ;
  assign n2280 = ( n2122 & n2127 ) | ( n2122 & n2151 ) | ( n2127 & n2151 ) ;
  assign n2281 = ( n2151 & n2279 ) | ( n2151 & ~n2280 ) | ( n2279 & ~n2280 ) ;
  assign n2282 = ( n2187 & ~n2278 ) | ( n2187 & n2281 ) | ( ~n2278 & n2281 ) ;
  assign n2283 = ( n2187 & n2278 ) | ( n2187 & n2281 ) | ( n2278 & n2281 ) ;
  assign n2284 = ( n2278 & n2282 ) | ( n2278 & ~n2283 ) | ( n2282 & ~n2283 ) ;
  assign n2285 = ( n2177 & n2190 ) | ( n2177 & ~n2284 ) | ( n2190 & ~n2284 ) ;
  assign n2286 = ( n2177 & n2190 ) | ( n2177 & n2284 ) | ( n2190 & n2284 ) ;
  assign n2287 = ( n2284 & n2285 ) | ( n2284 & ~n2286 ) | ( n2285 & ~n2286 ) ;
  assign n2288 = ( n2192 & n2195 ) | ( n2192 & n2287 ) | ( n2195 & n2287 ) ;
  assign n2289 = ( n2192 & ~n2195 ) | ( n2192 & n2287 ) | ( ~n2195 & n2287 ) ;
  assign n2290 = ( n2195 & ~n2288 ) | ( n2195 & n2289 ) | ( ~n2288 & n2289 ) ;
  assign n2291 = ( n2198 & n2264 ) | ( n2198 & n2290 ) | ( n2264 & n2290 ) ;
  assign n2292 = ( ~n2198 & n2264 ) | ( ~n2198 & n2290 ) | ( n2264 & n2290 ) ;
  assign n2293 = ( n2198 & ~n2291 ) | ( n2198 & n2292 ) | ( ~n2291 & n2292 ) ;
  assign n2294 = x13 & x34 ;
  assign n2295 = x7 & x40 ;
  assign n2296 = x12 & x35 ;
  assign n2297 = ( ~n2294 & n2295 ) | ( ~n2294 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = ( n2294 & n2295 ) | ( n2294 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2299 = ( n2294 & n2297 ) | ( n2294 & ~n2298 ) | ( n2297 & ~n2298 ) ;
  assign n2300 = ( n2214 & ~n2280 ) | ( n2214 & n2299 ) | ( ~n2280 & n2299 ) ;
  assign n2301 = ( n2214 & n2280 ) | ( n2214 & n2299 ) | ( n2280 & n2299 ) ;
  assign n2302 = ( n2280 & n2300 ) | ( n2280 & ~n2301 ) | ( n2300 & ~n2301 ) ;
  assign n2303 = ( n2202 & n2216 ) | ( n2202 & n2302 ) | ( n2216 & n2302 ) ;
  assign n2304 = ( ~n2202 & n2216 ) | ( ~n2202 & n2302 ) | ( n2216 & n2302 ) ;
  assign n2305 = ( n2202 & ~n2303 ) | ( n2202 & n2304 ) | ( ~n2303 & n2304 ) ;
  assign n2306 = ~x1 & x24 ;
  assign n2307 = ( x1 & x24 ) | ( x1 & x46 ) | ( x24 & x46 ) ;
  assign n2308 = x24 & x46 ;
  assign n2309 = ( n2306 & n2307 ) | ( n2306 & ~n2308 ) | ( n2307 & ~n2308 ) ;
  assign n2310 = ( n2227 & ~n2248 ) | ( n2227 & n2309 ) | ( ~n2248 & n2309 ) ;
  assign n2311 = ( n2227 & n2248 ) | ( n2227 & n2309 ) | ( n2248 & n2309 ) ;
  assign n2312 = ( n2248 & n2310 ) | ( n2248 & ~n2311 ) | ( n2310 & ~n2311 ) ;
  assign n2313 = ( n2205 & n2236 ) | ( n2205 & ~n2312 ) | ( n2236 & ~n2312 ) ;
  assign n2314 = ( n2205 & n2236 ) | ( n2205 & n2312 ) | ( n2236 & n2312 ) ;
  assign n2315 = ( n2312 & n2313 ) | ( n2312 & ~n2314 ) | ( n2313 & ~n2314 ) ;
  assign n2316 = x2 & x45 ;
  assign n2317 = x0 & x47 ;
  assign n2318 = ( ~n2209 & n2316 ) | ( ~n2209 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2319 = ( n2209 & n2316 ) | ( n2209 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2320 = ( n2209 & n2318 ) | ( n2209 & ~n2319 ) | ( n2318 & ~n2319 ) ;
  assign n2321 = x17 & x30 ;
  assign n2322 = x16 & x31 ;
  assign n2323 = x18 & x29 ;
  assign n2324 = ( ~n2321 & n2322 ) | ( ~n2321 & n2323 ) | ( n2322 & n2323 ) ;
  assign n2325 = ( n2321 & n2322 ) | ( n2321 & n2323 ) | ( n2322 & n2323 ) ;
  assign n2326 = ( n2321 & n2324 ) | ( n2321 & ~n2325 ) | ( n2324 & ~n2325 ) ;
  assign n2327 = x19 & x28 ;
  assign n2328 = x20 & x27 ;
  assign n2329 = x21 & x26 ;
  assign n2330 = ( ~n2327 & n2328 ) | ( ~n2327 & n2329 ) | ( n2328 & n2329 ) ;
  assign n2331 = ( n2327 & n2328 ) | ( n2327 & n2329 ) | ( n2328 & n2329 ) ;
  assign n2332 = ( n2327 & n2330 ) | ( n2327 & ~n2331 ) | ( n2330 & ~n2331 ) ;
  assign n2333 = ( ~n2320 & n2326 ) | ( ~n2320 & n2332 ) | ( n2326 & n2332 ) ;
  assign n2334 = ( n2320 & n2326 ) | ( n2320 & n2332 ) | ( n2326 & n2332 ) ;
  assign n2335 = ( n2320 & n2333 ) | ( n2320 & ~n2334 ) | ( n2333 & ~n2334 ) ;
  assign n2336 = x15 & x32 ;
  assign n2337 = x4 & x43 ;
  assign n2338 = x3 & x44 ;
  assign n2339 = ( ~n2336 & n2337 ) | ( ~n2336 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2340 = ( n2336 & n2337 ) | ( n2336 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2341 = ( n2336 & n2339 ) | ( n2336 & ~n2340 ) | ( n2339 & ~n2340 ) ;
  assign n2342 = ( n2233 & n2274 ) | ( n2233 & ~n2341 ) | ( n2274 & ~n2341 ) ;
  assign n2343 = ( n2233 & n2274 ) | ( n2233 & n2341 ) | ( n2274 & n2341 ) ;
  assign n2344 = ( n2341 & n2342 ) | ( n2341 & ~n2343 ) | ( n2342 & ~n2343 ) ;
  assign n2345 = x8 & x39 ;
  assign n2346 = x11 & x36 ;
  assign n2347 = x9 & x38 ;
  assign n2348 = ( ~n2345 & n2346 ) | ( ~n2345 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2349 = ( n2345 & n2346 ) | ( n2345 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2350 = ( n2345 & n2348 ) | ( n2345 & ~n2349 ) | ( n2348 & ~n2349 ) ;
  assign n2351 = x23 & x24 ;
  assign n2352 = x10 & x37 ;
  assign n2353 = x22 & x25 ;
  assign n2354 = ( ~n2351 & n2352 ) | ( ~n2351 & n2353 ) | ( n2352 & n2353 ) ;
  assign n2355 = ( n2351 & n2352 ) | ( n2351 & n2353 ) | ( n2352 & n2353 ) ;
  assign n2356 = ( n2351 & n2354 ) | ( n2351 & ~n2355 ) | ( n2354 & ~n2355 ) ;
  assign n2357 = x5 & x42 ;
  assign n2358 = x6 & x41 ;
  assign n2359 = x14 & x33 ;
  assign n2360 = ( ~n2357 & n2358 ) | ( ~n2357 & n2359 ) | ( n2358 & n2359 ) ;
  assign n2361 = ( n2357 & n2358 ) | ( n2357 & n2359 ) | ( n2358 & n2359 ) ;
  assign n2362 = ( n2357 & n2360 ) | ( n2357 & ~n2361 ) | ( n2360 & ~n2361 ) ;
  assign n2363 = ( ~n2350 & n2356 ) | ( ~n2350 & n2362 ) | ( n2356 & n2362 ) ;
  assign n2364 = ( n2350 & n2356 ) | ( n2350 & n2362 ) | ( n2356 & n2362 ) ;
  assign n2365 = ( n2350 & n2363 ) | ( n2350 & ~n2364 ) | ( n2363 & ~n2364 ) ;
  assign n2366 = ( ~n2335 & n2344 ) | ( ~n2335 & n2365 ) | ( n2344 & n2365 ) ;
  assign n2367 = ( n2335 & n2344 ) | ( n2335 & n2365 ) | ( n2344 & n2365 ) ;
  assign n2368 = ( n2335 & n2366 ) | ( n2335 & ~n2367 ) | ( n2366 & ~n2367 ) ;
  assign n2369 = ( n2305 & n2315 ) | ( n2305 & n2368 ) | ( n2315 & n2368 ) ;
  assign n2370 = ( ~n2305 & n2315 ) | ( ~n2305 & n2368 ) | ( n2315 & n2368 ) ;
  assign n2371 = ( n2305 & ~n2369 ) | ( n2305 & n2370 ) | ( ~n2369 & n2370 ) ;
  assign n2372 = ( n2242 & n2254 ) | ( n2242 & ~n2268 ) | ( n2254 & ~n2268 ) ;
  assign n2373 = ( n2242 & n2254 ) | ( n2242 & n2268 ) | ( n2254 & n2268 ) ;
  assign n2374 = ( n2268 & n2372 ) | ( n2268 & ~n2373 ) | ( n2372 & ~n2373 ) ;
  assign n2375 = ( n2257 & n2277 ) | ( n2257 & n2374 ) | ( n2277 & n2374 ) ;
  assign n2376 = ( n2257 & ~n2277 ) | ( n2257 & n2374 ) | ( ~n2277 & n2374 ) ;
  assign n2377 = ( n2277 & ~n2375 ) | ( n2277 & n2376 ) | ( ~n2375 & n2376 ) ;
  assign n2378 = ( n2259 & n2283 ) | ( n2259 & n2377 ) | ( n2283 & n2377 ) ;
  assign n2379 = ( n2259 & ~n2283 ) | ( n2259 & n2377 ) | ( ~n2283 & n2377 ) ;
  assign n2380 = ( n2283 & ~n2378 ) | ( n2283 & n2379 ) | ( ~n2378 & n2379 ) ;
  assign n2381 = ( n2219 & n2286 ) | ( n2219 & n2380 ) | ( n2286 & n2380 ) ;
  assign n2382 = ( n2219 & ~n2286 ) | ( n2219 & n2380 ) | ( ~n2286 & n2380 ) ;
  assign n2383 = ( n2286 & ~n2381 ) | ( n2286 & n2382 ) | ( ~n2381 & n2382 ) ;
  assign n2384 = ( n2263 & n2371 ) | ( n2263 & n2383 ) | ( n2371 & n2383 ) ;
  assign n2385 = ( ~n2263 & n2371 ) | ( ~n2263 & n2383 ) | ( n2371 & n2383 ) ;
  assign n2386 = ( n2263 & ~n2384 ) | ( n2263 & n2385 ) | ( ~n2384 & n2385 ) ;
  assign n2387 = ( n2288 & n2291 ) | ( n2288 & n2386 ) | ( n2291 & n2386 ) ;
  assign n2388 = ( n2288 & ~n2291 ) | ( n2288 & n2386 ) | ( ~n2291 & n2386 ) ;
  assign n2389 = ( n2291 & ~n2387 ) | ( n2291 & n2388 ) | ( ~n2387 & n2388 ) ;
  assign n2390 = x23 & x25 ;
  assign n2391 = x1 & x47 ;
  assign n2392 = n2390 | n2391 ;
  assign n2393 = x25 & x47 ;
  assign n2394 = n648 & n2393 ;
  assign n2395 = n2392 & ~n2394 ;
  assign n2396 = x46 & n695 ;
  assign n2397 = x0 & x48 ;
  assign n2398 = ( n2395 & n2396 ) | ( n2395 & n2397 ) | ( n2396 & n2397 ) ;
  assign n2399 = ( ~n2395 & n2396 ) | ( ~n2395 & n2397 ) | ( n2396 & n2397 ) ;
  assign n2400 = ( n2395 & ~n2398 ) | ( n2395 & n2399 ) | ( ~n2398 & n2399 ) ;
  assign n2401 = ( n2343 & n2373 ) | ( n2343 & n2400 ) | ( n2373 & n2400 ) ;
  assign n2402 = ( n2343 & n2373 ) | ( n2343 & ~n2400 ) | ( n2373 & ~n2400 ) ;
  assign n2403 = ( n2400 & ~n2401 ) | ( n2400 & n2402 ) | ( ~n2401 & n2402 ) ;
  assign n2404 = ( ~n2314 & n2375 ) | ( ~n2314 & n2403 ) | ( n2375 & n2403 ) ;
  assign n2405 = ( n2314 & n2375 ) | ( n2314 & n2403 ) | ( n2375 & n2403 ) ;
  assign n2406 = ( n2314 & n2404 ) | ( n2314 & ~n2405 ) | ( n2404 & ~n2405 ) ;
  assign n2407 = ( ~n2319 & n2325 ) | ( ~n2319 & n2340 ) | ( n2325 & n2340 ) ;
  assign n2408 = ( n2319 & n2325 ) | ( n2319 & n2340 ) | ( n2325 & n2340 ) ;
  assign n2409 = ( n2319 & n2407 ) | ( n2319 & ~n2408 ) | ( n2407 & ~n2408 ) ;
  assign n2410 = ( n2311 & n2334 ) | ( n2311 & n2409 ) | ( n2334 & n2409 ) ;
  assign n2411 = ( n2311 & n2334 ) | ( n2311 & ~n2409 ) | ( n2334 & ~n2409 ) ;
  assign n2412 = ( n2409 & ~n2410 ) | ( n2409 & n2411 ) | ( ~n2410 & n2411 ) ;
  assign n2413 = x3 & x45 ;
  assign n2414 = x2 & x46 ;
  assign n2415 = x16 & x32 ;
  assign n2416 = ( ~n2413 & n2414 ) | ( ~n2413 & n2415 ) | ( n2414 & n2415 ) ;
  assign n2417 = ( n2413 & n2414 ) | ( n2413 & n2415 ) | ( n2414 & n2415 ) ;
  assign n2418 = ( n2413 & n2416 ) | ( n2413 & ~n2417 ) | ( n2416 & ~n2417 ) ;
  assign n2419 = ( n2298 & n2355 ) | ( n2298 & ~n2418 ) | ( n2355 & ~n2418 ) ;
  assign n2420 = ( n2298 & n2355 ) | ( n2298 & n2418 ) | ( n2355 & n2418 ) ;
  assign n2421 = ( n2418 & n2419 ) | ( n2418 & ~n2420 ) | ( n2419 & ~n2420 ) ;
  assign n2422 = ( n2331 & ~n2349 ) | ( n2331 & n2361 ) | ( ~n2349 & n2361 ) ;
  assign n2423 = ( n2331 & n2349 ) | ( n2331 & n2361 ) | ( n2349 & n2361 ) ;
  assign n2424 = ( n2349 & n2422 ) | ( n2349 & ~n2423 ) | ( n2422 & ~n2423 ) ;
  assign n2425 = ( n2364 & n2421 ) | ( n2364 & n2424 ) | ( n2421 & n2424 ) ;
  assign n2426 = ( n2364 & ~n2421 ) | ( n2364 & n2424 ) | ( ~n2421 & n2424 ) ;
  assign n2427 = ( n2421 & ~n2425 ) | ( n2421 & n2426 ) | ( ~n2425 & n2426 ) ;
  assign n2428 = ( ~n2367 & n2412 ) | ( ~n2367 & n2427 ) | ( n2412 & n2427 ) ;
  assign n2429 = ( n2367 & n2412 ) | ( n2367 & n2427 ) | ( n2412 & n2427 ) ;
  assign n2430 = ( n2367 & n2428 ) | ( n2367 & ~n2429 ) | ( n2428 & ~n2429 ) ;
  assign n2431 = ( n2369 & n2406 ) | ( n2369 & n2430 ) | ( n2406 & n2430 ) ;
  assign n2432 = ( ~n2369 & n2406 ) | ( ~n2369 & n2430 ) | ( n2406 & n2430 ) ;
  assign n2433 = ( n2369 & ~n2431 ) | ( n2369 & n2432 ) | ( ~n2431 & n2432 ) ;
  assign n2434 = x12 & x36 ;
  assign n2435 = x8 & x40 ;
  assign n2436 = x7 & x41 ;
  assign n2437 = ( ~n2434 & n2435 ) | ( ~n2434 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2438 = ( n2434 & n2435 ) | ( n2434 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2439 = ( n2434 & n2437 ) | ( n2434 & ~n2438 ) | ( n2437 & ~n2438 ) ;
  assign n2440 = x9 & x39 ;
  assign n2441 = x10 & x38 ;
  assign n2442 = x11 & x37 ;
  assign n2443 = ( ~n2440 & n2441 ) | ( ~n2440 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2444 = ( n2440 & n2441 ) | ( n2440 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2445 = ( n2440 & n2443 ) | ( n2440 & ~n2444 ) | ( n2443 & ~n2444 ) ;
  assign n2446 = x14 & x34 ;
  assign n2447 = x13 & x35 ;
  assign n2448 = x6 & x42 ;
  assign n2449 = ( ~n2446 & n2447 ) | ( ~n2446 & n2448 ) | ( n2447 & n2448 ) ;
  assign n2450 = ( n2446 & n2447 ) | ( n2446 & n2448 ) | ( n2447 & n2448 ) ;
  assign n2451 = ( n2446 & n2449 ) | ( n2446 & ~n2450 ) | ( n2449 & ~n2450 ) ;
  assign n2452 = ( ~n2439 & n2445 ) | ( ~n2439 & n2451 ) | ( n2445 & n2451 ) ;
  assign n2453 = ( n2439 & n2445 ) | ( n2439 & n2451 ) | ( n2445 & n2451 ) ;
  assign n2454 = ( n2439 & n2452 ) | ( n2439 & ~n2453 ) | ( n2452 & ~n2453 ) ;
  assign n2455 = x4 & x44 ;
  assign n2456 = x15 & x33 ;
  assign n2457 = x5 & x43 ;
  assign n2458 = ( ~n2455 & n2456 ) | ( ~n2455 & n2457 ) | ( n2456 & n2457 ) ;
  assign n2459 = ( n2455 & n2456 ) | ( n2455 & n2457 ) | ( n2456 & n2457 ) ;
  assign n2460 = ( n2455 & n2458 ) | ( n2455 & ~n2459 ) | ( n2458 & ~n2459 ) ;
  assign n2461 = x17 & x31 ;
  assign n2462 = x19 & x29 ;
  assign n2463 = x18 & x30 ;
  assign n2464 = ( ~n2461 & n2462 ) | ( ~n2461 & n2463 ) | ( n2462 & n2463 ) ;
  assign n2465 = ( n2461 & n2462 ) | ( n2461 & n2463 ) | ( n2462 & n2463 ) ;
  assign n2466 = ( n2461 & n2464 ) | ( n2461 & ~n2465 ) | ( n2464 & ~n2465 ) ;
  assign n2467 = x22 & x26 ;
  assign n2468 = x20 & x28 ;
  assign n2469 = x21 & x27 ;
  assign n2470 = ( ~n2467 & n2468 ) | ( ~n2467 & n2469 ) | ( n2468 & n2469 ) ;
  assign n2471 = ( n2467 & n2468 ) | ( n2467 & n2469 ) | ( n2468 & n2469 ) ;
  assign n2472 = ( n2467 & n2470 ) | ( n2467 & ~n2471 ) | ( n2470 & ~n2471 ) ;
  assign n2473 = ( ~n2460 & n2466 ) | ( ~n2460 & n2472 ) | ( n2466 & n2472 ) ;
  assign n2474 = ( n2460 & n2466 ) | ( n2460 & n2472 ) | ( n2466 & n2472 ) ;
  assign n2475 = ( n2460 & n2473 ) | ( n2460 & ~n2474 ) | ( n2473 & ~n2474 ) ;
  assign n2476 = ( n2301 & n2454 ) | ( n2301 & n2475 ) | ( n2454 & n2475 ) ;
  assign n2477 = ( ~n2301 & n2454 ) | ( ~n2301 & n2475 ) | ( n2454 & n2475 ) ;
  assign n2478 = ( n2301 & ~n2476 ) | ( n2301 & n2477 ) | ( ~n2476 & n2477 ) ;
  assign n2479 = ( n2303 & n2378 ) | ( n2303 & n2478 ) | ( n2378 & n2478 ) ;
  assign n2480 = ( n2303 & ~n2378 ) | ( n2303 & n2478 ) | ( ~n2378 & n2478 ) ;
  assign n2481 = ( n2378 & ~n2479 ) | ( n2378 & n2480 ) | ( ~n2479 & n2480 ) ;
  assign n2482 = ( n2381 & n2433 ) | ( n2381 & n2481 ) | ( n2433 & n2481 ) ;
  assign n2483 = ( ~n2381 & n2433 ) | ( ~n2381 & n2481 ) | ( n2433 & n2481 ) ;
  assign n2484 = ( n2381 & ~n2482 ) | ( n2381 & n2483 ) | ( ~n2482 & n2483 ) ;
  assign n2485 = ( n2384 & n2387 ) | ( n2384 & n2484 ) | ( n2387 & n2484 ) ;
  assign n2486 = ( n2384 & ~n2387 ) | ( n2384 & n2484 ) | ( ~n2387 & n2484 ) ;
  assign n2487 = ( n2387 & ~n2485 ) | ( n2387 & n2486 ) | ( ~n2485 & n2486 ) ;
  assign n2488 = ( n2408 & n2420 ) | ( n2408 & n2423 ) | ( n2420 & n2423 ) ;
  assign n2489 = ( ~n2408 & n2420 ) | ( ~n2408 & n2423 ) | ( n2420 & n2423 ) ;
  assign n2490 = ( n2408 & ~n2488 ) | ( n2408 & n2489 ) | ( ~n2488 & n2489 ) ;
  assign n2491 = ( n2410 & n2425 ) | ( n2410 & n2490 ) | ( n2425 & n2490 ) ;
  assign n2492 = ( n2410 & ~n2425 ) | ( n2410 & n2490 ) | ( ~n2425 & n2490 ) ;
  assign n2493 = ( n2425 & ~n2491 ) | ( n2425 & n2492 ) | ( ~n2491 & n2492 ) ;
  assign n2494 = ( n2438 & ~n2450 ) | ( n2438 & n2465 ) | ( ~n2450 & n2465 ) ;
  assign n2495 = ( n2438 & n2450 ) | ( n2438 & n2465 ) | ( n2450 & n2465 ) ;
  assign n2496 = ( n2450 & n2494 ) | ( n2450 & ~n2495 ) | ( n2494 & ~n2495 ) ;
  assign n2497 = ( n2401 & n2474 ) | ( n2401 & ~n2496 ) | ( n2474 & ~n2496 ) ;
  assign n2498 = ( n2401 & n2474 ) | ( n2401 & n2496 ) | ( n2474 & n2496 ) ;
  assign n2499 = ( n2496 & n2497 ) | ( n2496 & ~n2498 ) | ( n2497 & ~n2498 ) ;
  assign n2500 = ( x25 & ~n2391 ) | ( x25 & n2395 ) | ( ~n2391 & n2395 ) ;
  assign n2501 = x1 & x48 ;
  assign n2502 = ( n2444 & n2500 ) | ( n2444 & ~n2501 ) | ( n2500 & ~n2501 ) ;
  assign n2503 = ( ~n2444 & n2500 ) | ( ~n2444 & n2501 ) | ( n2500 & n2501 ) ;
  assign n2504 = ( ~n2500 & n2502 ) | ( ~n2500 & n2503 ) | ( n2502 & n2503 ) ;
  assign n2505 = ( n2417 & ~n2459 ) | ( n2417 & n2471 ) | ( ~n2459 & n2471 ) ;
  assign n2506 = ( n2417 & n2459 ) | ( n2417 & n2471 ) | ( n2459 & n2471 ) ;
  assign n2507 = ( n2459 & n2505 ) | ( n2459 & ~n2506 ) | ( n2505 & ~n2506 ) ;
  assign n2508 = ( n2453 & n2504 ) | ( n2453 & n2507 ) | ( n2504 & n2507 ) ;
  assign n2509 = ( n2453 & ~n2504 ) | ( n2453 & n2507 ) | ( ~n2504 & n2507 ) ;
  assign n2510 = ( n2504 & ~n2508 ) | ( n2504 & n2509 ) | ( ~n2508 & n2509 ) ;
  assign n2511 = ( n2476 & n2499 ) | ( n2476 & n2510 ) | ( n2499 & n2510 ) ;
  assign n2512 = ( n2476 & ~n2499 ) | ( n2476 & n2510 ) | ( ~n2499 & n2510 ) ;
  assign n2513 = ( n2499 & ~n2511 ) | ( n2499 & n2512 ) | ( ~n2511 & n2512 ) ;
  assign n2514 = ( n2479 & n2493 ) | ( n2479 & n2513 ) | ( n2493 & n2513 ) ;
  assign n2515 = ( ~n2479 & n2493 ) | ( ~n2479 & n2513 ) | ( n2493 & n2513 ) ;
  assign n2516 = ( n2479 & ~n2514 ) | ( n2479 & n2515 ) | ( ~n2514 & n2515 ) ;
  assign n2517 = x16 & x33 ;
  assign n2518 = x18 & x31 ;
  assign n2519 = x17 & x32 ;
  assign n2520 = ( ~n2517 & n2518 ) | ( ~n2517 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2521 = ( n2517 & n2518 ) | ( n2517 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2522 = ( n2517 & n2520 ) | ( n2517 & ~n2521 ) | ( n2520 & ~n2521 ) ;
  assign n2523 = x5 & x44 ;
  assign n2524 = x4 & x45 ;
  assign n2525 = x0 & x49 ;
  assign n2526 = ( ~n2523 & n2524 ) | ( ~n2523 & n2525 ) | ( n2524 & n2525 ) ;
  assign n2527 = ( n2523 & n2524 ) | ( n2523 & n2525 ) | ( n2524 & n2525 ) ;
  assign n2528 = ( n2523 & n2526 ) | ( n2523 & ~n2527 ) | ( n2526 & ~n2527 ) ;
  assign n2529 = ( ~n2398 & n2522 ) | ( ~n2398 & n2528 ) | ( n2522 & n2528 ) ;
  assign n2530 = ( n2398 & n2522 ) | ( n2398 & n2528 ) | ( n2522 & n2528 ) ;
  assign n2531 = ( n2398 & n2529 ) | ( n2398 & ~n2530 ) | ( n2529 & ~n2530 ) ;
  assign n2532 = x8 & x41 ;
  assign n2533 = x7 & x42 ;
  assign n2534 = x13 & x36 ;
  assign n2535 = ( ~n2532 & n2533 ) | ( ~n2532 & n2534 ) | ( n2533 & n2534 ) ;
  assign n2536 = ( n2532 & n2533 ) | ( n2532 & n2534 ) | ( n2533 & n2534 ) ;
  assign n2537 = ( n2532 & n2535 ) | ( n2532 & ~n2536 ) | ( n2535 & ~n2536 ) ;
  assign n2538 = x15 & x34 ;
  assign n2539 = x6 & x43 ;
  assign n2540 = x14 & x35 ;
  assign n2541 = ( ~n2538 & n2539 ) | ( ~n2538 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = ( n2538 & n2539 ) | ( n2538 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2543 = ( n2538 & n2541 ) | ( n2538 & ~n2542 ) | ( n2541 & ~n2542 ) ;
  assign n2544 = x24 & x25 ;
  assign n2545 = x23 & x26 ;
  assign n2546 = x11 & x38 ;
  assign n2547 = ( ~n2544 & n2545 ) | ( ~n2544 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2548 = ( n2544 & n2545 ) | ( n2544 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2549 = ( n2544 & n2547 ) | ( n2544 & ~n2548 ) | ( n2547 & ~n2548 ) ;
  assign n2550 = ( ~n2537 & n2543 ) | ( ~n2537 & n2549 ) | ( n2543 & n2549 ) ;
  assign n2551 = ( n2537 & n2543 ) | ( n2537 & n2549 ) | ( n2543 & n2549 ) ;
  assign n2552 = ( n2537 & n2550 ) | ( n2537 & ~n2551 ) | ( n2550 & ~n2551 ) ;
  assign n2553 = x12 & x37 ;
  assign n2554 = x9 & x40 ;
  assign n2555 = x10 & x39 ;
  assign n2556 = ( ~n2553 & n2554 ) | ( ~n2553 & n2555 ) | ( n2554 & n2555 ) ;
  assign n2557 = ( n2553 & n2554 ) | ( n2553 & n2555 ) | ( n2554 & n2555 ) ;
  assign n2558 = ( n2553 & n2556 ) | ( n2553 & ~n2557 ) | ( n2556 & ~n2557 ) ;
  assign n2559 = x21 & x28 ;
  assign n2560 = x19 & x30 ;
  assign n2561 = x20 & x29 ;
  assign n2562 = ( ~n2559 & n2560 ) | ( ~n2559 & n2561 ) | ( n2560 & n2561 ) ;
  assign n2563 = ( n2559 & n2560 ) | ( n2559 & n2561 ) | ( n2560 & n2561 ) ;
  assign n2564 = ( n2559 & n2562 ) | ( n2559 & ~n2563 ) | ( n2562 & ~n2563 ) ;
  assign n2565 = x2 & x47 ;
  assign n2566 = x22 & x27 ;
  assign n2567 = x3 & x46 ;
  assign n2568 = ( ~n2565 & n2566 ) | ( ~n2565 & n2567 ) | ( n2566 & n2567 ) ;
  assign n2569 = ( n2565 & n2566 ) | ( n2565 & n2567 ) | ( n2566 & n2567 ) ;
  assign n2570 = ( n2565 & n2568 ) | ( n2565 & ~n2569 ) | ( n2568 & ~n2569 ) ;
  assign n2571 = ( ~n2558 & n2564 ) | ( ~n2558 & n2570 ) | ( n2564 & n2570 ) ;
  assign n2572 = ( n2558 & n2564 ) | ( n2558 & n2570 ) | ( n2564 & n2570 ) ;
  assign n2573 = ( n2558 & n2571 ) | ( n2558 & ~n2572 ) | ( n2571 & ~n2572 ) ;
  assign n2574 = ( ~n2531 & n2552 ) | ( ~n2531 & n2573 ) | ( n2552 & n2573 ) ;
  assign n2575 = ( n2531 & n2552 ) | ( n2531 & n2573 ) | ( n2552 & n2573 ) ;
  assign n2576 = ( n2531 & n2574 ) | ( n2531 & ~n2575 ) | ( n2574 & ~n2575 ) ;
  assign n2577 = ( ~n2405 & n2429 ) | ( ~n2405 & n2576 ) | ( n2429 & n2576 ) ;
  assign n2578 = ( n2405 & n2429 ) | ( n2405 & n2576 ) | ( n2429 & n2576 ) ;
  assign n2579 = ( n2405 & n2577 ) | ( n2405 & ~n2578 ) | ( n2577 & ~n2578 ) ;
  assign n2580 = ( n2431 & n2516 ) | ( n2431 & n2579 ) | ( n2516 & n2579 ) ;
  assign n2581 = ( n2431 & ~n2516 ) | ( n2431 & n2579 ) | ( ~n2516 & n2579 ) ;
  assign n2582 = ( n2516 & ~n2580 ) | ( n2516 & n2581 ) | ( ~n2580 & n2581 ) ;
  assign n2583 = ( n2482 & ~n2485 ) | ( n2482 & n2582 ) | ( ~n2485 & n2582 ) ;
  assign n2584 = ( n2482 & n2485 ) | ( n2482 & n2582 ) | ( n2485 & n2582 ) ;
  assign n2585 = ( n2485 & n2583 ) | ( n2485 & ~n2584 ) | ( n2583 & ~n2584 ) ;
  assign n2586 = ( n2527 & ~n2542 ) | ( n2527 & n2569 ) | ( ~n2542 & n2569 ) ;
  assign n2587 = ( n2527 & n2542 ) | ( n2527 & n2569 ) | ( n2542 & n2569 ) ;
  assign n2588 = ( n2542 & n2586 ) | ( n2542 & ~n2587 ) | ( n2586 & ~n2587 ) ;
  assign n2589 = ( n2495 & n2506 ) | ( n2495 & n2588 ) | ( n2506 & n2588 ) ;
  assign n2590 = ( n2495 & n2506 ) | ( n2495 & ~n2588 ) | ( n2506 & ~n2588 ) ;
  assign n2591 = ( n2588 & ~n2589 ) | ( n2588 & n2590 ) | ( ~n2589 & n2590 ) ;
  assign n2592 = ( ~n2498 & n2508 ) | ( ~n2498 & n2591 ) | ( n2508 & n2591 ) ;
  assign n2593 = ( n2498 & n2508 ) | ( n2498 & n2591 ) | ( n2508 & n2591 ) ;
  assign n2594 = ( n2498 & n2592 ) | ( n2498 & ~n2593 ) | ( n2592 & ~n2593 ) ;
  assign n2595 = x24 & x26 ;
  assign n2596 = x1 & x49 ;
  assign n2597 = n2595 | n2596 ;
  assign n2598 = x26 & x49 ;
  assign n2599 = n695 & n2598 ;
  assign n2600 = n2597 & ~n2599 ;
  assign n2601 = ( n2548 & ~n2557 ) | ( n2548 & n2600 ) | ( ~n2557 & n2600 ) ;
  assign n2602 = ( n2548 & n2557 ) | ( n2548 & n2600 ) | ( n2557 & n2600 ) ;
  assign n2603 = ( n2557 & n2601 ) | ( n2557 & ~n2602 ) | ( n2601 & ~n2602 ) ;
  assign n2604 = ( ~n2530 & n2572 ) | ( ~n2530 & n2603 ) | ( n2572 & n2603 ) ;
  assign n2605 = ( n2530 & n2572 ) | ( n2530 & n2603 ) | ( n2572 & n2603 ) ;
  assign n2606 = ( n2530 & n2604 ) | ( n2530 & ~n2605 ) | ( n2604 & ~n2605 ) ;
  assign n2607 = ( n2521 & ~n2536 ) | ( n2521 & n2563 ) | ( ~n2536 & n2563 ) ;
  assign n2608 = ( n2521 & n2536 ) | ( n2521 & n2563 ) | ( n2536 & n2563 ) ;
  assign n2609 = ( n2536 & n2607 ) | ( n2536 & ~n2608 ) | ( n2607 & ~n2608 ) ;
  assign n2610 = ( n2488 & n2551 ) | ( n2488 & n2609 ) | ( n2551 & n2609 ) ;
  assign n2611 = ( ~n2488 & n2551 ) | ( ~n2488 & n2609 ) | ( n2551 & n2609 ) ;
  assign n2612 = ( n2488 & ~n2610 ) | ( n2488 & n2611 ) | ( ~n2610 & n2611 ) ;
  assign n2613 = ( ~n2575 & n2606 ) | ( ~n2575 & n2612 ) | ( n2606 & n2612 ) ;
  assign n2614 = ( n2575 & n2606 ) | ( n2575 & n2612 ) | ( n2606 & n2612 ) ;
  assign n2615 = ( n2575 & n2613 ) | ( n2575 & ~n2614 ) | ( n2613 & ~n2614 ) ;
  assign n2616 = ( ~n2578 & n2594 ) | ( ~n2578 & n2615 ) | ( n2594 & n2615 ) ;
  assign n2617 = ( n2578 & n2594 ) | ( n2578 & n2615 ) | ( n2594 & n2615 ) ;
  assign n2618 = ( n2578 & n2616 ) | ( n2578 & ~n2617 ) | ( n2616 & ~n2617 ) ;
  assign n2619 = ( n2394 & n2444 ) | ( n2394 & ~n2504 ) | ( n2444 & ~n2504 ) ;
  assign n2620 = x23 & x27 ;
  assign n2621 = x18 & x32 ;
  assign n2622 = x22 & x28 ;
  assign n2623 = ( ~n2620 & n2621 ) | ( ~n2620 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2624 = ( n2620 & n2621 ) | ( n2620 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2625 = ( n2620 & n2623 ) | ( n2620 & ~n2624 ) | ( n2623 & ~n2624 ) ;
  assign n2626 = x16 & x34 ;
  assign n2627 = x15 & x35 ;
  assign n2628 = x5 & x45 ;
  assign n2629 = ( ~n2626 & n2627 ) | ( ~n2626 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2630 = ( n2626 & n2627 ) | ( n2626 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2631 = ( n2626 & n2629 ) | ( n2626 & ~n2630 ) | ( n2629 & ~n2630 ) ;
  assign n2632 = ( ~n2619 & n2625 ) | ( ~n2619 & n2631 ) | ( n2625 & n2631 ) ;
  assign n2633 = ( n2619 & n2625 ) | ( n2619 & n2631 ) | ( n2625 & n2631 ) ;
  assign n2634 = ( n2619 & n2632 ) | ( n2619 & ~n2633 ) | ( n2632 & ~n2633 ) ;
  assign n2635 = ( x2 & ~x48 ) | ( x2 & n782 ) | ( ~x48 & n782 ) ;
  assign n2636 = x0 & x50 ;
  assign n2637 = x2 | n782 ;
  assign n2638 = ( ~n2635 & n2636 ) | ( ~n2635 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2639 = ( n2635 & n2636 ) | ( n2635 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2640 = ( n2635 & n2638 ) | ( n2635 & ~n2639 ) | ( n2638 & ~n2639 ) ;
  assign n2641 = x4 & x46 ;
  assign n2642 = x3 & x47 ;
  assign n2643 = x17 & x33 ;
  assign n2644 = ( ~n2641 & n2642 ) | ( ~n2641 & n2643 ) | ( n2642 & n2643 ) ;
  assign n2645 = ( n2641 & n2642 ) | ( n2641 & n2643 ) | ( n2642 & n2643 ) ;
  assign n2646 = ( n2641 & n2644 ) | ( n2641 & ~n2645 ) | ( n2644 & ~n2645 ) ;
  assign n2647 = x19 & x31 ;
  assign n2648 = x20 & x30 ;
  assign n2649 = x21 & x29 ;
  assign n2650 = ( ~n2647 & n2648 ) | ( ~n2647 & n2649 ) | ( n2648 & n2649 ) ;
  assign n2651 = ( n2647 & n2648 ) | ( n2647 & n2649 ) | ( n2648 & n2649 ) ;
  assign n2652 = ( n2647 & n2650 ) | ( n2647 & ~n2651 ) | ( n2650 & ~n2651 ) ;
  assign n2653 = ( ~n2640 & n2646 ) | ( ~n2640 & n2652 ) | ( n2646 & n2652 ) ;
  assign n2654 = ( n2640 & n2646 ) | ( n2640 & n2652 ) | ( n2646 & n2652 ) ;
  assign n2655 = ( n2640 & n2653 ) | ( n2640 & ~n2654 ) | ( n2653 & ~n2654 ) ;
  assign n2656 = x13 & x37 ;
  assign n2657 = x9 & x41 ;
  assign n2658 = x8 & x42 ;
  assign n2659 = ( ~n2656 & n2657 ) | ( ~n2656 & n2658 ) | ( n2657 & n2658 ) ;
  assign n2660 = ( n2656 & n2657 ) | ( n2656 & n2658 ) | ( n2657 & n2658 ) ;
  assign n2661 = ( n2656 & n2659 ) | ( n2656 & ~n2660 ) | ( n2659 & ~n2660 ) ;
  assign n2662 = x11 & x39 ;
  assign n2663 = x10 & x40 ;
  assign n2664 = x12 & x38 ;
  assign n2665 = ( ~n2662 & n2663 ) | ( ~n2662 & n2664 ) | ( n2663 & n2664 ) ;
  assign n2666 = ( n2662 & n2663 ) | ( n2662 & n2664 ) | ( n2663 & n2664 ) ;
  assign n2667 = ( n2662 & n2665 ) | ( n2662 & ~n2666 ) | ( n2665 & ~n2666 ) ;
  assign n2668 = x14 & x36 ;
  assign n2669 = x6 & x44 ;
  assign n2670 = x7 & x43 ;
  assign n2671 = ( ~n2668 & n2669 ) | ( ~n2668 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2672 = ( n2668 & n2669 ) | ( n2668 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2673 = ( n2668 & n2671 ) | ( n2668 & ~n2672 ) | ( n2671 & ~n2672 ) ;
  assign n2674 = ( ~n2661 & n2667 ) | ( ~n2661 & n2673 ) | ( n2667 & n2673 ) ;
  assign n2675 = ( n2661 & n2667 ) | ( n2661 & n2673 ) | ( n2667 & n2673 ) ;
  assign n2676 = ( n2661 & n2674 ) | ( n2661 & ~n2675 ) | ( n2674 & ~n2675 ) ;
  assign n2677 = ( ~n2634 & n2655 ) | ( ~n2634 & n2676 ) | ( n2655 & n2676 ) ;
  assign n2678 = ( n2634 & n2655 ) | ( n2634 & n2676 ) | ( n2655 & n2676 ) ;
  assign n2679 = ( n2634 & n2677 ) | ( n2634 & ~n2678 ) | ( n2677 & ~n2678 ) ;
  assign n2680 = ( n2491 & n2511 ) | ( n2491 & ~n2679 ) | ( n2511 & ~n2679 ) ;
  assign n2681 = ( n2491 & n2511 ) | ( n2491 & n2679 ) | ( n2511 & n2679 ) ;
  assign n2682 = ( n2679 & n2680 ) | ( n2679 & ~n2681 ) | ( n2680 & ~n2681 ) ;
  assign n2683 = ( n2514 & n2618 ) | ( n2514 & n2682 ) | ( n2618 & n2682 ) ;
  assign n2684 = ( n2514 & ~n2618 ) | ( n2514 & n2682 ) | ( ~n2618 & n2682 ) ;
  assign n2685 = ( n2618 & ~n2683 ) | ( n2618 & n2684 ) | ( ~n2683 & n2684 ) ;
  assign n2686 = ( n2580 & n2584 ) | ( n2580 & n2685 ) | ( n2584 & n2685 ) ;
  assign n2687 = ( n2580 & ~n2584 ) | ( n2580 & n2685 ) | ( ~n2584 & n2685 ) ;
  assign n2688 = ( n2584 & ~n2686 ) | ( n2584 & n2687 ) | ( ~n2686 & n2687 ) ;
  assign n2689 = x7 & x44 ;
  assign n2690 = x13 & x38 ;
  assign n2691 = x8 & x43 ;
  assign n2692 = ( ~n2689 & n2690 ) | ( ~n2689 & n2691 ) | ( n2690 & n2691 ) ;
  assign n2693 = ( n2689 & n2690 ) | ( n2689 & n2691 ) | ( n2690 & n2691 ) ;
  assign n2694 = ( n2689 & n2692 ) | ( n2689 & ~n2693 ) | ( n2692 & ~n2693 ) ;
  assign n2695 = x9 & x42 ;
  assign n2696 = x10 & x41 ;
  assign n2697 = x12 & x39 ;
  assign n2698 = ( ~n2695 & n2696 ) | ( ~n2695 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2699 = ( n2695 & n2696 ) | ( n2695 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2700 = ( n2695 & n2698 ) | ( n2695 & ~n2699 ) | ( n2698 & ~n2699 ) ;
  assign n2701 = x25 & x26 ;
  assign n2702 = x24 & x27 ;
  assign n2703 = x11 & x40 ;
  assign n2704 = ( ~n2701 & n2702 ) | ( ~n2701 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2705 = ( n2701 & n2702 ) | ( n2701 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2706 = ( n2701 & n2704 ) | ( n2701 & ~n2705 ) | ( n2704 & ~n2705 ) ;
  assign n2707 = ( ~n2694 & n2700 ) | ( ~n2694 & n2706 ) | ( n2700 & n2706 ) ;
  assign n2708 = ( n2694 & n2700 ) | ( n2694 & n2706 ) | ( n2700 & n2706 ) ;
  assign n2709 = ( n2694 & n2707 ) | ( n2694 & ~n2708 ) | ( n2707 & ~n2708 ) ;
  assign n2710 = x21 & x30 ;
  assign n2711 = x22 & x29 ;
  assign n2712 = x23 & x28 ;
  assign n2713 = ( ~n2710 & n2711 ) | ( ~n2710 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2714 = ( n2710 & n2711 ) | ( n2710 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2715 = ( n2710 & n2713 ) | ( n2710 & ~n2714 ) | ( n2713 & ~n2714 ) ;
  assign n2716 = x5 & x46 ;
  assign n2717 = x16 & x35 ;
  assign n2718 = ( ~n1279 & n2716 ) | ( ~n1279 & n2717 ) | ( n2716 & n2717 ) ;
  assign n2719 = ( n1279 & n2716 ) | ( n1279 & n2717 ) | ( n2716 & n2717 ) ;
  assign n2720 = ( n1279 & n2718 ) | ( n1279 & ~n2719 ) | ( n2718 & ~n2719 ) ;
  assign n2721 = x6 & x45 ;
  assign n2722 = x14 & x37 ;
  assign n2723 = x15 & x36 ;
  assign n2724 = ( ~n2721 & n2722 ) | ( ~n2721 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2725 = ( n2721 & n2722 ) | ( n2721 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2726 = ( n2721 & n2724 ) | ( n2721 & ~n2725 ) | ( n2724 & ~n2725 ) ;
  assign n2727 = ( ~n2715 & n2720 ) | ( ~n2715 & n2726 ) | ( n2720 & n2726 ) ;
  assign n2728 = ( n2715 & n2720 ) | ( n2715 & n2726 ) | ( n2720 & n2726 ) ;
  assign n2729 = ( n2715 & n2727 ) | ( n2715 & ~n2728 ) | ( n2727 & ~n2728 ) ;
  assign n2730 = x1 & x50 ;
  assign n2731 = x26 & x50 ;
  assign n2732 = ( n2599 & n2730 ) | ( n2599 & ~n2731 ) | ( n2730 & ~n2731 ) ;
  assign n2733 = x26 & ~n2730 ;
  assign n2734 = x0 & x51 ;
  assign n2735 = ( n2732 & n2733 ) | ( n2732 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2736 = ( ~n2732 & n2733 ) | ( ~n2732 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2737 = ( n2732 & ~n2735 ) | ( n2732 & n2736 ) | ( ~n2735 & n2736 ) ;
  assign n2738 = x20 & x31 ;
  assign n2739 = x19 & x32 ;
  assign n2740 = x17 & x34 ;
  assign n2741 = ( ~n2738 & n2739 ) | ( ~n2738 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2742 = ( n2738 & n2739 ) | ( n2738 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2743 = ( n2738 & n2741 ) | ( n2738 & ~n2742 ) | ( n2741 & ~n2742 ) ;
  assign n2744 = ( n2608 & n2737 ) | ( n2608 & n2743 ) | ( n2737 & n2743 ) ;
  assign n2745 = ( ~n2608 & n2737 ) | ( ~n2608 & n2743 ) | ( n2737 & n2743 ) ;
  assign n2746 = ( n2608 & ~n2744 ) | ( n2608 & n2745 ) | ( ~n2744 & n2745 ) ;
  assign n2747 = ( ~n2709 & n2729 ) | ( ~n2709 & n2746 ) | ( n2729 & n2746 ) ;
  assign n2748 = ( n2709 & n2729 ) | ( n2709 & n2746 ) | ( n2729 & n2746 ) ;
  assign n2749 = ( n2709 & n2747 ) | ( n2709 & ~n2748 ) | ( n2747 & ~n2748 ) ;
  assign n2750 = ( n2593 & ~n2614 ) | ( n2593 & n2749 ) | ( ~n2614 & n2749 ) ;
  assign n2751 = ( n2593 & n2614 ) | ( n2593 & n2749 ) | ( n2614 & n2749 ) ;
  assign n2752 = ( n2614 & n2750 ) | ( n2614 & ~n2751 ) | ( n2750 & ~n2751 ) ;
  assign n2753 = x3 & x48 ;
  assign n2754 = x4 & x47 ;
  assign n2755 = x2 & x49 ;
  assign n2756 = ( ~n2753 & n2754 ) | ( ~n2753 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2757 = ( n2753 & n2754 ) | ( n2753 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2758 = ( n2753 & n2756 ) | ( n2753 & ~n2757 ) | ( n2756 & ~n2757 ) ;
  assign n2759 = ( n2630 & n2666 ) | ( n2630 & ~n2758 ) | ( n2666 & ~n2758 ) ;
  assign n2760 = ( n2630 & n2666 ) | ( n2630 & n2758 ) | ( n2666 & n2758 ) ;
  assign n2761 = ( n2758 & n2759 ) | ( n2758 & ~n2760 ) | ( n2759 & ~n2760 ) ;
  assign n2762 = ( n2589 & n2633 ) | ( n2589 & n2761 ) | ( n2633 & n2761 ) ;
  assign n2763 = ( n2589 & n2633 ) | ( n2589 & ~n2761 ) | ( n2633 & ~n2761 ) ;
  assign n2764 = ( n2761 & ~n2762 ) | ( n2761 & n2763 ) | ( ~n2762 & n2763 ) ;
  assign n2765 = ( x2 & n782 ) | ( x2 & n2636 ) | ( n782 & n2636 ) ;
  assign n2766 = x48 & n2765 ;
  assign n2767 = ( n2645 & n2651 ) | ( n2645 & n2766 ) | ( n2651 & n2766 ) ;
  assign n2768 = ( n2645 & n2651 ) | ( n2645 & ~n2766 ) | ( n2651 & ~n2766 ) ;
  assign n2769 = ( n2766 & ~n2767 ) | ( n2766 & n2768 ) | ( ~n2767 & n2768 ) ;
  assign n2770 = ( n2624 & ~n2660 ) | ( n2624 & n2672 ) | ( ~n2660 & n2672 ) ;
  assign n2771 = ( n2624 & n2660 ) | ( n2624 & n2672 ) | ( n2660 & n2672 ) ;
  assign n2772 = ( n2660 & n2770 ) | ( n2660 & ~n2771 ) | ( n2770 & ~n2771 ) ;
  assign n2773 = ( n2675 & n2769 ) | ( n2675 & n2772 ) | ( n2769 & n2772 ) ;
  assign n2774 = ( n2675 & ~n2769 ) | ( n2675 & n2772 ) | ( ~n2769 & n2772 ) ;
  assign n2775 = ( n2769 & ~n2773 ) | ( n2769 & n2774 ) | ( ~n2773 & n2774 ) ;
  assign n2776 = ( n2678 & n2764 ) | ( n2678 & n2775 ) | ( n2764 & n2775 ) ;
  assign n2777 = ( n2678 & ~n2764 ) | ( n2678 & n2775 ) | ( ~n2764 & n2775 ) ;
  assign n2778 = ( n2764 & ~n2776 ) | ( n2764 & n2777 ) | ( ~n2776 & n2777 ) ;
  assign n2779 = ( n2587 & n2602 ) | ( n2587 & ~n2654 ) | ( n2602 & ~n2654 ) ;
  assign n2780 = ( n2587 & n2602 ) | ( n2587 & n2654 ) | ( n2602 & n2654 ) ;
  assign n2781 = ( n2654 & n2779 ) | ( n2654 & ~n2780 ) | ( n2779 & ~n2780 ) ;
  assign n2782 = ( n2605 & n2610 ) | ( n2605 & n2781 ) | ( n2610 & n2781 ) ;
  assign n2783 = ( n2605 & ~n2610 ) | ( n2605 & n2781 ) | ( ~n2610 & n2781 ) ;
  assign n2784 = ( n2610 & ~n2782 ) | ( n2610 & n2783 ) | ( ~n2782 & n2783 ) ;
  assign n2785 = ( ~n2681 & n2778 ) | ( ~n2681 & n2784 ) | ( n2778 & n2784 ) ;
  assign n2786 = ( n2681 & n2778 ) | ( n2681 & n2784 ) | ( n2778 & n2784 ) ;
  assign n2787 = ( n2681 & n2785 ) | ( n2681 & ~n2786 ) | ( n2785 & ~n2786 ) ;
  assign n2788 = ( n2617 & ~n2752 ) | ( n2617 & n2787 ) | ( ~n2752 & n2787 ) ;
  assign n2789 = ( n2617 & n2752 ) | ( n2617 & n2787 ) | ( n2752 & n2787 ) ;
  assign n2790 = ( n2752 & n2788 ) | ( n2752 & ~n2789 ) | ( n2788 & ~n2789 ) ;
  assign n2791 = ( n2683 & n2686 ) | ( n2683 & n2790 ) | ( n2686 & n2790 ) ;
  assign n2792 = ( n2683 & ~n2686 ) | ( n2683 & n2790 ) | ( ~n2686 & n2790 ) ;
  assign n2793 = ( n2686 & ~n2791 ) | ( n2686 & n2792 ) | ( ~n2791 & n2792 ) ;
  assign n2794 = x5 & x47 ;
  assign n2795 = x16 & x36 ;
  assign n2796 = x6 & x46 ;
  assign n2797 = ( ~n2794 & n2795 ) | ( ~n2794 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2798 = ( n2794 & n2795 ) | ( n2794 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2799 = ( n2794 & n2797 ) | ( n2794 & ~n2798 ) | ( n2797 & ~n2798 ) ;
  assign n2800 = x7 & x45 ;
  assign n2801 = x8 & x44 ;
  assign n2802 = x15 & x37 ;
  assign n2803 = ( ~n2800 & n2801 ) | ( ~n2800 & n2802 ) | ( n2801 & n2802 ) ;
  assign n2804 = ( n2800 & n2801 ) | ( n2800 & n2802 ) | ( n2801 & n2802 ) ;
  assign n2805 = ( n2800 & n2803 ) | ( n2800 & ~n2804 ) | ( n2803 & ~n2804 ) ;
  assign n2806 = x11 & x41 ;
  assign n2807 = x10 & x42 ;
  assign n2808 = x12 & x40 ;
  assign n2809 = ( ~n2806 & n2807 ) | ( ~n2806 & n2808 ) | ( n2807 & n2808 ) ;
  assign n2810 = ( n2806 & n2807 ) | ( n2806 & n2808 ) | ( n2807 & n2808 ) ;
  assign n2811 = ( n2806 & n2809 ) | ( n2806 & ~n2810 ) | ( n2809 & ~n2810 ) ;
  assign n2812 = ( ~n2799 & n2805 ) | ( ~n2799 & n2811 ) | ( n2805 & n2811 ) ;
  assign n2813 = ( n2799 & n2805 ) | ( n2799 & n2811 ) | ( n2805 & n2811 ) ;
  assign n2814 = ( n2799 & n2812 ) | ( n2799 & ~n2813 ) | ( n2812 & ~n2813 ) ;
  assign n2815 = x21 & x31 ;
  assign n2816 = x20 & x32 ;
  assign n2817 = ( ~n1349 & n2815 ) | ( ~n1349 & n2816 ) | ( n2815 & n2816 ) ;
  assign n2818 = ( n1349 & n2815 ) | ( n1349 & n2816 ) | ( n2815 & n2816 ) ;
  assign n2819 = ( n1349 & n2817 ) | ( n1349 & ~n2818 ) | ( n2817 & ~n2818 ) ;
  assign n2820 = x24 & x28 ;
  assign n2821 = x22 & x30 ;
  assign n2822 = x23 & x29 ;
  assign n2823 = ( ~n2820 & n2821 ) | ( ~n2820 & n2822 ) | ( n2821 & n2822 ) ;
  assign n2824 = ( n2820 & n2821 ) | ( n2820 & n2822 ) | ( n2821 & n2822 ) ;
  assign n2825 = ( n2820 & n2823 ) | ( n2820 & ~n2824 ) | ( n2823 & ~n2824 ) ;
  assign n2826 = x13 & x39 ;
  assign n2827 = x14 & x38 ;
  assign n2828 = x9 & x43 ;
  assign n2829 = ( ~n2826 & n2827 ) | ( ~n2826 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2830 = ( n2826 & n2827 ) | ( n2826 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2831 = ( n2826 & n2829 ) | ( n2826 & ~n2830 ) | ( n2829 & ~n2830 ) ;
  assign n2832 = ( ~n2819 & n2825 ) | ( ~n2819 & n2831 ) | ( n2825 & n2831 ) ;
  assign n2833 = ( n2819 & n2825 ) | ( n2819 & n2831 ) | ( n2825 & n2831 ) ;
  assign n2834 = ( n2819 & n2832 ) | ( n2819 & ~n2833 ) | ( n2832 & ~n2833 ) ;
  assign n2835 = ( n2773 & n2814 ) | ( n2773 & n2834 ) | ( n2814 & n2834 ) ;
  assign n2836 = ( ~n2773 & n2814 ) | ( ~n2773 & n2834 ) | ( n2814 & n2834 ) ;
  assign n2837 = ( n2773 & ~n2835 ) | ( n2773 & n2836 ) | ( ~n2835 & n2836 ) ;
  assign n2838 = ( n2776 & n2782 ) | ( n2776 & n2837 ) | ( n2782 & n2837 ) ;
  assign n2839 = ( n2776 & n2782 ) | ( n2776 & ~n2837 ) | ( n2782 & ~n2837 ) ;
  assign n2840 = ( n2837 & ~n2838 ) | ( n2837 & n2839 ) | ( ~n2838 & n2839 ) ;
  assign n2841 = x25 & x27 ;
  assign n2842 = x1 & x51 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = x27 & x51 ;
  assign n2845 = n782 & n2844 ;
  assign n2846 = n2843 & ~n2845 ;
  assign n2847 = x50 & n820 ;
  assign n2848 = ( n2705 & ~n2846 ) | ( n2705 & n2847 ) | ( ~n2846 & n2847 ) ;
  assign n2849 = ( n2705 & n2846 ) | ( n2705 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2850 = ( n2846 & n2848 ) | ( n2846 & ~n2849 ) | ( n2848 & ~n2849 ) ;
  assign n2851 = ( n2708 & n2760 ) | ( n2708 & n2850 ) | ( n2760 & n2850 ) ;
  assign n2852 = ( n2708 & ~n2760 ) | ( n2708 & n2850 ) | ( ~n2760 & n2850 ) ;
  assign n2853 = ( n2760 & ~n2851 ) | ( n2760 & n2852 ) | ( ~n2851 & n2852 ) ;
  assign n2854 = x2 & x50 ;
  assign n2855 = x19 & x33 ;
  assign n2856 = x3 & x49 ;
  assign n2857 = ( ~n2854 & n2855 ) | ( ~n2854 & n2856 ) | ( n2855 & n2856 ) ;
  assign n2858 = ( n2854 & n2855 ) | ( n2854 & n2856 ) | ( n2855 & n2856 ) ;
  assign n2859 = ( n2854 & n2857 ) | ( n2854 & ~n2858 ) | ( n2857 & ~n2858 ) ;
  assign n2860 = ( ~n2767 & n2771 ) | ( ~n2767 & n2859 ) | ( n2771 & n2859 ) ;
  assign n2861 = ( n2767 & n2771 ) | ( n2767 & n2859 ) | ( n2771 & n2859 ) ;
  assign n2862 = ( n2767 & n2860 ) | ( n2767 & ~n2861 ) | ( n2860 & ~n2861 ) ;
  assign n2863 = ( n2762 & ~n2853 ) | ( n2762 & n2862 ) | ( ~n2853 & n2862 ) ;
  assign n2864 = ( n2762 & n2853 ) | ( n2762 & n2862 ) | ( n2853 & n2862 ) ;
  assign n2865 = ( n2853 & n2863 ) | ( n2853 & ~n2864 ) | ( n2863 & ~n2864 ) ;
  assign n2866 = x0 & x52 ;
  assign n2867 = x4 & x48 ;
  assign n2868 = ( ~n1372 & n2866 ) | ( ~n1372 & n2867 ) | ( n2866 & n2867 ) ;
  assign n2869 = ( n1372 & n2866 ) | ( n1372 & n2867 ) | ( n2866 & n2867 ) ;
  assign n2870 = ( n1372 & n2868 ) | ( n1372 & ~n2869 ) | ( n2868 & ~n2869 ) ;
  assign n2871 = ( n2699 & ~n2735 ) | ( n2699 & n2870 ) | ( ~n2735 & n2870 ) ;
  assign n2872 = ( n2699 & n2735 ) | ( n2699 & n2870 ) | ( n2735 & n2870 ) ;
  assign n2873 = ( n2735 & n2871 ) | ( n2735 & ~n2872 ) | ( n2871 & ~n2872 ) ;
  assign n2874 = ( n2744 & ~n2780 ) | ( n2744 & n2873 ) | ( ~n2780 & n2873 ) ;
  assign n2875 = ( n2744 & n2780 ) | ( n2744 & n2873 ) | ( n2780 & n2873 ) ;
  assign n2876 = ( n2780 & n2874 ) | ( n2780 & ~n2875 ) | ( n2874 & ~n2875 ) ;
  assign n2877 = ( n2725 & n2742 ) | ( n2725 & ~n2757 ) | ( n2742 & ~n2757 ) ;
  assign n2878 = ( n2725 & n2742 ) | ( n2725 & n2757 ) | ( n2742 & n2757 ) ;
  assign n2879 = ( n2757 & n2877 ) | ( n2757 & ~n2878 ) | ( n2877 & ~n2878 ) ;
  assign n2880 = ( ~n2693 & n2714 ) | ( ~n2693 & n2719 ) | ( n2714 & n2719 ) ;
  assign n2881 = ( n2693 & n2714 ) | ( n2693 & n2719 ) | ( n2714 & n2719 ) ;
  assign n2882 = ( n2693 & n2880 ) | ( n2693 & ~n2881 ) | ( n2880 & ~n2881 ) ;
  assign n2883 = ( n2728 & n2879 ) | ( n2728 & n2882 ) | ( n2879 & n2882 ) ;
  assign n2884 = ( ~n2728 & n2879 ) | ( ~n2728 & n2882 ) | ( n2879 & n2882 ) ;
  assign n2885 = ( n2728 & ~n2883 ) | ( n2728 & n2884 ) | ( ~n2883 & n2884 ) ;
  assign n2886 = ( n2748 & n2876 ) | ( n2748 & n2885 ) | ( n2876 & n2885 ) ;
  assign n2887 = ( n2748 & ~n2876 ) | ( n2748 & n2885 ) | ( ~n2876 & n2885 ) ;
  assign n2888 = ( n2876 & ~n2886 ) | ( n2876 & n2887 ) | ( ~n2886 & n2887 ) ;
  assign n2889 = ( n2751 & ~n2865 ) | ( n2751 & n2888 ) | ( ~n2865 & n2888 ) ;
  assign n2890 = ( n2751 & n2865 ) | ( n2751 & n2888 ) | ( n2865 & n2888 ) ;
  assign n2891 = ( n2865 & n2889 ) | ( n2865 & ~n2890 ) | ( n2889 & ~n2890 ) ;
  assign n2892 = ( n2786 & n2840 ) | ( n2786 & n2891 ) | ( n2840 & n2891 ) ;
  assign n2893 = ( n2786 & ~n2840 ) | ( n2786 & n2891 ) | ( ~n2840 & n2891 ) ;
  assign n2894 = ( n2840 & ~n2892 ) | ( n2840 & n2893 ) | ( ~n2892 & n2893 ) ;
  assign n2895 = ( n2789 & n2791 ) | ( n2789 & n2894 ) | ( n2791 & n2894 ) ;
  assign n2896 = ( n2789 & ~n2791 ) | ( n2789 & n2894 ) | ( ~n2791 & n2894 ) ;
  assign n2897 = ( n2791 & ~n2895 ) | ( n2791 & n2896 ) | ( ~n2895 & n2896 ) ;
  assign n2898 = ( ~n2824 & n2858 ) | ( ~n2824 & n2869 ) | ( n2858 & n2869 ) ;
  assign n2899 = ( n2824 & n2858 ) | ( n2824 & n2869 ) | ( n2858 & n2869 ) ;
  assign n2900 = ( n2824 & n2898 ) | ( n2824 & ~n2899 ) | ( n2898 & ~n2899 ) ;
  assign n2901 = ( n2833 & n2872 ) | ( n2833 & n2900 ) | ( n2872 & n2900 ) ;
  assign n2902 = ( n2833 & ~n2872 ) | ( n2833 & n2900 ) | ( ~n2872 & n2900 ) ;
  assign n2903 = ( n2872 & ~n2901 ) | ( n2872 & n2902 ) | ( ~n2901 & n2902 ) ;
  assign n2904 = ~x1 & x27 ;
  assign n2905 = ( x1 & x27 ) | ( x1 & x52 ) | ( x27 & x52 ) ;
  assign n2906 = x27 & x52 ;
  assign n2907 = ( n2904 & n2905 ) | ( n2904 & ~n2906 ) | ( n2905 & ~n2906 ) ;
  assign n2908 = ( n2810 & n2830 ) | ( n2810 & ~n2907 ) | ( n2830 & ~n2907 ) ;
  assign n2909 = ( n2810 & n2830 ) | ( n2810 & n2907 ) | ( n2830 & n2907 ) ;
  assign n2910 = ( n2907 & n2908 ) | ( n2907 & ~n2909 ) | ( n2908 & ~n2909 ) ;
  assign n2911 = ( n2798 & ~n2804 ) | ( n2798 & n2818 ) | ( ~n2804 & n2818 ) ;
  assign n2912 = ( n2798 & n2804 ) | ( n2798 & n2818 ) | ( n2804 & n2818 ) ;
  assign n2913 = ( n2804 & n2911 ) | ( n2804 & ~n2912 ) | ( n2911 & ~n2912 ) ;
  assign n2914 = ( n2813 & n2910 ) | ( n2813 & n2913 ) | ( n2910 & n2913 ) ;
  assign n2915 = ( n2813 & ~n2910 ) | ( n2813 & n2913 ) | ( ~n2910 & n2913 ) ;
  assign n2916 = ( n2910 & ~n2914 ) | ( n2910 & n2915 ) | ( ~n2914 & n2915 ) ;
  assign n2917 = ( n2864 & ~n2903 ) | ( n2864 & n2916 ) | ( ~n2903 & n2916 ) ;
  assign n2918 = ( n2864 & n2903 ) | ( n2864 & n2916 ) | ( n2903 & n2916 ) ;
  assign n2919 = ( n2903 & n2917 ) | ( n2903 & ~n2918 ) | ( n2917 & ~n2918 ) ;
  assign n2920 = ( n2849 & ~n2878 ) | ( n2849 & n2881 ) | ( ~n2878 & n2881 ) ;
  assign n2921 = ( n2849 & n2878 ) | ( n2849 & n2881 ) | ( n2878 & n2881 ) ;
  assign n2922 = ( n2878 & n2920 ) | ( n2878 & ~n2921 ) | ( n2920 & ~n2921 ) ;
  assign n2923 = ( n2835 & n2875 ) | ( n2835 & n2922 ) | ( n2875 & n2922 ) ;
  assign n2924 = ( ~n2835 & n2875 ) | ( ~n2835 & n2922 ) | ( n2875 & n2922 ) ;
  assign n2925 = ( n2835 & ~n2923 ) | ( n2835 & n2924 ) | ( ~n2923 & n2924 ) ;
  assign n2926 = ( n2838 & n2919 ) | ( n2838 & n2925 ) | ( n2919 & n2925 ) ;
  assign n2927 = ( ~n2838 & n2919 ) | ( ~n2838 & n2925 ) | ( n2919 & n2925 ) ;
  assign n2928 = ( n2838 & ~n2926 ) | ( n2838 & n2927 ) | ( ~n2926 & n2927 ) ;
  assign n2929 = x2 & x51 ;
  assign n2930 = x3 & x50 ;
  assign n2931 = ( ~n2845 & n2929 ) | ( ~n2845 & n2930 ) | ( n2929 & n2930 ) ;
  assign n2932 = ( n2845 & n2929 ) | ( n2845 & n2930 ) | ( n2929 & n2930 ) ;
  assign n2933 = ( n2845 & n2931 ) | ( n2845 & ~n2932 ) | ( n2931 & ~n2932 ) ;
  assign n2934 = x20 & x33 ;
  assign n2935 = x19 & x34 ;
  assign n2936 = x21 & x32 ;
  assign n2937 = ( ~n2934 & n2935 ) | ( ~n2934 & n2936 ) | ( n2935 & n2936 ) ;
  assign n2938 = ( n2934 & n2935 ) | ( n2934 & n2936 ) | ( n2935 & n2936 ) ;
  assign n2939 = ( n2934 & n2937 ) | ( n2934 & ~n2938 ) | ( n2937 & ~n2938 ) ;
  assign n2940 = x4 & x49 ;
  assign n2941 = x18 & x35 ;
  assign n2942 = x17 & x36 ;
  assign n2943 = ( ~n2940 & n2941 ) | ( ~n2940 & n2942 ) | ( n2941 & n2942 ) ;
  assign n2944 = ( n2940 & n2941 ) | ( n2940 & n2942 ) | ( n2941 & n2942 ) ;
  assign n2945 = ( n2940 & n2943 ) | ( n2940 & ~n2944 ) | ( n2943 & ~n2944 ) ;
  assign n2946 = ( ~n2933 & n2939 ) | ( ~n2933 & n2945 ) | ( n2939 & n2945 ) ;
  assign n2947 = ( n2933 & n2939 ) | ( n2933 & n2945 ) | ( n2939 & n2945 ) ;
  assign n2948 = ( n2933 & n2946 ) | ( n2933 & ~n2947 ) | ( n2946 & ~n2947 ) ;
  assign n2949 = x9 & x44 ;
  assign n2950 = x8 & x45 ;
  assign n2951 = x14 & x39 ;
  assign n2952 = ( ~n2949 & n2950 ) | ( ~n2949 & n2951 ) | ( n2950 & n2951 ) ;
  assign n2953 = ( n2949 & n2950 ) | ( n2949 & n2951 ) | ( n2950 & n2951 ) ;
  assign n2954 = ( n2949 & n2952 ) | ( n2949 & ~n2953 ) | ( n2952 & ~n2953 ) ;
  assign n2955 = x5 & x48 ;
  assign n2956 = x0 & x53 ;
  assign n2957 = x16 & x37 ;
  assign n2958 = ( ~n2955 & n2956 ) | ( ~n2955 & n2957 ) | ( n2956 & n2957 ) ;
  assign n2959 = ( n2955 & n2956 ) | ( n2955 & n2957 ) | ( n2956 & n2957 ) ;
  assign n2960 = ( n2955 & n2958 ) | ( n2955 & ~n2959 ) | ( n2958 & ~n2959 ) ;
  assign n2961 = x7 & x46 ;
  assign n2962 = x6 & x47 ;
  assign n2963 = x15 & x38 ;
  assign n2964 = ( ~n2961 & n2962 ) | ( ~n2961 & n2963 ) | ( n2962 & n2963 ) ;
  assign n2965 = ( n2961 & n2962 ) | ( n2961 & n2963 ) | ( n2962 & n2963 ) ;
  assign n2966 = ( n2961 & n2964 ) | ( n2961 & ~n2965 ) | ( n2964 & ~n2965 ) ;
  assign n2967 = ( ~n2954 & n2960 ) | ( ~n2954 & n2966 ) | ( n2960 & n2966 ) ;
  assign n2968 = ( n2954 & n2960 ) | ( n2954 & n2966 ) | ( n2960 & n2966 ) ;
  assign n2969 = ( n2954 & n2967 ) | ( n2954 & ~n2968 ) | ( n2967 & ~n2968 ) ;
  assign n2970 = ( n2861 & n2948 ) | ( n2861 & n2969 ) | ( n2948 & n2969 ) ;
  assign n2971 = ( ~n2861 & n2948 ) | ( ~n2861 & n2969 ) | ( n2948 & n2969 ) ;
  assign n2972 = ( n2861 & ~n2970 ) | ( n2861 & n2971 ) | ( ~n2970 & n2971 ) ;
  assign n2973 = x22 & x31 ;
  assign n2974 = x23 & x30 ;
  assign n2975 = x24 & x29 ;
  assign n2976 = ( ~n2973 & n2974 ) | ( ~n2973 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2977 = ( n2973 & n2974 ) | ( n2973 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2978 = ( n2973 & n2976 ) | ( n2973 & ~n2977 ) | ( n2976 & ~n2977 ) ;
  assign n2979 = x12 & x41 ;
  assign n2980 = x10 & x43 ;
  assign n2981 = x13 & x40 ;
  assign n2982 = ( ~n2979 & n2980 ) | ( ~n2979 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2983 = ( n2979 & n2980 ) | ( n2979 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2984 = ( n2979 & n2982 ) | ( n2979 & ~n2983 ) | ( n2982 & ~n2983 ) ;
  assign n2985 = x26 & x27 ;
  assign n2986 = x25 & x28 ;
  assign n2987 = x11 & x42 ;
  assign n2988 = ( ~n2985 & n2986 ) | ( ~n2985 & n2987 ) | ( n2986 & n2987 ) ;
  assign n2989 = ( n2985 & n2986 ) | ( n2985 & n2987 ) | ( n2986 & n2987 ) ;
  assign n2990 = ( n2985 & n2988 ) | ( n2985 & ~n2989 ) | ( n2988 & ~n2989 ) ;
  assign n2991 = ( ~n2978 & n2984 ) | ( ~n2978 & n2990 ) | ( n2984 & n2990 ) ;
  assign n2992 = ( n2978 & n2984 ) | ( n2978 & n2990 ) | ( n2984 & n2990 ) ;
  assign n2993 = ( n2978 & n2991 ) | ( n2978 & ~n2992 ) | ( n2991 & ~n2992 ) ;
  assign n2994 = ( n2851 & n2883 ) | ( n2851 & n2993 ) | ( n2883 & n2993 ) ;
  assign n2995 = ( n2851 & ~n2883 ) | ( n2851 & n2993 ) | ( ~n2883 & n2993 ) ;
  assign n2996 = ( n2883 & ~n2994 ) | ( n2883 & n2995 ) | ( ~n2994 & n2995 ) ;
  assign n2997 = ( n2886 & n2972 ) | ( n2886 & n2996 ) | ( n2972 & n2996 ) ;
  assign n2998 = ( ~n2886 & n2972 ) | ( ~n2886 & n2996 ) | ( n2972 & n2996 ) ;
  assign n2999 = ( n2886 & ~n2997 ) | ( n2886 & n2998 ) | ( ~n2997 & n2998 ) ;
  assign n3000 = ( n2890 & n2928 ) | ( n2890 & n2999 ) | ( n2928 & n2999 ) ;
  assign n3001 = ( n2890 & ~n2928 ) | ( n2890 & n2999 ) | ( ~n2928 & n2999 ) ;
  assign n3002 = ( n2928 & ~n3000 ) | ( n2928 & n3001 ) | ( ~n3000 & n3001 ) ;
  assign n3003 = ( n2892 & ~n2895 ) | ( n2892 & n3002 ) | ( ~n2895 & n3002 ) ;
  assign n3004 = ( n2892 & n2895 ) | ( n2892 & n3002 ) | ( n2895 & n3002 ) ;
  assign n3005 = ( n2895 & n3003 ) | ( n2895 & ~n3004 ) | ( n3003 & ~n3004 ) ;
  assign n3006 = x26 & x28 ;
  assign n3007 = x1 & x53 ;
  assign n3008 = n3006 | n3007 ;
  assign n3009 = x28 & x53 ;
  assign n3010 = n820 & n3009 ;
  assign n3011 = n3008 & ~n3010 ;
  assign n3012 = x52 & n892 ;
  assign n3013 = x0 & x54 ;
  assign n3014 = ( n3011 & n3012 ) | ( n3011 & n3013 ) | ( n3012 & n3013 ) ;
  assign n3015 = ( ~n3011 & n3012 ) | ( ~n3011 & n3013 ) | ( n3012 & n3013 ) ;
  assign n3016 = ( n3011 & ~n3014 ) | ( n3011 & n3015 ) | ( ~n3014 & n3015 ) ;
  assign n3017 = x24 & x30 ;
  assign n3018 = x25 & x29 ;
  assign n3019 = x23 & x31 ;
  assign n3020 = ( ~n3017 & n3018 ) | ( ~n3017 & n3019 ) | ( n3018 & n3019 ) ;
  assign n3021 = ( n3017 & n3018 ) | ( n3017 & n3019 ) | ( n3018 & n3019 ) ;
  assign n3022 = ( n3017 & n3020 ) | ( n3017 & ~n3021 ) | ( n3020 & ~n3021 ) ;
  assign n3023 = x19 & x35 ;
  assign n3024 = x21 & x33 ;
  assign n3025 = x22 & x32 ;
  assign n3026 = ( ~n3023 & n3024 ) | ( ~n3023 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3027 = ( n3023 & n3024 ) | ( n3023 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3028 = ( n3023 & n3026 ) | ( n3023 & ~n3027 ) | ( n3026 & ~n3027 ) ;
  assign n3029 = ( n3016 & n3022 ) | ( n3016 & n3028 ) | ( n3022 & n3028 ) ;
  assign n3030 = ( ~n3016 & n3022 ) | ( ~n3016 & n3028 ) | ( n3022 & n3028 ) ;
  assign n3031 = ( n3016 & ~n3029 ) | ( n3016 & n3030 ) | ( ~n3029 & n3030 ) ;
  assign n3032 = ( ~n2901 & n2914 ) | ( ~n2901 & n3031 ) | ( n2914 & n3031 ) ;
  assign n3033 = ( n2901 & n2914 ) | ( n2901 & n3031 ) | ( n2914 & n3031 ) ;
  assign n3034 = ( n2901 & n3032 ) | ( n2901 & ~n3033 ) | ( n3032 & ~n3033 ) ;
  assign n3035 = ( n2918 & n2923 ) | ( n2918 & ~n3034 ) | ( n2923 & ~n3034 ) ;
  assign n3036 = ( n2918 & n2923 ) | ( n2918 & n3034 ) | ( n2923 & n3034 ) ;
  assign n3037 = ( n3034 & n3035 ) | ( n3034 & ~n3036 ) | ( n3035 & ~n3036 ) ;
  assign n3038 = ( n2899 & ~n2909 ) | ( n2899 & n2912 ) | ( ~n2909 & n2912 ) ;
  assign n3039 = ( n2899 & n2909 ) | ( n2899 & n2912 ) | ( n2909 & n2912 ) ;
  assign n3040 = ( n2909 & n3038 ) | ( n2909 & ~n3039 ) | ( n3038 & ~n3039 ) ;
  assign n3041 = ( n2938 & n2944 ) | ( n2938 & ~n2977 ) | ( n2944 & ~n2977 ) ;
  assign n3042 = ( n2938 & n2944 ) | ( n2938 & n2977 ) | ( n2944 & n2977 ) ;
  assign n3043 = ( n2977 & n3041 ) | ( n2977 & ~n3042 ) | ( n3041 & ~n3042 ) ;
  assign n3044 = ( ~n2959 & n2965 ) | ( ~n2959 & n2989 ) | ( n2965 & n2989 ) ;
  assign n3045 = ( n2959 & n2965 ) | ( n2959 & n2989 ) | ( n2965 & n2989 ) ;
  assign n3046 = ( n2959 & n3044 ) | ( n2959 & ~n3045 ) | ( n3044 & ~n3045 ) ;
  assign n3047 = ( n2968 & n3043 ) | ( n2968 & n3046 ) | ( n3043 & n3046 ) ;
  assign n3048 = ( n2968 & ~n3043 ) | ( n2968 & n3046 ) | ( ~n3043 & n3046 ) ;
  assign n3049 = ( n3043 & ~n3047 ) | ( n3043 & n3048 ) | ( ~n3047 & n3048 ) ;
  assign n3050 = ( ~n2970 & n3040 ) | ( ~n2970 & n3049 ) | ( n3040 & n3049 ) ;
  assign n3051 = ( n2970 & n3040 ) | ( n2970 & n3049 ) | ( n3040 & n3049 ) ;
  assign n3052 = ( n2970 & n3050 ) | ( n2970 & ~n3051 ) | ( n3050 & ~n3051 ) ;
  assign n3053 = ( ~n2932 & n2953 ) | ( ~n2932 & n2983 ) | ( n2953 & n2983 ) ;
  assign n3054 = ( n2932 & n2953 ) | ( n2932 & n2983 ) | ( n2953 & n2983 ) ;
  assign n3055 = ( n2932 & n3053 ) | ( n2932 & ~n3054 ) | ( n3053 & ~n3054 ) ;
  assign n3056 = ( n2947 & n2992 ) | ( n2947 & n3055 ) | ( n2992 & n3055 ) ;
  assign n3057 = ( n2947 & n2992 ) | ( n2947 & ~n3055 ) | ( n2992 & ~n3055 ) ;
  assign n3058 = ( n3055 & ~n3056 ) | ( n3055 & n3057 ) | ( ~n3056 & n3057 ) ;
  assign n3059 = x15 & x39 ;
  assign n3060 = x7 & x47 ;
  assign n3061 = x8 & x46 ;
  assign n3062 = ( ~n3059 & n3060 ) | ( ~n3059 & n3061 ) | ( n3060 & n3061 ) ;
  assign n3063 = ( n3059 & n3060 ) | ( n3059 & n3061 ) | ( n3060 & n3061 ) ;
  assign n3064 = ( n3059 & n3062 ) | ( n3059 & ~n3063 ) | ( n3062 & ~n3063 ) ;
  assign n3065 = x3 & x51 ;
  assign n3066 = x4 & x50 ;
  assign n3067 = x2 & x52 ;
  assign n3068 = ( ~n3065 & n3066 ) | ( ~n3065 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3069 = ( n3065 & n3066 ) | ( n3065 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3070 = ( n3065 & n3068 ) | ( n3065 & ~n3069 ) | ( n3068 & ~n3069 ) ;
  assign n3071 = x10 & x44 ;
  assign n3072 = x14 & x40 ;
  assign n3073 = x9 & x45 ;
  assign n3074 = ( ~n3071 & n3072 ) | ( ~n3071 & n3073 ) | ( n3072 & n3073 ) ;
  assign n3075 = ( n3071 & n3072 ) | ( n3071 & n3073 ) | ( n3072 & n3073 ) ;
  assign n3076 = ( n3071 & n3074 ) | ( n3071 & ~n3075 ) | ( n3074 & ~n3075 ) ;
  assign n3077 = ( ~n3064 & n3070 ) | ( ~n3064 & n3076 ) | ( n3070 & n3076 ) ;
  assign n3078 = ( n3064 & n3070 ) | ( n3064 & n3076 ) | ( n3070 & n3076 ) ;
  assign n3079 = ( n3064 & n3077 ) | ( n3064 & ~n3078 ) | ( n3077 & ~n3078 ) ;
  assign n3080 = x11 & x43 ;
  assign n3081 = x13 & x41 ;
  assign n3082 = x12 & x42 ;
  assign n3083 = ( ~n3080 & n3081 ) | ( ~n3080 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = ( n3080 & n3081 ) | ( n3080 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3085 = ( n3080 & n3083 ) | ( n3080 & ~n3084 ) | ( n3083 & ~n3084 ) ;
  assign n3086 = x16 & x38 ;
  assign n3087 = x6 & x48 ;
  assign n3088 = x17 & x37 ;
  assign n3089 = ( ~n3086 & n3087 ) | ( ~n3086 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3090 = ( n3086 & n3087 ) | ( n3086 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3091 = ( n3086 & n3089 ) | ( n3086 & ~n3090 ) | ( n3089 & ~n3090 ) ;
  assign n3092 = x18 & x36 ;
  assign n3093 = x5 & x49 ;
  assign n3094 = x20 & x34 ;
  assign n3095 = ( ~n3092 & n3093 ) | ( ~n3092 & n3094 ) | ( n3093 & n3094 ) ;
  assign n3096 = ( n3092 & n3093 ) | ( n3092 & n3094 ) | ( n3093 & n3094 ) ;
  assign n3097 = ( n3092 & n3095 ) | ( n3092 & ~n3096 ) | ( n3095 & ~n3096 ) ;
  assign n3098 = ( ~n3085 & n3091 ) | ( ~n3085 & n3097 ) | ( n3091 & n3097 ) ;
  assign n3099 = ( n3085 & n3091 ) | ( n3085 & n3097 ) | ( n3091 & n3097 ) ;
  assign n3100 = ( n3085 & n3098 ) | ( n3085 & ~n3099 ) | ( n3098 & ~n3099 ) ;
  assign n3101 = ( n2921 & n3079 ) | ( n2921 & n3100 ) | ( n3079 & n3100 ) ;
  assign n3102 = ( ~n2921 & n3079 ) | ( ~n2921 & n3100 ) | ( n3079 & n3100 ) ;
  assign n3103 = ( n2921 & ~n3101 ) | ( n2921 & n3102 ) | ( ~n3101 & n3102 ) ;
  assign n3104 = ( n2994 & n3058 ) | ( n2994 & n3103 ) | ( n3058 & n3103 ) ;
  assign n3105 = ( n2994 & ~n3058 ) | ( n2994 & n3103 ) | ( ~n3058 & n3103 ) ;
  assign n3106 = ( n3058 & ~n3104 ) | ( n3058 & n3105 ) | ( ~n3104 & n3105 ) ;
  assign n3107 = ( n2997 & n3052 ) | ( n2997 & n3106 ) | ( n3052 & n3106 ) ;
  assign n3108 = ( ~n2997 & n3052 ) | ( ~n2997 & n3106 ) | ( n3052 & n3106 ) ;
  assign n3109 = ( n2997 & ~n3107 ) | ( n2997 & n3108 ) | ( ~n3107 & n3108 ) ;
  assign n3110 = ( n2926 & n3037 ) | ( n2926 & n3109 ) | ( n3037 & n3109 ) ;
  assign n3111 = ( ~n2926 & n3037 ) | ( ~n2926 & n3109 ) | ( n3037 & n3109 ) ;
  assign n3112 = ( n2926 & ~n3110 ) | ( n2926 & n3111 ) | ( ~n3110 & n3111 ) ;
  assign n3113 = ( n3000 & n3004 ) | ( n3000 & n3112 ) | ( n3004 & n3112 ) ;
  assign n3114 = ( n3000 & ~n3004 ) | ( n3000 & n3112 ) | ( ~n3004 & n3112 ) ;
  assign n3115 = ( n3004 & ~n3113 ) | ( n3004 & n3114 ) | ( ~n3113 & n3114 ) ;
  assign n3116 = x6 & x49 ;
  assign n3117 = x17 & x38 ;
  assign n3118 = x3 & x52 ;
  assign n3119 = ( ~n3116 & n3117 ) | ( ~n3116 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3120 = ( n3116 & n3117 ) | ( n3116 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3121 = ( n3116 & n3119 ) | ( n3116 & ~n3120 ) | ( n3119 & ~n3120 ) ;
  assign n3122 = x9 & x46 ;
  assign n3123 = x14 & x41 ;
  assign n3124 = x15 & x40 ;
  assign n3125 = ( ~n3122 & n3123 ) | ( ~n3122 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3126 = ( n3122 & n3123 ) | ( n3122 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3127 = ( n3122 & n3125 ) | ( n3122 & ~n3126 ) | ( n3125 & ~n3126 ) ;
  assign n3128 = ( ~n3042 & n3121 ) | ( ~n3042 & n3127 ) | ( n3121 & n3127 ) ;
  assign n3129 = ( n3042 & n3121 ) | ( n3042 & n3127 ) | ( n3121 & n3127 ) ;
  assign n3130 = ( n3042 & n3128 ) | ( n3042 & ~n3129 ) | ( n3128 & ~n3129 ) ;
  assign n3131 = ( n3047 & n3056 ) | ( n3047 & n3130 ) | ( n3056 & n3130 ) ;
  assign n3132 = ( n3047 & ~n3056 ) | ( n3047 & n3130 ) | ( ~n3056 & n3130 ) ;
  assign n3133 = ( n3056 & ~n3131 ) | ( n3056 & n3132 ) | ( ~n3131 & n3132 ) ;
  assign n3134 = ( n3051 & n3104 ) | ( n3051 & n3133 ) | ( n3104 & n3133 ) ;
  assign n3135 = ( n3051 & ~n3104 ) | ( n3051 & n3133 ) | ( ~n3104 & n3133 ) ;
  assign n3136 = ( n3104 & ~n3134 ) | ( n3104 & n3135 ) | ( ~n3134 & n3135 ) ;
  assign n3137 = x13 & x42 ;
  assign n3138 = x10 & x45 ;
  assign n3139 = x11 & x44 ;
  assign n3140 = ( ~n3137 & n3138 ) | ( ~n3137 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3141 = ( n3137 & n3138 ) | ( n3137 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3142 = ( n3137 & n3140 ) | ( n3137 & ~n3141 ) | ( n3140 & ~n3141 ) ;
  assign n3143 = x27 & x28 ;
  assign n3144 = x26 & x29 ;
  assign n3145 = x12 & x43 ;
  assign n3146 = ( ~n3143 & n3144 ) | ( ~n3143 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3147 = ( n3143 & n3144 ) | ( n3143 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3148 = ( n3143 & n3146 ) | ( n3143 & ~n3147 ) | ( n3146 & ~n3147 ) ;
  assign n3149 = x8 & x47 ;
  assign n3150 = x16 & x39 ;
  assign n3151 = x7 & x48 ;
  assign n3152 = ( ~n3149 & n3150 ) | ( ~n3149 & n3151 ) | ( n3150 & n3151 ) ;
  assign n3153 = ( n3149 & n3150 ) | ( n3149 & n3151 ) | ( n3150 & n3151 ) ;
  assign n3154 = ( n3149 & n3152 ) | ( n3149 & ~n3153 ) | ( n3152 & ~n3153 ) ;
  assign n3155 = ( ~n3142 & n3148 ) | ( ~n3142 & n3154 ) | ( n3148 & n3154 ) ;
  assign n3156 = ( n3142 & n3148 ) | ( n3142 & n3154 ) | ( n3148 & n3154 ) ;
  assign n3157 = ( n3142 & n3155 ) | ( n3142 & ~n3156 ) | ( n3155 & ~n3156 ) ;
  assign n3158 = x20 & x35 ;
  assign n3159 = x22 & x33 ;
  assign n3160 = x21 & x34 ;
  assign n3161 = ( ~n3158 & n3159 ) | ( ~n3158 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3162 = ( n3158 & n3159 ) | ( n3158 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3163 = ( n3158 & n3161 ) | ( n3158 & ~n3162 ) | ( n3161 & ~n3162 ) ;
  assign n3164 = x2 & x53 ;
  assign n3165 = x0 & x55 ;
  assign n3166 = x4 & x51 ;
  assign n3167 = ( ~n3164 & n3165 ) | ( ~n3164 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3168 = ( n3164 & n3165 ) | ( n3164 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3169 = ( n3164 & n3167 ) | ( n3164 & ~n3168 ) | ( n3167 & ~n3168 ) ;
  assign n3170 = x24 & x31 ;
  assign n3171 = x25 & x30 ;
  assign n3172 = x23 & x32 ;
  assign n3173 = ( ~n3170 & n3171 ) | ( ~n3170 & n3172 ) | ( n3171 & n3172 ) ;
  assign n3174 = ( n3170 & n3171 ) | ( n3170 & n3172 ) | ( n3171 & n3172 ) ;
  assign n3175 = ( n3170 & n3173 ) | ( n3170 & ~n3174 ) | ( n3173 & ~n3174 ) ;
  assign n3176 = ( ~n3163 & n3169 ) | ( ~n3163 & n3175 ) | ( n3169 & n3175 ) ;
  assign n3177 = ( n3163 & n3169 ) | ( n3163 & n3175 ) | ( n3169 & n3175 ) ;
  assign n3178 = ( n3163 & n3176 ) | ( n3163 & ~n3177 ) | ( n3176 & ~n3177 ) ;
  assign n3179 = ( n3039 & n3157 ) | ( n3039 & n3178 ) | ( n3157 & n3178 ) ;
  assign n3180 = ( ~n3039 & n3157 ) | ( ~n3039 & n3178 ) | ( n3157 & n3178 ) ;
  assign n3181 = ( n3039 & ~n3179 ) | ( n3039 & n3180 ) | ( ~n3179 & n3180 ) ;
  assign n3182 = ( ~n3021 & n3027 ) | ( ~n3021 & n3090 ) | ( n3027 & n3090 ) ;
  assign n3183 = ( n3021 & n3027 ) | ( n3021 & n3090 ) | ( n3027 & n3090 ) ;
  assign n3184 = ( n3021 & n3182 ) | ( n3021 & ~n3183 ) | ( n3182 & ~n3183 ) ;
  assign n3185 = ( n3078 & n3099 ) | ( n3078 & n3184 ) | ( n3099 & n3184 ) ;
  assign n3186 = ( n3078 & n3099 ) | ( n3078 & ~n3184 ) | ( n3099 & ~n3184 ) ;
  assign n3187 = ( n3184 & ~n3185 ) | ( n3184 & n3186 ) | ( ~n3185 & n3186 ) ;
  assign n3188 = ( n3033 & n3181 ) | ( n3033 & n3187 ) | ( n3181 & n3187 ) ;
  assign n3189 = ( ~n3033 & n3181 ) | ( ~n3033 & n3187 ) | ( n3181 & n3187 ) ;
  assign n3190 = ( n3033 & ~n3188 ) | ( n3033 & n3189 ) | ( ~n3188 & n3189 ) ;
  assign n3191 = ( x28 & ~n3007 ) | ( x28 & n3011 ) | ( ~n3007 & n3011 ) ;
  assign n3192 = x1 & x54 ;
  assign n3193 = ( n3084 & n3191 ) | ( n3084 & ~n3192 ) | ( n3191 & ~n3192 ) ;
  assign n3194 = ( ~n3084 & n3191 ) | ( ~n3084 & n3192 ) | ( n3191 & n3192 ) ;
  assign n3195 = ( ~n3191 & n3193 ) | ( ~n3191 & n3194 ) | ( n3193 & n3194 ) ;
  assign n3196 = ( n3045 & n3054 ) | ( n3045 & ~n3195 ) | ( n3054 & ~n3195 ) ;
  assign n3197 = ( n3045 & n3054 ) | ( n3045 & n3195 ) | ( n3054 & n3195 ) ;
  assign n3198 = ( n3195 & n3196 ) | ( n3195 & ~n3197 ) | ( n3196 & ~n3197 ) ;
  assign n3199 = x19 & x36 ;
  assign n3200 = x5 & x50 ;
  assign n3201 = ( ~n1580 & n3199 ) | ( ~n1580 & n3200 ) | ( n3199 & n3200 ) ;
  assign n3202 = ( n1580 & n3199 ) | ( n1580 & n3200 ) | ( n3199 & n3200 ) ;
  assign n3203 = ( n1580 & n3201 ) | ( n1580 & ~n3202 ) | ( n3201 & ~n3202 ) ;
  assign n3204 = ( ~n3014 & n3063 ) | ( ~n3014 & n3203 ) | ( n3063 & n3203 ) ;
  assign n3205 = ( n3014 & n3063 ) | ( n3014 & n3203 ) | ( n3063 & n3203 ) ;
  assign n3206 = ( n3014 & n3204 ) | ( n3014 & ~n3205 ) | ( n3204 & ~n3205 ) ;
  assign n3207 = ( n3069 & ~n3075 ) | ( n3069 & n3096 ) | ( ~n3075 & n3096 ) ;
  assign n3208 = ( n3069 & n3075 ) | ( n3069 & n3096 ) | ( n3075 & n3096 ) ;
  assign n3209 = ( n3075 & n3207 ) | ( n3075 & ~n3208 ) | ( n3207 & ~n3208 ) ;
  assign n3210 = ( n3029 & ~n3206 ) | ( n3029 & n3209 ) | ( ~n3206 & n3209 ) ;
  assign n3211 = ( n3029 & n3206 ) | ( n3029 & n3209 ) | ( n3206 & n3209 ) ;
  assign n3212 = ( n3206 & n3210 ) | ( n3206 & ~n3211 ) | ( n3210 & ~n3211 ) ;
  assign n3213 = ( n3101 & ~n3198 ) | ( n3101 & n3212 ) | ( ~n3198 & n3212 ) ;
  assign n3214 = ( n3101 & n3198 ) | ( n3101 & n3212 ) | ( n3198 & n3212 ) ;
  assign n3215 = ( n3198 & n3213 ) | ( n3198 & ~n3214 ) | ( n3213 & ~n3214 ) ;
  assign n3216 = ( n3036 & ~n3190 ) | ( n3036 & n3215 ) | ( ~n3190 & n3215 ) ;
  assign n3217 = ( n3036 & n3190 ) | ( n3036 & n3215 ) | ( n3190 & n3215 ) ;
  assign n3218 = ( n3190 & n3216 ) | ( n3190 & ~n3217 ) | ( n3216 & ~n3217 ) ;
  assign n3219 = ( n3107 & ~n3136 ) | ( n3107 & n3218 ) | ( ~n3136 & n3218 ) ;
  assign n3220 = ( n3107 & n3136 ) | ( n3107 & n3218 ) | ( n3136 & n3218 ) ;
  assign n3221 = ( n3136 & n3219 ) | ( n3136 & ~n3220 ) | ( n3219 & ~n3220 ) ;
  assign n3222 = ( n3110 & ~n3113 ) | ( n3110 & n3221 ) | ( ~n3113 & n3221 ) ;
  assign n3223 = ( n3110 & n3113 ) | ( n3110 & n3221 ) | ( n3113 & n3221 ) ;
  assign n3224 = ( n3113 & n3222 ) | ( n3113 & ~n3223 ) | ( n3222 & ~n3223 ) ;
  assign n3225 = ( x2 & ~x54 ) | ( x2 & n933 ) | ( ~x54 & n933 ) ;
  assign n3226 = x0 & x56 ;
  assign n3227 = x2 | n933 ;
  assign n3228 = ( ~n3225 & n3226 ) | ( ~n3225 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3229 = ( n3225 & n3226 ) | ( n3225 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3230 = ( n3225 & n3228 ) | ( n3225 & ~n3229 ) | ( n3228 & ~n3229 ) ;
  assign n3231 = x4 & x52 ;
  assign n3232 = x19 & x37 ;
  assign n3233 = x3 & x53 ;
  assign n3234 = ( ~n3231 & n3232 ) | ( ~n3231 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3235 = ( n3231 & n3232 ) | ( n3231 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3236 = ( n3231 & n3234 ) | ( n3231 & ~n3235 ) | ( n3234 & ~n3235 ) ;
  assign n3237 = ( n3153 & ~n3230 ) | ( n3153 & n3236 ) | ( ~n3230 & n3236 ) ;
  assign n3238 = ( n3153 & n3230 ) | ( n3153 & n3236 ) | ( n3230 & n3236 ) ;
  assign n3239 = ( n3230 & n3237 ) | ( n3230 & ~n3238 ) | ( n3237 & ~n3238 ) ;
  assign n3240 = x11 & x45 ;
  assign n3241 = x13 & x43 ;
  assign n3242 = x12 & x44 ;
  assign n3243 = ( ~n3240 & n3241 ) | ( ~n3240 & n3242 ) | ( n3241 & n3242 ) ;
  assign n3244 = ( n3240 & n3241 ) | ( n3240 & n3242 ) | ( n3241 & n3242 ) ;
  assign n3245 = ( n3240 & n3243 ) | ( n3240 & ~n3244 ) | ( n3243 & ~n3244 ) ;
  assign n3246 = x6 & x50 ;
  assign n3247 = x7 & x49 ;
  assign n3248 = x17 & x39 ;
  assign n3249 = ( ~n3246 & n3247 ) | ( ~n3246 & n3248 ) | ( n3247 & n3248 ) ;
  assign n3250 = ( n3246 & n3247 ) | ( n3246 & n3248 ) | ( n3247 & n3248 ) ;
  assign n3251 = ( n3246 & n3249 ) | ( n3246 & ~n3250 ) | ( n3249 & ~n3250 ) ;
  assign n3252 = x15 & x41 ;
  assign n3253 = x8 & x48 ;
  assign n3254 = x16 & x40 ;
  assign n3255 = ( ~n3252 & n3253 ) | ( ~n3252 & n3254 ) | ( n3253 & n3254 ) ;
  assign n3256 = ( n3252 & n3253 ) | ( n3252 & n3254 ) | ( n3253 & n3254 ) ;
  assign n3257 = ( n3252 & n3255 ) | ( n3252 & ~n3256 ) | ( n3255 & ~n3256 ) ;
  assign n3258 = ( ~n3245 & n3251 ) | ( ~n3245 & n3257 ) | ( n3251 & n3257 ) ;
  assign n3259 = ( n3245 & n3251 ) | ( n3245 & n3257 ) | ( n3251 & n3257 ) ;
  assign n3260 = ( n3245 & n3258 ) | ( n3245 & ~n3259 ) | ( n3258 & ~n3259 ) ;
  assign n3261 = x20 & x36 ;
  assign n3262 = x22 & x34 ;
  assign n3263 = x23 & x33 ;
  assign n3264 = ( ~n3261 & n3262 ) | ( ~n3261 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3265 = ( n3261 & n3262 ) | ( n3261 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3266 = ( n3261 & n3264 ) | ( n3261 & ~n3265 ) | ( n3264 & ~n3265 ) ;
  assign n3267 = x14 & x42 ;
  assign n3268 = x10 & x46 ;
  assign n3269 = x9 & x47 ;
  assign n3270 = ( ~n3267 & n3268 ) | ( ~n3267 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3271 = ( n3267 & n3268 ) | ( n3267 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3272 = ( n3267 & n3270 ) | ( n3267 & ~n3271 ) | ( n3270 & ~n3271 ) ;
  assign n3273 = x25 & x31 ;
  assign n3274 = x24 & x32 ;
  assign n3275 = x26 & x30 ;
  assign n3276 = ( ~n3273 & n3274 ) | ( ~n3273 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3277 = ( n3273 & n3274 ) | ( n3273 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3278 = ( n3273 & n3276 ) | ( n3273 & ~n3277 ) | ( n3276 & ~n3277 ) ;
  assign n3279 = ( ~n3266 & n3272 ) | ( ~n3266 & n3278 ) | ( n3272 & n3278 ) ;
  assign n3280 = ( n3266 & n3272 ) | ( n3266 & n3278 ) | ( n3272 & n3278 ) ;
  assign n3281 = ( n3266 & n3279 ) | ( n3266 & ~n3280 ) | ( n3279 & ~n3280 ) ;
  assign n3282 = ( n3239 & n3260 ) | ( n3239 & n3281 ) | ( n3260 & n3281 ) ;
  assign n3283 = ( ~n3239 & n3260 ) | ( ~n3239 & n3281 ) | ( n3260 & n3281 ) ;
  assign n3284 = ( n3239 & ~n3282 ) | ( n3239 & n3283 ) | ( ~n3282 & n3283 ) ;
  assign n3285 = ( ~n3120 & n3162 ) | ( ~n3120 & n3174 ) | ( n3162 & n3174 ) ;
  assign n3286 = ( n3120 & n3162 ) | ( n3120 & n3174 ) | ( n3162 & n3174 ) ;
  assign n3287 = ( n3120 & n3285 ) | ( n3120 & ~n3286 ) | ( n3285 & ~n3286 ) ;
  assign n3288 = x27 & x29 ;
  assign n3289 = x1 & x55 ;
  assign n3290 = n3288 | n3289 ;
  assign n3291 = x29 & x55 ;
  assign n3292 = n892 & n3291 ;
  assign n3293 = n3290 & ~n3292 ;
  assign n3294 = ( ~n3141 & n3147 ) | ( ~n3141 & n3293 ) | ( n3147 & n3293 ) ;
  assign n3295 = ( n3141 & n3147 ) | ( n3141 & n3293 ) | ( n3147 & n3293 ) ;
  assign n3296 = ( n3141 & n3294 ) | ( n3141 & ~n3295 ) | ( n3294 & ~n3295 ) ;
  assign n3297 = ( n3156 & n3287 ) | ( n3156 & n3296 ) | ( n3287 & n3296 ) ;
  assign n3298 = ( ~n3156 & n3287 ) | ( ~n3156 & n3296 ) | ( n3287 & n3296 ) ;
  assign n3299 = ( n3156 & ~n3297 ) | ( n3156 & n3298 ) | ( ~n3297 & n3298 ) ;
  assign n3300 = ( n3131 & n3284 ) | ( n3131 & n3299 ) | ( n3284 & n3299 ) ;
  assign n3301 = ( ~n3131 & n3284 ) | ( ~n3131 & n3299 ) | ( n3284 & n3299 ) ;
  assign n3302 = ( n3131 & ~n3300 ) | ( n3131 & n3301 ) | ( ~n3300 & n3301 ) ;
  assign n3303 = ( n3177 & n3183 ) | ( n3177 & ~n3205 ) | ( n3183 & ~n3205 ) ;
  assign n3304 = ( n3177 & n3183 ) | ( n3177 & n3205 ) | ( n3183 & n3205 ) ;
  assign n3305 = ( n3205 & n3303 ) | ( n3205 & ~n3304 ) | ( n3303 & ~n3304 ) ;
  assign n3306 = ( ~n3126 & n3168 ) | ( ~n3126 & n3202 ) | ( n3168 & n3202 ) ;
  assign n3307 = ( n3126 & n3168 ) | ( n3126 & n3202 ) | ( n3168 & n3202 ) ;
  assign n3308 = ( n3126 & n3306 ) | ( n3126 & ~n3307 ) | ( n3306 & ~n3307 ) ;
  assign n3309 = ( n3129 & n3197 ) | ( n3129 & ~n3308 ) | ( n3197 & ~n3308 ) ;
  assign n3310 = ( n3129 & n3197 ) | ( n3129 & n3308 ) | ( n3197 & n3308 ) ;
  assign n3311 = ( n3308 & n3309 ) | ( n3308 & ~n3310 ) | ( n3309 & ~n3310 ) ;
  assign n3312 = ( n3179 & ~n3305 ) | ( n3179 & n3311 ) | ( ~n3305 & n3311 ) ;
  assign n3313 = ( n3179 & n3305 ) | ( n3179 & n3311 ) | ( n3305 & n3311 ) ;
  assign n3314 = ( n3305 & n3312 ) | ( n3305 & ~n3313 ) | ( n3312 & ~n3313 ) ;
  assign n3315 = ( n3134 & ~n3302 ) | ( n3134 & n3314 ) | ( ~n3302 & n3314 ) ;
  assign n3316 = ( n3134 & n3302 ) | ( n3134 & n3314 ) | ( n3302 & n3314 ) ;
  assign n3317 = ( n3302 & n3315 ) | ( n3302 & ~n3316 ) | ( n3315 & ~n3316 ) ;
  assign n3318 = ( n3010 & n3084 ) | ( n3010 & ~n3195 ) | ( n3084 & ~n3195 ) ;
  assign n3319 = x18 & x38 ;
  assign n3320 = x21 & x35 ;
  assign n3321 = x5 & x51 ;
  assign n3322 = ( ~n3319 & n3320 ) | ( ~n3319 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = ( n3319 & n3320 ) | ( n3319 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3324 = ( n3319 & n3322 ) | ( n3319 & ~n3323 ) | ( n3322 & ~n3323 ) ;
  assign n3325 = ( n3208 & ~n3318 ) | ( n3208 & n3324 ) | ( ~n3318 & n3324 ) ;
  assign n3326 = ( n3208 & n3318 ) | ( n3208 & n3324 ) | ( n3318 & n3324 ) ;
  assign n3327 = ( n3318 & n3325 ) | ( n3318 & ~n3326 ) | ( n3325 & ~n3326 ) ;
  assign n3328 = ( n3185 & n3211 ) | ( n3185 & n3327 ) | ( n3211 & n3327 ) ;
  assign n3329 = ( n3185 & n3211 ) | ( n3185 & ~n3327 ) | ( n3211 & ~n3327 ) ;
  assign n3330 = ( n3327 & ~n3328 ) | ( n3327 & n3329 ) | ( ~n3328 & n3329 ) ;
  assign n3331 = ( n3188 & n3214 ) | ( n3188 & n3330 ) | ( n3214 & n3330 ) ;
  assign n3332 = ( ~n3188 & n3214 ) | ( ~n3188 & n3330 ) | ( n3214 & n3330 ) ;
  assign n3333 = ( n3188 & ~n3331 ) | ( n3188 & n3332 ) | ( ~n3331 & n3332 ) ;
  assign n3334 = ( n3217 & n3317 ) | ( n3217 & n3333 ) | ( n3317 & n3333 ) ;
  assign n3335 = ( ~n3217 & n3317 ) | ( ~n3217 & n3333 ) | ( n3317 & n3333 ) ;
  assign n3336 = ( n3217 & ~n3334 ) | ( n3217 & n3335 ) | ( ~n3334 & n3335 ) ;
  assign n3337 = ( n3220 & n3223 ) | ( n3220 & n3336 ) | ( n3223 & n3336 ) ;
  assign n3338 = ( n3220 & ~n3223 ) | ( n3220 & n3336 ) | ( ~n3223 & n3336 ) ;
  assign n3339 = ( n3223 & ~n3337 ) | ( n3223 & n3338 ) | ( ~n3337 & n3338 ) ;
  assign n3340 = x1 & x56 ;
  assign n3341 = x29 & x56 ;
  assign n3342 = ( n3292 & n3340 ) | ( n3292 & ~n3341 ) | ( n3340 & ~n3341 ) ;
  assign n3343 = x29 & ~n3340 ;
  assign n3344 = x0 & x57 ;
  assign n3345 = ( n3342 & n3343 ) | ( n3342 & n3344 ) | ( n3343 & n3344 ) ;
  assign n3346 = ( ~n3342 & n3343 ) | ( ~n3342 & n3344 ) | ( n3343 & n3344 ) ;
  assign n3347 = ( n3342 & ~n3345 ) | ( n3342 & n3346 ) | ( ~n3345 & n3346 ) ;
  assign n3348 = ( n3286 & n3307 ) | ( n3286 & n3347 ) | ( n3307 & n3347 ) ;
  assign n3349 = ( n3286 & n3307 ) | ( n3286 & ~n3347 ) | ( n3307 & ~n3347 ) ;
  assign n3350 = ( n3347 & ~n3348 ) | ( n3347 & n3349 ) | ( ~n3348 & n3349 ) ;
  assign n3351 = ( n3297 & ~n3310 ) | ( n3297 & n3350 ) | ( ~n3310 & n3350 ) ;
  assign n3352 = ( n3297 & n3310 ) | ( n3297 & n3350 ) | ( n3310 & n3350 ) ;
  assign n3353 = ( n3310 & n3351 ) | ( n3310 & ~n3352 ) | ( n3351 & ~n3352 ) ;
  assign n3354 = ( n3300 & n3313 ) | ( n3300 & ~n3353 ) | ( n3313 & ~n3353 ) ;
  assign n3355 = ( n3300 & n3313 ) | ( n3300 & n3353 ) | ( n3313 & n3353 ) ;
  assign n3356 = ( n3353 & n3354 ) | ( n3353 & ~n3355 ) | ( n3354 & ~n3355 ) ;
  assign n3357 = ( ~n3238 & n3280 ) | ( ~n3238 & n3295 ) | ( n3280 & n3295 ) ;
  assign n3358 = ( n3238 & n3280 ) | ( n3238 & n3295 ) | ( n3280 & n3295 ) ;
  assign n3359 = ( n3238 & n3357 ) | ( n3238 & ~n3358 ) | ( n3357 & ~n3358 ) ;
  assign n3360 = ( x2 & n933 ) | ( x2 & n3226 ) | ( n933 & n3226 ) ;
  assign n3361 = x54 & n3360 ;
  assign n3362 = ( n3235 & n3265 ) | ( n3235 & n3361 ) | ( n3265 & n3361 ) ;
  assign n3363 = ( n3235 & n3265 ) | ( n3235 & ~n3361 ) | ( n3265 & ~n3361 ) ;
  assign n3364 = ( n3361 & ~n3362 ) | ( n3361 & n3363 ) | ( ~n3362 & n3363 ) ;
  assign n3365 = ( n3250 & n3256 ) | ( n3250 & ~n3277 ) | ( n3256 & ~n3277 ) ;
  assign n3366 = ( n3250 & n3256 ) | ( n3250 & n3277 ) | ( n3256 & n3277 ) ;
  assign n3367 = ( n3277 & n3365 ) | ( n3277 & ~n3366 ) | ( n3365 & ~n3366 ) ;
  assign n3368 = ( n3259 & n3364 ) | ( n3259 & n3367 ) | ( n3364 & n3367 ) ;
  assign n3369 = ( n3259 & ~n3364 ) | ( n3259 & n3367 ) | ( ~n3364 & n3367 ) ;
  assign n3370 = ( n3364 & ~n3368 ) | ( n3364 & n3369 ) | ( ~n3368 & n3369 ) ;
  assign n3371 = ( n3282 & n3359 ) | ( n3282 & n3370 ) | ( n3359 & n3370 ) ;
  assign n3372 = ( ~n3282 & n3359 ) | ( ~n3282 & n3370 ) | ( n3359 & n3370 ) ;
  assign n3373 = ( n3282 & ~n3371 ) | ( n3282 & n3372 ) | ( ~n3371 & n3372 ) ;
  assign n3374 = ( n3244 & n3271 ) | ( n3244 & ~n3323 ) | ( n3271 & ~n3323 ) ;
  assign n3375 = ( n3244 & n3271 ) | ( n3244 & n3323 ) | ( n3271 & n3323 ) ;
  assign n3376 = ( n3323 & n3374 ) | ( n3323 & ~n3375 ) | ( n3374 & ~n3375 ) ;
  assign n3377 = x22 & x35 ;
  assign n3378 = x23 & x34 ;
  assign n3379 = x21 & x36 ;
  assign n3380 = ( ~n3377 & n3378 ) | ( ~n3377 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = ( n3377 & n3378 ) | ( n3377 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3382 = ( n3377 & n3380 ) | ( n3377 & ~n3381 ) | ( n3380 & ~n3381 ) ;
  assign n3383 = x7 & x50 ;
  assign n3384 = x16 & x41 ;
  assign n3385 = x8 & x49 ;
  assign n3386 = ( ~n3383 & n3384 ) | ( ~n3383 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3387 = ( n3383 & n3384 ) | ( n3383 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3388 = ( n3383 & n3386 ) | ( n3383 & ~n3387 ) | ( n3386 & ~n3387 ) ;
  assign n3389 = x26 & x31 ;
  assign n3390 = x24 & x33 ;
  assign n3391 = x25 & x32 ;
  assign n3392 = ( ~n3389 & n3390 ) | ( ~n3389 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = ( n3389 & n3390 ) | ( n3389 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3394 = ( n3389 & n3392 ) | ( n3389 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = ( ~n3382 & n3388 ) | ( ~n3382 & n3394 ) | ( n3388 & n3394 ) ;
  assign n3396 = ( n3382 & n3388 ) | ( n3382 & n3394 ) | ( n3388 & n3394 ) ;
  assign n3397 = ( n3382 & n3395 ) | ( n3382 & ~n3396 ) | ( n3395 & ~n3396 ) ;
  assign n3398 = ( n3326 & n3376 ) | ( n3326 & n3397 ) | ( n3376 & n3397 ) ;
  assign n3399 = ( ~n3326 & n3376 ) | ( ~n3326 & n3397 ) | ( n3376 & n3397 ) ;
  assign n3400 = ( n3326 & ~n3398 ) | ( n3326 & n3399 ) | ( ~n3398 & n3399 ) ;
  assign n3401 = x10 & x47 ;
  assign n3402 = x15 & x42 ;
  assign n3403 = x9 & x48 ;
  assign n3404 = ( ~n3401 & n3402 ) | ( ~n3401 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3405 = ( n3401 & n3402 ) | ( n3401 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3406 = ( n3401 & n3404 ) | ( n3401 & ~n3405 ) | ( n3404 & ~n3405 ) ;
  assign n3407 = x20 & x37 ;
  assign n3408 = x19 & x38 ;
  assign n3409 = x5 & x52 ;
  assign n3410 = ( ~n3407 & n3408 ) | ( ~n3407 & n3409 ) | ( n3408 & n3409 ) ;
  assign n3411 = ( n3407 & n3408 ) | ( n3407 & n3409 ) | ( n3408 & n3409 ) ;
  assign n3412 = ( n3407 & n3410 ) | ( n3407 & ~n3411 ) | ( n3410 & ~n3411 ) ;
  assign n3413 = x4 & x53 ;
  assign n3414 = x2 & x55 ;
  assign n3415 = x3 & x54 ;
  assign n3416 = ( ~n3413 & n3414 ) | ( ~n3413 & n3415 ) | ( n3414 & n3415 ) ;
  assign n3417 = ( n3413 & n3414 ) | ( n3413 & n3415 ) | ( n3414 & n3415 ) ;
  assign n3418 = ( n3413 & n3416 ) | ( n3413 & ~n3417 ) | ( n3416 & ~n3417 ) ;
  assign n3419 = ( ~n3406 & n3412 ) | ( ~n3406 & n3418 ) | ( n3412 & n3418 ) ;
  assign n3420 = ( n3406 & n3412 ) | ( n3406 & n3418 ) | ( n3412 & n3418 ) ;
  assign n3421 = ( n3406 & n3419 ) | ( n3406 & ~n3420 ) | ( n3419 & ~n3420 ) ;
  assign n3422 = x28 & x29 ;
  assign n3423 = x12 & x45 ;
  assign n3424 = x27 & x30 ;
  assign n3425 = ( ~n3422 & n3423 ) | ( ~n3422 & n3424 ) | ( n3423 & n3424 ) ;
  assign n3426 = ( n3422 & n3423 ) | ( n3422 & n3424 ) | ( n3423 & n3424 ) ;
  assign n3427 = ( n3422 & n3425 ) | ( n3422 & ~n3426 ) | ( n3425 & ~n3426 ) ;
  assign n3428 = x13 & x44 ;
  assign n3429 = x11 & x46 ;
  assign n3430 = x14 & x43 ;
  assign n3431 = ( ~n3428 & n3429 ) | ( ~n3428 & n3430 ) | ( n3429 & n3430 ) ;
  assign n3432 = ( n3428 & n3429 ) | ( n3428 & n3430 ) | ( n3429 & n3430 ) ;
  assign n3433 = ( n3428 & n3431 ) | ( n3428 & ~n3432 ) | ( n3431 & ~n3432 ) ;
  assign n3434 = x18 & x39 ;
  assign n3435 = x6 & x51 ;
  assign n3436 = x17 & x40 ;
  assign n3437 = ( ~n3434 & n3435 ) | ( ~n3434 & n3436 ) | ( n3435 & n3436 ) ;
  assign n3438 = ( n3434 & n3435 ) | ( n3434 & n3436 ) | ( n3435 & n3436 ) ;
  assign n3439 = ( n3434 & n3437 ) | ( n3434 & ~n3438 ) | ( n3437 & ~n3438 ) ;
  assign n3440 = ( ~n3427 & n3433 ) | ( ~n3427 & n3439 ) | ( n3433 & n3439 ) ;
  assign n3441 = ( n3427 & n3433 ) | ( n3427 & n3439 ) | ( n3433 & n3439 ) ;
  assign n3442 = ( n3427 & n3440 ) | ( n3427 & ~n3441 ) | ( n3440 & ~n3441 ) ;
  assign n3443 = ( n3304 & n3421 ) | ( n3304 & n3442 ) | ( n3421 & n3442 ) ;
  assign n3444 = ( ~n3304 & n3421 ) | ( ~n3304 & n3442 ) | ( n3421 & n3442 ) ;
  assign n3445 = ( n3304 & ~n3443 ) | ( n3304 & n3444 ) | ( ~n3443 & n3444 ) ;
  assign n3446 = ( n3328 & n3400 ) | ( n3328 & n3445 ) | ( n3400 & n3445 ) ;
  assign n3447 = ( n3328 & ~n3400 ) | ( n3328 & n3445 ) | ( ~n3400 & n3445 ) ;
  assign n3448 = ( n3400 & ~n3446 ) | ( n3400 & n3447 ) | ( ~n3446 & n3447 ) ;
  assign n3449 = ( ~n3331 & n3373 ) | ( ~n3331 & n3448 ) | ( n3373 & n3448 ) ;
  assign n3450 = ( n3331 & n3373 ) | ( n3331 & n3448 ) | ( n3373 & n3448 ) ;
  assign n3451 = ( n3331 & n3449 ) | ( n3331 & ~n3450 ) | ( n3449 & ~n3450 ) ;
  assign n3452 = ( n3316 & ~n3356 ) | ( n3316 & n3451 ) | ( ~n3356 & n3451 ) ;
  assign n3453 = ( n3316 & n3356 ) | ( n3316 & n3451 ) | ( n3356 & n3451 ) ;
  assign n3454 = ( n3356 & n3452 ) | ( n3356 & ~n3453 ) | ( n3452 & ~n3453 ) ;
  assign n3455 = ( n3334 & n3337 ) | ( n3334 & n3454 ) | ( n3337 & n3454 ) ;
  assign n3456 = ( n3334 & ~n3337 ) | ( n3334 & n3454 ) | ( ~n3337 & n3454 ) ;
  assign n3457 = ( n3337 & ~n3455 ) | ( n3337 & n3456 ) | ( ~n3455 & n3456 ) ;
  assign n3458 = ( ~n3345 & n3387 ) | ( ~n3345 & n3438 ) | ( n3387 & n3438 ) ;
  assign n3459 = ( n3345 & n3387 ) | ( n3345 & n3438 ) | ( n3387 & n3438 ) ;
  assign n3460 = ( n3345 & n3458 ) | ( n3345 & ~n3459 ) | ( n3458 & ~n3459 ) ;
  assign n3461 = x14 & x44 ;
  assign n3462 = x12 & x46 ;
  assign n3463 = x13 & x45 ;
  assign n3464 = ( ~n3461 & n3462 ) | ( ~n3461 & n3463 ) | ( n3462 & n3463 ) ;
  assign n3465 = ( n3461 & n3462 ) | ( n3461 & n3463 ) | ( n3462 & n3463 ) ;
  assign n3466 = ( n3461 & n3464 ) | ( n3461 & ~n3465 ) | ( n3464 & ~n3465 ) ;
  assign n3467 = x11 & x47 ;
  assign n3468 = x10 & x48 ;
  assign n3469 = x15 & x43 ;
  assign n3470 = ( ~n3467 & n3468 ) | ( ~n3467 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = ( n3467 & n3468 ) | ( n3467 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3472 = ( n3467 & n3470 ) | ( n3467 & ~n3471 ) | ( n3470 & ~n3471 ) ;
  assign n3473 = x3 & x55 ;
  assign n3474 = x6 & x52 ;
  assign n3475 = x19 & x39 ;
  assign n3476 = ( ~n3473 & n3474 ) | ( ~n3473 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3477 = ( n3473 & n3474 ) | ( n3473 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3478 = ( n3473 & n3476 ) | ( n3473 & ~n3477 ) | ( n3476 & ~n3477 ) ;
  assign n3479 = ( ~n3466 & n3472 ) | ( ~n3466 & n3478 ) | ( n3472 & n3478 ) ;
  assign n3480 = ( n3466 & n3472 ) | ( n3466 & n3478 ) | ( n3472 & n3478 ) ;
  assign n3481 = ( n3466 & n3479 ) | ( n3466 & ~n3480 ) | ( n3479 & ~n3480 ) ;
  assign n3482 = ( ~n3348 & n3460 ) | ( ~n3348 & n3481 ) | ( n3460 & n3481 ) ;
  assign n3483 = ( n3348 & n3460 ) | ( n3348 & n3481 ) | ( n3460 & n3481 ) ;
  assign n3484 = ( n3348 & n3482 ) | ( n3348 & ~n3483 ) | ( n3482 & ~n3483 ) ;
  assign n3485 = x25 & x33 ;
  assign n3486 = x26 & x32 ;
  assign n3487 = x27 & x31 ;
  assign n3488 = ( ~n3485 & n3486 ) | ( ~n3485 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = ( n3485 & n3486 ) | ( n3485 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3490 = ( n3485 & n3488 ) | ( n3485 & ~n3489 ) | ( n3488 & ~n3489 ) ;
  assign n3491 = x22 & x36 ;
  assign n3492 = x23 & x35 ;
  assign n3493 = x24 & x34 ;
  assign n3494 = ( ~n3491 & n3492 ) | ( ~n3491 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3495 = ( n3491 & n3492 ) | ( n3491 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3496 = ( n3491 & n3494 ) | ( n3491 & ~n3495 ) | ( n3494 & ~n3495 ) ;
  assign n3497 = x8 & x50 ;
  assign n3498 = x7 & x51 ;
  assign n3499 = x18 & x40 ;
  assign n3500 = ( ~n3497 & n3498 ) | ( ~n3497 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = ( n3497 & n3498 ) | ( n3497 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3502 = ( n3497 & n3500 ) | ( n3497 & ~n3501 ) | ( n3500 & ~n3501 ) ;
  assign n3503 = ( ~n3490 & n3496 ) | ( ~n3490 & n3502 ) | ( n3496 & n3502 ) ;
  assign n3504 = ( n3490 & n3496 ) | ( n3490 & n3502 ) | ( n3496 & n3502 ) ;
  assign n3505 = ( n3490 & n3503 ) | ( n3490 & ~n3504 ) | ( n3503 & ~n3504 ) ;
  assign n3506 = x16 & x42 ;
  assign n3507 = x17 & x41 ;
  assign n3508 = x9 & x49 ;
  assign n3509 = ( ~n3506 & n3507 ) | ( ~n3506 & n3508 ) | ( n3507 & n3508 ) ;
  assign n3510 = ( n3506 & n3507 ) | ( n3506 & n3508 ) | ( n3507 & n3508 ) ;
  assign n3511 = ( n3506 & n3509 ) | ( n3506 & ~n3510 ) | ( n3509 & ~n3510 ) ;
  assign n3512 = x4 & x54 ;
  assign n3513 = x0 & x58 ;
  assign n3514 = x2 & x56 ;
  assign n3515 = ( ~n3512 & n3513 ) | ( ~n3512 & n3514 ) | ( n3513 & n3514 ) ;
  assign n3516 = ( n3512 & n3513 ) | ( n3512 & n3514 ) | ( n3513 & n3514 ) ;
  assign n3517 = ( n3512 & n3515 ) | ( n3512 & ~n3516 ) | ( n3515 & ~n3516 ) ;
  assign n3518 = x21 & x37 ;
  assign n3519 = x5 & x53 ;
  assign n3520 = ( ~n1677 & n3518 ) | ( ~n1677 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3521 = ( n1677 & n3518 ) | ( n1677 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3522 = ( n1677 & n3520 ) | ( n1677 & ~n3521 ) | ( n3520 & ~n3521 ) ;
  assign n3523 = ( ~n3511 & n3517 ) | ( ~n3511 & n3522 ) | ( n3517 & n3522 ) ;
  assign n3524 = ( n3511 & n3517 ) | ( n3511 & n3522 ) | ( n3517 & n3522 ) ;
  assign n3525 = ( n3511 & n3523 ) | ( n3511 & ~n3524 ) | ( n3523 & ~n3524 ) ;
  assign n3526 = ( n3358 & n3505 ) | ( n3358 & n3525 ) | ( n3505 & n3525 ) ;
  assign n3527 = ( ~n3358 & n3505 ) | ( ~n3358 & n3525 ) | ( n3505 & n3525 ) ;
  assign n3528 = ( n3358 & ~n3526 ) | ( n3358 & n3527 ) | ( ~n3526 & n3527 ) ;
  assign n3529 = ( n3352 & n3484 ) | ( n3352 & n3528 ) | ( n3484 & n3528 ) ;
  assign n3530 = ( ~n3352 & n3484 ) | ( ~n3352 & n3528 ) | ( n3484 & n3528 ) ;
  assign n3531 = ( n3352 & ~n3529 ) | ( n3352 & n3530 ) | ( ~n3529 & n3530 ) ;
  assign n3532 = x28 & x30 ;
  assign n3533 = x1 & x57 ;
  assign n3534 = n3532 | n3533 ;
  assign n3535 = x30 & x57 ;
  assign n3536 = n933 & n3535 ;
  assign n3537 = n3534 & ~n3536 ;
  assign n3538 = x56 & n970 ;
  assign n3539 = ( n3426 & n3537 ) | ( n3426 & n3538 ) | ( n3537 & n3538 ) ;
  assign n3540 = ( n3426 & ~n3537 ) | ( n3426 & n3538 ) | ( ~n3537 & n3538 ) ;
  assign n3541 = ( n3537 & ~n3539 ) | ( n3537 & n3540 ) | ( ~n3539 & n3540 ) ;
  assign n3542 = ( n3420 & n3441 ) | ( n3420 & n3541 ) | ( n3441 & n3541 ) ;
  assign n3543 = ( n3420 & n3441 ) | ( n3420 & ~n3541 ) | ( n3441 & ~n3541 ) ;
  assign n3544 = ( n3541 & ~n3542 ) | ( n3541 & n3543 ) | ( ~n3542 & n3543 ) ;
  assign n3545 = ( ~n3411 & n3417 ) | ( ~n3411 & n3432 ) | ( n3417 & n3432 ) ;
  assign n3546 = ( n3411 & n3417 ) | ( n3411 & n3432 ) | ( n3417 & n3432 ) ;
  assign n3547 = ( n3411 & n3545 ) | ( n3411 & ~n3546 ) | ( n3545 & ~n3546 ) ;
  assign n3548 = ( ~n3381 & n3393 ) | ( ~n3381 & n3405 ) | ( n3393 & n3405 ) ;
  assign n3549 = ( n3381 & n3393 ) | ( n3381 & n3405 ) | ( n3393 & n3405 ) ;
  assign n3550 = ( n3381 & n3548 ) | ( n3381 & ~n3549 ) | ( n3548 & ~n3549 ) ;
  assign n3551 = ( n3396 & n3547 ) | ( n3396 & n3550 ) | ( n3547 & n3550 ) ;
  assign n3552 = ( ~n3396 & n3547 ) | ( ~n3396 & n3550 ) | ( n3547 & n3550 ) ;
  assign n3553 = ( n3396 & ~n3551 ) | ( n3396 & n3552 ) | ( ~n3551 & n3552 ) ;
  assign n3554 = ( n3443 & n3544 ) | ( n3443 & n3553 ) | ( n3544 & n3553 ) ;
  assign n3555 = ( ~n3443 & n3544 ) | ( ~n3443 & n3553 ) | ( n3544 & n3553 ) ;
  assign n3556 = ( n3443 & ~n3554 ) | ( n3443 & n3555 ) | ( ~n3554 & n3555 ) ;
  assign n3557 = ( n3355 & n3531 ) | ( n3355 & n3556 ) | ( n3531 & n3556 ) ;
  assign n3558 = ( ~n3355 & n3531 ) | ( ~n3355 & n3556 ) | ( n3531 & n3556 ) ;
  assign n3559 = ( n3355 & ~n3557 ) | ( n3355 & n3558 ) | ( ~n3557 & n3558 ) ;
  assign n3560 = ( ~n3362 & n3366 ) | ( ~n3362 & n3375 ) | ( n3366 & n3375 ) ;
  assign n3561 = ( n3362 & n3366 ) | ( n3362 & n3375 ) | ( n3366 & n3375 ) ;
  assign n3562 = ( n3362 & n3560 ) | ( n3362 & ~n3561 ) | ( n3560 & ~n3561 ) ;
  assign n3563 = ( n3368 & ~n3398 ) | ( n3368 & n3562 ) | ( ~n3398 & n3562 ) ;
  assign n3564 = ( n3368 & n3398 ) | ( n3368 & n3562 ) | ( n3398 & n3562 ) ;
  assign n3565 = ( n3398 & n3563 ) | ( n3398 & ~n3564 ) | ( n3563 & ~n3564 ) ;
  assign n3566 = ( n3371 & n3446 ) | ( n3371 & n3565 ) | ( n3446 & n3565 ) ;
  assign n3567 = ( n3371 & n3446 ) | ( n3371 & ~n3565 ) | ( n3446 & ~n3565 ) ;
  assign n3568 = ( n3565 & ~n3566 ) | ( n3565 & n3567 ) | ( ~n3566 & n3567 ) ;
  assign n3569 = ( n3450 & ~n3559 ) | ( n3450 & n3568 ) | ( ~n3559 & n3568 ) ;
  assign n3570 = ( n3450 & n3559 ) | ( n3450 & n3568 ) | ( n3559 & n3568 ) ;
  assign n3571 = ( n3559 & n3569 ) | ( n3559 & ~n3570 ) | ( n3569 & ~n3570 ) ;
  assign n3572 = ( n3453 & n3455 ) | ( n3453 & n3571 ) | ( n3455 & n3571 ) ;
  assign n3573 = ( n3453 & ~n3455 ) | ( n3453 & n3571 ) | ( ~n3455 & n3571 ) ;
  assign n3574 = ( n3455 & ~n3572 ) | ( n3455 & n3573 ) | ( ~n3572 & n3573 ) ;
  assign n3575 = x6 & x53 ;
  assign n3576 = x18 & x41 ;
  assign n3577 = x7 & x52 ;
  assign n3578 = ( ~n3575 & n3576 ) | ( ~n3575 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3579 = ( n3575 & n3576 ) | ( n3575 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3580 = ( n3575 & n3578 ) | ( n3575 & ~n3579 ) | ( n3578 & ~n3579 ) ;
  assign n3581 = x9 & x50 ;
  assign n3582 = x15 & x44 ;
  assign n3583 = x10 & x49 ;
  assign n3584 = ( ~n3581 & n3582 ) | ( ~n3581 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3585 = ( n3581 & n3582 ) | ( n3581 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3586 = ( n3581 & n3584 ) | ( n3581 & ~n3585 ) | ( n3584 & ~n3585 ) ;
  assign n3587 = ( ~n3539 & n3580 ) | ( ~n3539 & n3586 ) | ( n3580 & n3586 ) ;
  assign n3588 = ( n3539 & n3580 ) | ( n3539 & n3586 ) | ( n3580 & n3586 ) ;
  assign n3589 = ( n3539 & n3587 ) | ( n3539 & ~n3588 ) | ( n3587 & ~n3588 ) ;
  assign n3590 = x0 & x59 ;
  assign n3591 = x27 & x32 ;
  assign n3592 = x26 & x33 ;
  assign n3593 = ( ~n3590 & n3591 ) | ( ~n3590 & n3592 ) | ( n3591 & n3592 ) ;
  assign n3594 = ( n3590 & n3591 ) | ( n3590 & n3592 ) | ( n3591 & n3592 ) ;
  assign n3595 = ( n3590 & n3593 ) | ( n3590 & ~n3594 ) | ( n3593 & ~n3594 ) ;
  assign n3596 = x24 & x35 ;
  assign n3597 = x25 & x34 ;
  assign n3598 = x23 & x36 ;
  assign n3599 = ( ~n3596 & n3597 ) | ( ~n3596 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3600 = ( n3596 & n3597 ) | ( n3596 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3601 = ( n3596 & n3599 ) | ( n3596 & ~n3600 ) | ( n3599 & ~n3600 ) ;
  assign n3602 = x20 & x39 ;
  assign n3603 = x21 & x38 ;
  assign n3604 = x22 & x37 ;
  assign n3605 = ( ~n3602 & n3603 ) | ( ~n3602 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3606 = ( n3602 & n3603 ) | ( n3602 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3607 = ( n3602 & n3605 ) | ( n3602 & ~n3606 ) | ( n3605 & ~n3606 ) ;
  assign n3608 = ( ~n3595 & n3601 ) | ( ~n3595 & n3607 ) | ( n3601 & n3607 ) ;
  assign n3609 = ( n3595 & n3601 ) | ( n3595 & n3607 ) | ( n3601 & n3607 ) ;
  assign n3610 = ( n3595 & n3608 ) | ( n3595 & ~n3609 ) | ( n3608 & ~n3609 ) ;
  assign n3611 = ( n3561 & n3589 ) | ( n3561 & n3610 ) | ( n3589 & n3610 ) ;
  assign n3612 = ( n3561 & ~n3589 ) | ( n3561 & n3610 ) | ( ~n3589 & n3610 ) ;
  assign n3613 = ( n3589 & ~n3611 ) | ( n3589 & n3612 ) | ( ~n3611 & n3612 ) ;
  assign n3614 = x2 & x57 ;
  assign n3615 = x3 & x56 ;
  assign n3616 = ( ~n3536 & n3614 ) | ( ~n3536 & n3615 ) | ( n3614 & n3615 ) ;
  assign n3617 = ( n3536 & n3614 ) | ( n3536 & n3615 ) | ( n3614 & n3615 ) ;
  assign n3618 = ( n3536 & n3616 ) | ( n3536 & ~n3617 ) | ( n3616 & ~n3617 ) ;
  assign n3619 = x5 & x54 ;
  assign n3620 = x4 & x55 ;
  assign n3621 = x19 & x40 ;
  assign n3622 = ( ~n3619 & n3620 ) | ( ~n3619 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3623 = ( n3619 & n3620 ) | ( n3619 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3624 = ( n3619 & n3622 ) | ( n3619 & ~n3623 ) | ( n3622 & ~n3623 ) ;
  assign n3625 = ( n3489 & ~n3618 ) | ( n3489 & n3624 ) | ( ~n3618 & n3624 ) ;
  assign n3626 = ( n3489 & n3618 ) | ( n3489 & n3624 ) | ( n3618 & n3624 ) ;
  assign n3627 = ( n3618 & n3625 ) | ( n3618 & ~n3626 ) | ( n3625 & ~n3626 ) ;
  assign n3628 = x17 & x42 ;
  assign n3629 = x16 & x43 ;
  assign n3630 = x8 & x51 ;
  assign n3631 = ( ~n3628 & n3629 ) | ( ~n3628 & n3630 ) | ( n3629 & n3630 ) ;
  assign n3632 = ( n3628 & n3629 ) | ( n3628 & n3630 ) | ( n3629 & n3630 ) ;
  assign n3633 = ( n3628 & n3631 ) | ( n3628 & ~n3632 ) | ( n3631 & ~n3632 ) ;
  assign n3634 = x12 & x47 ;
  assign n3635 = x14 & x45 ;
  assign n3636 = x11 & x48 ;
  assign n3637 = ( ~n3634 & n3635 ) | ( ~n3634 & n3636 ) | ( n3635 & n3636 ) ;
  assign n3638 = ( n3634 & n3635 ) | ( n3634 & n3636 ) | ( n3635 & n3636 ) ;
  assign n3639 = ( n3634 & n3637 ) | ( n3634 & ~n3638 ) | ( n3637 & ~n3638 ) ;
  assign n3640 = x29 & x30 ;
  assign n3641 = x13 & x46 ;
  assign n3642 = x28 & x31 ;
  assign n3643 = ( ~n3640 & n3641 ) | ( ~n3640 & n3642 ) | ( n3641 & n3642 ) ;
  assign n3644 = ( n3640 & n3641 ) | ( n3640 & n3642 ) | ( n3641 & n3642 ) ;
  assign n3645 = ( n3640 & n3643 ) | ( n3640 & ~n3644 ) | ( n3643 & ~n3644 ) ;
  assign n3646 = ( ~n3633 & n3639 ) | ( ~n3633 & n3645 ) | ( n3639 & n3645 ) ;
  assign n3647 = ( n3633 & n3639 ) | ( n3633 & n3645 ) | ( n3639 & n3645 ) ;
  assign n3648 = ( n3633 & n3646 ) | ( n3633 & ~n3647 ) | ( n3646 & ~n3647 ) ;
  assign n3649 = ( n3542 & n3627 ) | ( n3542 & n3648 ) | ( n3627 & n3648 ) ;
  assign n3650 = ( ~n3542 & n3627 ) | ( ~n3542 & n3648 ) | ( n3627 & n3648 ) ;
  assign n3651 = ( n3542 & ~n3649 ) | ( n3542 & n3650 ) | ( ~n3649 & n3650 ) ;
  assign n3652 = ( n3564 & ~n3613 ) | ( n3564 & n3651 ) | ( ~n3613 & n3651 ) ;
  assign n3653 = ( n3564 & n3613 ) | ( n3564 & n3651 ) | ( n3613 & n3651 ) ;
  assign n3654 = ( n3613 & n3652 ) | ( n3613 & ~n3653 ) | ( n3652 & ~n3653 ) ;
  assign n3655 = ( ~n3480 & n3504 ) | ( ~n3480 & n3524 ) | ( n3504 & n3524 ) ;
  assign n3656 = ( n3480 & n3504 ) | ( n3480 & n3524 ) | ( n3504 & n3524 ) ;
  assign n3657 = ( n3480 & n3655 ) | ( n3480 & ~n3656 ) | ( n3655 & ~n3656 ) ;
  assign n3658 = ( ~n3477 & n3510 ) | ( ~n3477 & n3516 ) | ( n3510 & n3516 ) ;
  assign n3659 = ( n3477 & n3510 ) | ( n3477 & n3516 ) | ( n3510 & n3516 ) ;
  assign n3660 = ( n3477 & n3658 ) | ( n3477 & ~n3659 ) | ( n3658 & ~n3659 ) ;
  assign n3661 = ( ~n3495 & n3501 ) | ( ~n3495 & n3521 ) | ( n3501 & n3521 ) ;
  assign n3662 = ( n3495 & n3501 ) | ( n3495 & n3521 ) | ( n3501 & n3521 ) ;
  assign n3663 = ( n3495 & n3661 ) | ( n3495 & ~n3662 ) | ( n3661 & ~n3662 ) ;
  assign n3664 = ~x1 & x30 ;
  assign n3665 = ( x1 & x30 ) | ( x1 & x58 ) | ( x30 & x58 ) ;
  assign n3666 = x30 & x58 ;
  assign n3667 = ( n3664 & n3665 ) | ( n3664 & ~n3666 ) | ( n3665 & ~n3666 ) ;
  assign n3668 = ( ~n3465 & n3471 ) | ( ~n3465 & n3667 ) | ( n3471 & n3667 ) ;
  assign n3669 = ( n3465 & n3471 ) | ( n3465 & n3667 ) | ( n3471 & n3667 ) ;
  assign n3670 = ( n3465 & n3668 ) | ( n3465 & ~n3669 ) | ( n3668 & ~n3669 ) ;
  assign n3671 = ( n3660 & n3663 ) | ( n3660 & n3670 ) | ( n3663 & n3670 ) ;
  assign n3672 = ( ~n3660 & n3663 ) | ( ~n3660 & n3670 ) | ( n3663 & n3670 ) ;
  assign n3673 = ( n3660 & ~n3671 ) | ( n3660 & n3672 ) | ( ~n3671 & n3672 ) ;
  assign n3674 = ( n3526 & n3657 ) | ( n3526 & n3673 ) | ( n3657 & n3673 ) ;
  assign n3675 = ( ~n3526 & n3657 ) | ( ~n3526 & n3673 ) | ( n3657 & n3673 ) ;
  assign n3676 = ( n3526 & ~n3674 ) | ( n3526 & n3675 ) | ( ~n3674 & n3675 ) ;
  assign n3677 = ( ~n3566 & n3654 ) | ( ~n3566 & n3676 ) | ( n3654 & n3676 ) ;
  assign n3678 = ( n3566 & n3654 ) | ( n3566 & n3676 ) | ( n3654 & n3676 ) ;
  assign n3679 = ( n3566 & n3677 ) | ( n3566 & ~n3678 ) | ( n3677 & ~n3678 ) ;
  assign n3680 = ( ~n3459 & n3546 ) | ( ~n3459 & n3549 ) | ( n3546 & n3549 ) ;
  assign n3681 = ( n3459 & n3546 ) | ( n3459 & n3549 ) | ( n3546 & n3549 ) ;
  assign n3682 = ( n3459 & n3680 ) | ( n3459 & ~n3681 ) | ( n3680 & ~n3681 ) ;
  assign n3683 = ( n3483 & n3551 ) | ( n3483 & n3682 ) | ( n3551 & n3682 ) ;
  assign n3684 = ( n3483 & n3551 ) | ( n3483 & ~n3682 ) | ( n3551 & ~n3682 ) ;
  assign n3685 = ( n3682 & ~n3683 ) | ( n3682 & n3684 ) | ( ~n3683 & n3684 ) ;
  assign n3686 = ( ~n3529 & n3554 ) | ( ~n3529 & n3685 ) | ( n3554 & n3685 ) ;
  assign n3687 = ( n3529 & n3554 ) | ( n3529 & n3685 ) | ( n3554 & n3685 ) ;
  assign n3688 = ( n3529 & n3686 ) | ( n3529 & ~n3687 ) | ( n3686 & ~n3687 ) ;
  assign n3689 = ( n3557 & ~n3679 ) | ( n3557 & n3688 ) | ( ~n3679 & n3688 ) ;
  assign n3690 = ( n3557 & n3679 ) | ( n3557 & n3688 ) | ( n3679 & n3688 ) ;
  assign n3691 = ( n3679 & n3689 ) | ( n3679 & ~n3690 ) | ( n3689 & ~n3690 ) ;
  assign n3692 = ( n3570 & n3572 ) | ( n3570 & n3691 ) | ( n3572 & n3691 ) ;
  assign n3693 = ( n3570 & ~n3572 ) | ( n3570 & n3691 ) | ( ~n3572 & n3691 ) ;
  assign n3694 = ( n3572 & ~n3692 ) | ( n3572 & n3693 ) | ( ~n3692 & n3693 ) ;
  assign n3695 = x4 & x56 ;
  assign n3696 = x2 & x58 ;
  assign n3697 = x3 & x57 ;
  assign n3698 = ( ~n3695 & n3696 ) | ( ~n3695 & n3697 ) | ( n3696 & n3697 ) ;
  assign n3699 = ( n3695 & n3696 ) | ( n3695 & n3697 ) | ( n3696 & n3697 ) ;
  assign n3700 = ( n3695 & n3698 ) | ( n3695 & ~n3699 ) | ( n3698 & ~n3699 ) ;
  assign n3701 = x22 & x38 ;
  assign n3702 = x20 & x40 ;
  assign n3703 = ( ~n1911 & n3701 ) | ( ~n1911 & n3702 ) | ( n3701 & n3702 ) ;
  assign n3704 = ( n1911 & n3701 ) | ( n1911 & n3702 ) | ( n3701 & n3702 ) ;
  assign n3705 = ( n1911 & n3703 ) | ( n1911 & ~n3704 ) | ( n3703 & ~n3704 ) ;
  assign n3706 = x26 & x34 ;
  assign n3707 = x25 & x35 ;
  assign n3708 = x24 & x36 ;
  assign n3709 = ( ~n3706 & n3707 ) | ( ~n3706 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3710 = ( n3706 & n3707 ) | ( n3706 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3711 = ( n3706 & n3709 ) | ( n3706 & ~n3710 ) | ( n3709 & ~n3710 ) ;
  assign n3712 = ( ~n3700 & n3705 ) | ( ~n3700 & n3711 ) | ( n3705 & n3711 ) ;
  assign n3713 = ( n3700 & n3705 ) | ( n3700 & n3711 ) | ( n3705 & n3711 ) ;
  assign n3714 = ( n3700 & n3712 ) | ( n3700 & ~n3713 ) | ( n3712 & ~n3713 ) ;
  assign n3715 = x15 & x45 ;
  assign n3716 = x10 & x50 ;
  assign n3717 = x11 & x49 ;
  assign n3718 = ( ~n3715 & n3716 ) | ( ~n3715 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3719 = ( n3715 & n3716 ) | ( n3715 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3720 = ( n3715 & n3718 ) | ( n3715 & ~n3719 ) | ( n3718 & ~n3719 ) ;
  assign n3721 = x16 & x44 ;
  assign n3722 = x9 & x51 ;
  assign n3723 = x17 & x43 ;
  assign n3724 = ( ~n3721 & n3722 ) | ( ~n3721 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = ( n3721 & n3722 ) | ( n3721 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3726 = ( n3721 & n3724 ) | ( n3721 & ~n3725 ) | ( n3724 & ~n3725 ) ;
  assign n3727 = ( ~n3638 & n3720 ) | ( ~n3638 & n3726 ) | ( n3720 & n3726 ) ;
  assign n3728 = ( n3638 & n3720 ) | ( n3638 & n3726 ) | ( n3720 & n3726 ) ;
  assign n3729 = ( n3638 & n3727 ) | ( n3638 & ~n3728 ) | ( n3727 & ~n3728 ) ;
  assign n3730 = ( n3681 & n3714 ) | ( n3681 & n3729 ) | ( n3714 & n3729 ) ;
  assign n3731 = ( ~n3681 & n3714 ) | ( ~n3681 & n3729 ) | ( n3714 & n3729 ) ;
  assign n3732 = ( n3681 & ~n3730 ) | ( n3681 & n3731 ) | ( ~n3730 & n3731 ) ;
  assign n3733 = x29 & x31 ;
  assign n3734 = x1 & x59 ;
  assign n3735 = n3733 | n3734 ;
  assign n3736 = x31 & x59 ;
  assign n3737 = n970 & n3736 ;
  assign n3738 = n3735 & ~n3737 ;
  assign n3739 = x58 & n1037 ;
  assign n3740 = x0 & x60 ;
  assign n3741 = ( n3738 & n3739 ) | ( n3738 & n3740 ) | ( n3739 & n3740 ) ;
  assign n3742 = ( ~n3738 & n3739 ) | ( ~n3738 & n3740 ) | ( n3739 & n3740 ) ;
  assign n3743 = ( n3738 & ~n3741 ) | ( n3738 & n3742 ) | ( ~n3741 & n3742 ) ;
  assign n3744 = x28 & x32 ;
  assign n3745 = x23 & x37 ;
  assign n3746 = x27 & x33 ;
  assign n3747 = ( ~n3744 & n3745 ) | ( ~n3744 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3748 = ( n3744 & n3745 ) | ( n3744 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3749 = ( n3744 & n3747 ) | ( n3744 & ~n3748 ) | ( n3747 & ~n3748 ) ;
  assign n3750 = ( n3669 & n3743 ) | ( n3669 & n3749 ) | ( n3743 & n3749 ) ;
  assign n3751 = ( n3669 & ~n3743 ) | ( n3669 & n3749 ) | ( ~n3743 & n3749 ) ;
  assign n3752 = ( n3743 & ~n3750 ) | ( n3743 & n3751 ) | ( ~n3750 & n3751 ) ;
  assign n3753 = x14 & x46 ;
  assign n3754 = x12 & x48 ;
  assign n3755 = x13 & x47 ;
  assign n3756 = ( ~n3753 & n3754 ) | ( ~n3753 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3757 = ( n3753 & n3754 ) | ( n3753 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3758 = ( n3753 & n3756 ) | ( n3753 & ~n3757 ) | ( n3756 & ~n3757 ) ;
  assign n3759 = x8 & x52 ;
  assign n3760 = x7 & x53 ;
  assign n3761 = x18 & x42 ;
  assign n3762 = ( ~n3759 & n3760 ) | ( ~n3759 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = ( n3759 & n3760 ) | ( n3759 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3764 = ( n3759 & n3762 ) | ( n3759 & ~n3763 ) | ( n3762 & ~n3763 ) ;
  assign n3765 = x6 & x54 ;
  assign n3766 = x5 & x55 ;
  assign n3767 = x19 & x41 ;
  assign n3768 = ( ~n3765 & n3766 ) | ( ~n3765 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3769 = ( n3765 & n3766 ) | ( n3765 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3770 = ( n3765 & n3768 ) | ( n3765 & ~n3769 ) | ( n3768 & ~n3769 ) ;
  assign n3771 = ( ~n3758 & n3764 ) | ( ~n3758 & n3770 ) | ( n3764 & n3770 ) ;
  assign n3772 = ( n3758 & n3764 ) | ( n3758 & n3770 ) | ( n3764 & n3770 ) ;
  assign n3773 = ( n3758 & n3771 ) | ( n3758 & ~n3772 ) | ( n3771 & ~n3772 ) ;
  assign n3774 = ( n3671 & n3752 ) | ( n3671 & n3773 ) | ( n3752 & n3773 ) ;
  assign n3775 = ( n3671 & ~n3752 ) | ( n3671 & n3773 ) | ( ~n3752 & n3773 ) ;
  assign n3776 = ( n3752 & ~n3774 ) | ( n3752 & n3775 ) | ( ~n3774 & n3775 ) ;
  assign n3777 = ( ~n3683 & n3732 ) | ( ~n3683 & n3776 ) | ( n3732 & n3776 ) ;
  assign n3778 = ( n3683 & n3732 ) | ( n3683 & n3776 ) | ( n3732 & n3776 ) ;
  assign n3779 = ( n3683 & n3777 ) | ( n3683 & ~n3778 ) | ( n3777 & ~n3778 ) ;
  assign n3780 = ( n3585 & n3594 ) | ( n3585 & ~n3617 ) | ( n3594 & ~n3617 ) ;
  assign n3781 = ( n3585 & n3594 ) | ( n3585 & n3617 ) | ( n3594 & n3617 ) ;
  assign n3782 = ( n3617 & n3780 ) | ( n3617 & ~n3781 ) | ( n3780 & ~n3781 ) ;
  assign n3783 = ( n3600 & n3606 ) | ( n3600 & ~n3623 ) | ( n3606 & ~n3623 ) ;
  assign n3784 = ( n3600 & n3606 ) | ( n3600 & n3623 ) | ( n3606 & n3623 ) ;
  assign n3785 = ( n3623 & n3783 ) | ( n3623 & ~n3784 ) | ( n3783 & ~n3784 ) ;
  assign n3786 = ( n3588 & n3782 ) | ( n3588 & n3785 ) | ( n3782 & n3785 ) ;
  assign n3787 = ( ~n3588 & n3782 ) | ( ~n3588 & n3785 ) | ( n3782 & n3785 ) ;
  assign n3788 = ( n3588 & ~n3786 ) | ( n3588 & n3787 ) | ( ~n3786 & n3787 ) ;
  assign n3789 = ( n3579 & ~n3632 ) | ( n3579 & n3644 ) | ( ~n3632 & n3644 ) ;
  assign n3790 = ( n3579 & n3632 ) | ( n3579 & n3644 ) | ( n3632 & n3644 ) ;
  assign n3791 = ( n3632 & n3789 ) | ( n3632 & ~n3790 ) | ( n3789 & ~n3790 ) ;
  assign n3792 = ( n3609 & n3647 ) | ( n3609 & n3791 ) | ( n3647 & n3791 ) ;
  assign n3793 = ( n3609 & ~n3647 ) | ( n3609 & n3791 ) | ( ~n3647 & n3791 ) ;
  assign n3794 = ( n3647 & ~n3792 ) | ( n3647 & n3793 ) | ( ~n3792 & n3793 ) ;
  assign n3795 = ( n3649 & n3788 ) | ( n3649 & n3794 ) | ( n3788 & n3794 ) ;
  assign n3796 = ( n3649 & ~n3788 ) | ( n3649 & n3794 ) | ( ~n3788 & n3794 ) ;
  assign n3797 = ( n3788 & ~n3795 ) | ( n3788 & n3796 ) | ( ~n3795 & n3796 ) ;
  assign n3798 = ( n3687 & n3779 ) | ( n3687 & n3797 ) | ( n3779 & n3797 ) ;
  assign n3799 = ( ~n3687 & n3779 ) | ( ~n3687 & n3797 ) | ( n3779 & n3797 ) ;
  assign n3800 = ( n3687 & ~n3798 ) | ( n3687 & n3799 ) | ( ~n3798 & n3799 ) ;
  assign n3801 = ( ~n3626 & n3659 ) | ( ~n3626 & n3662 ) | ( n3659 & n3662 ) ;
  assign n3802 = ( n3626 & n3659 ) | ( n3626 & n3662 ) | ( n3659 & n3662 ) ;
  assign n3803 = ( n3626 & n3801 ) | ( n3626 & ~n3802 ) | ( n3801 & ~n3802 ) ;
  assign n3804 = ( ~n3611 & n3656 ) | ( ~n3611 & n3803 ) | ( n3656 & n3803 ) ;
  assign n3805 = ( n3611 & n3656 ) | ( n3611 & n3803 ) | ( n3656 & n3803 ) ;
  assign n3806 = ( n3611 & n3804 ) | ( n3611 & ~n3805 ) | ( n3804 & ~n3805 ) ;
  assign n3807 = ( n3653 & n3674 ) | ( n3653 & ~n3806 ) | ( n3674 & ~n3806 ) ;
  assign n3808 = ( n3653 & n3674 ) | ( n3653 & n3806 ) | ( n3674 & n3806 ) ;
  assign n3809 = ( n3806 & n3807 ) | ( n3806 & ~n3808 ) | ( n3807 & ~n3808 ) ;
  assign n3810 = ( n3678 & n3800 ) | ( n3678 & n3809 ) | ( n3800 & n3809 ) ;
  assign n3811 = ( ~n3678 & n3800 ) | ( ~n3678 & n3809 ) | ( n3800 & n3809 ) ;
  assign n3812 = ( n3678 & ~n3810 ) | ( n3678 & n3811 ) | ( ~n3810 & n3811 ) ;
  assign n3813 = ( n3690 & n3692 ) | ( n3690 & n3812 ) | ( n3692 & n3812 ) ;
  assign n3814 = ( n3690 & ~n3692 ) | ( n3690 & n3812 ) | ( ~n3692 & n3812 ) ;
  assign n3815 = ( n3692 & ~n3813 ) | ( n3692 & n3814 ) | ( ~n3813 & n3814 ) ;
  assign n3816 = x1 & x60 ;
  assign n3817 = x31 & ~n3737 ;
  assign n3818 = ( n3737 & n3816 ) | ( n3737 & ~n3817 ) | ( n3816 & ~n3817 ) ;
  assign n3819 = x31 & ~n3816 ;
  assign n3820 = ( n3757 & n3818 ) | ( n3757 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3821 = ( n3757 & ~n3816 ) | ( n3757 & n3817 ) | ( ~n3816 & n3817 ) ;
  assign n3822 = ( n3818 & ~n3820 ) | ( n3818 & n3821 ) | ( ~n3820 & n3821 ) ;
  assign n3823 = ( n3728 & n3784 ) | ( n3728 & ~n3822 ) | ( n3784 & ~n3822 ) ;
  assign n3824 = ( n3728 & n3784 ) | ( n3728 & n3822 ) | ( n3784 & n3822 ) ;
  assign n3825 = ( n3822 & n3823 ) | ( n3822 & ~n3824 ) | ( n3823 & ~n3824 ) ;
  assign n3826 = x3 & x58 ;
  assign n3827 = x4 & x57 ;
  assign n3828 = x23 & x38 ;
  assign n3829 = ( ~n3826 & n3827 ) | ( ~n3826 & n3828 ) | ( n3827 & n3828 ) ;
  assign n3830 = ( n3826 & n3827 ) | ( n3826 & n3828 ) | ( n3827 & n3828 ) ;
  assign n3831 = ( n3826 & n3829 ) | ( n3826 & ~n3830 ) | ( n3829 & ~n3830 ) ;
  assign n3832 = ( ~n3781 & n3790 ) | ( ~n3781 & n3831 ) | ( n3790 & n3831 ) ;
  assign n3833 = ( n3781 & n3790 ) | ( n3781 & n3831 ) | ( n3790 & n3831 ) ;
  assign n3834 = ( n3781 & n3832 ) | ( n3781 & ~n3833 ) | ( n3832 & ~n3833 ) ;
  assign n3835 = ( n3730 & n3825 ) | ( n3730 & n3834 ) | ( n3825 & n3834 ) ;
  assign n3836 = ( ~n3730 & n3825 ) | ( ~n3730 & n3834 ) | ( n3825 & n3834 ) ;
  assign n3837 = ( n3730 & ~n3835 ) | ( n3730 & n3836 ) | ( ~n3835 & n3836 ) ;
  assign n3838 = x19 & x42 ;
  assign n3839 = x7 & x54 ;
  assign n3840 = x8 & x53 ;
  assign n3841 = ( ~n3838 & n3839 ) | ( ~n3838 & n3840 ) | ( n3839 & n3840 ) ;
  assign n3842 = ( n3838 & n3839 ) | ( n3838 & n3840 ) | ( n3839 & n3840 ) ;
  assign n3843 = ( n3838 & n3841 ) | ( n3838 & ~n3842 ) | ( n3841 & ~n3842 ) ;
  assign n3844 = x9 & x52 ;
  assign n3845 = x17 & x44 ;
  assign n3846 = x18 & x43 ;
  assign n3847 = ( ~n3844 & n3845 ) | ( ~n3844 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = ( n3844 & n3845 ) | ( n3844 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3849 = ( n3844 & n3847 ) | ( n3844 & ~n3848 ) | ( n3847 & ~n3848 ) ;
  assign n3850 = x28 & x33 ;
  assign n3851 = x27 & x34 ;
  assign n3852 = x26 & x35 ;
  assign n3853 = ( ~n3850 & n3851 ) | ( ~n3850 & n3852 ) | ( n3851 & n3852 ) ;
  assign n3854 = ( n3850 & n3851 ) | ( n3850 & n3852 ) | ( n3851 & n3852 ) ;
  assign n3855 = ( n3850 & n3853 ) | ( n3850 & ~n3854 ) | ( n3853 & ~n3854 ) ;
  assign n3856 = ( ~n3843 & n3849 ) | ( ~n3843 & n3855 ) | ( n3849 & n3855 ) ;
  assign n3857 = ( n3843 & n3849 ) | ( n3843 & n3855 ) | ( n3849 & n3855 ) ;
  assign n3858 = ( n3843 & n3856 ) | ( n3843 & ~n3857 ) | ( n3856 & ~n3857 ) ;
  assign n3859 = ( n3786 & n3792 ) | ( n3786 & n3858 ) | ( n3792 & n3858 ) ;
  assign n3860 = ( ~n3786 & n3792 ) | ( ~n3786 & n3858 ) | ( n3792 & n3858 ) ;
  assign n3861 = ( n3786 & ~n3859 ) | ( n3786 & n3860 ) | ( ~n3859 & n3860 ) ;
  assign n3862 = ( n3778 & n3837 ) | ( n3778 & n3861 ) | ( n3837 & n3861 ) ;
  assign n3863 = ( ~n3778 & n3837 ) | ( ~n3778 & n3861 ) | ( n3837 & n3861 ) ;
  assign n3864 = ( n3778 & ~n3862 ) | ( n3778 & n3863 ) | ( ~n3862 & n3863 ) ;
  assign n3865 = x24 & x37 ;
  assign n3866 = x22 & x39 ;
  assign n3867 = x25 & x36 ;
  assign n3868 = ( ~n3865 & n3866 ) | ( ~n3865 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = ( n3865 & n3866 ) | ( n3865 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3870 = ( n3865 & n3868 ) | ( n3865 & ~n3869 ) | ( n3868 & ~n3869 ) ;
  assign n3871 = x20 & x41 ;
  assign n3872 = x6 & x55 ;
  assign n3873 = ( ~n1826 & n3871 ) | ( ~n1826 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3874 = ( n1826 & n3871 ) | ( n1826 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3875 = ( n1826 & n3873 ) | ( n1826 & ~n3874 ) | ( n3873 & ~n3874 ) ;
  assign n3876 = x0 & x61 ;
  assign n3877 = x2 & x59 ;
  assign n3878 = x5 & x56 ;
  assign n3879 = ( ~n3876 & n3877 ) | ( ~n3876 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3880 = ( n3876 & n3877 ) | ( n3876 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3881 = ( n3876 & n3879 ) | ( n3876 & ~n3880 ) | ( n3879 & ~n3880 ) ;
  assign n3882 = ( ~n3870 & n3875 ) | ( ~n3870 & n3881 ) | ( n3875 & n3881 ) ;
  assign n3883 = ( n3870 & n3875 ) | ( n3870 & n3881 ) | ( n3875 & n3881 ) ;
  assign n3884 = ( n3870 & n3882 ) | ( n3870 & ~n3883 ) | ( n3882 & ~n3883 ) ;
  assign n3885 = x30 & x31 ;
  assign n3886 = x13 & x48 ;
  assign n3887 = x29 & x32 ;
  assign n3888 = ( ~n3885 & n3886 ) | ( ~n3885 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ( n3885 & n3886 ) | ( n3885 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3890 = ( n3885 & n3888 ) | ( n3885 & ~n3889 ) | ( n3888 & ~n3889 ) ;
  assign n3891 = x11 & x50 ;
  assign n3892 = x14 & x47 ;
  assign n3893 = x12 & x49 ;
  assign n3894 = ( ~n3891 & n3892 ) | ( ~n3891 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3895 = ( n3891 & n3892 ) | ( n3891 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3896 = ( n3891 & n3894 ) | ( n3891 & ~n3895 ) | ( n3894 & ~n3895 ) ;
  assign n3897 = x16 & x45 ;
  assign n3898 = x15 & x46 ;
  assign n3899 = x10 & x51 ;
  assign n3900 = ( ~n3897 & n3898 ) | ( ~n3897 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3901 = ( n3897 & n3898 ) | ( n3897 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3902 = ( n3897 & n3900 ) | ( n3897 & ~n3901 ) | ( n3900 & ~n3901 ) ;
  assign n3903 = ( ~n3890 & n3896 ) | ( ~n3890 & n3902 ) | ( n3896 & n3902 ) ;
  assign n3904 = ( n3890 & n3896 ) | ( n3890 & n3902 ) | ( n3896 & n3902 ) ;
  assign n3905 = ( n3890 & n3903 ) | ( n3890 & ~n3904 ) | ( n3903 & ~n3904 ) ;
  assign n3906 = ( n3802 & n3884 ) | ( n3802 & n3905 ) | ( n3884 & n3905 ) ;
  assign n3907 = ( ~n3802 & n3884 ) | ( ~n3802 & n3905 ) | ( n3884 & n3905 ) ;
  assign n3908 = ( n3802 & ~n3906 ) | ( n3802 & n3907 ) | ( ~n3906 & n3907 ) ;
  assign n3909 = ( n3795 & n3805 ) | ( n3795 & n3908 ) | ( n3805 & n3908 ) ;
  assign n3910 = ( ~n3795 & n3805 ) | ( ~n3795 & n3908 ) | ( n3805 & n3908 ) ;
  assign n3911 = ( n3795 & ~n3909 ) | ( n3795 & n3910 ) | ( ~n3909 & n3910 ) ;
  assign n3912 = ( n3725 & ~n3741 ) | ( n3725 & n3763 ) | ( ~n3741 & n3763 ) ;
  assign n3913 = ( n3725 & n3741 ) | ( n3725 & n3763 ) | ( n3741 & n3763 ) ;
  assign n3914 = ( n3741 & n3912 ) | ( n3741 & ~n3913 ) | ( n3912 & ~n3913 ) ;
  assign n3915 = ( n3750 & n3772 ) | ( n3750 & n3914 ) | ( n3772 & n3914 ) ;
  assign n3916 = ( n3750 & n3772 ) | ( n3750 & ~n3914 ) | ( n3772 & ~n3914 ) ;
  assign n3917 = ( n3914 & ~n3915 ) | ( n3914 & n3916 ) | ( ~n3915 & n3916 ) ;
  assign n3918 = ( n3704 & n3710 ) | ( n3704 & ~n3748 ) | ( n3710 & ~n3748 ) ;
  assign n3919 = ( n3704 & n3710 ) | ( n3704 & n3748 ) | ( n3710 & n3748 ) ;
  assign n3920 = ( n3748 & n3918 ) | ( n3748 & ~n3919 ) | ( n3918 & ~n3919 ) ;
  assign n3921 = ( n3699 & n3719 ) | ( n3699 & ~n3769 ) | ( n3719 & ~n3769 ) ;
  assign n3922 = ( n3699 & n3719 ) | ( n3699 & n3769 ) | ( n3719 & n3769 ) ;
  assign n3923 = ( n3769 & n3921 ) | ( n3769 & ~n3922 ) | ( n3921 & ~n3922 ) ;
  assign n3924 = ( n3713 & n3920 ) | ( n3713 & n3923 ) | ( n3920 & n3923 ) ;
  assign n3925 = ( n3713 & ~n3920 ) | ( n3713 & n3923 ) | ( ~n3920 & n3923 ) ;
  assign n3926 = ( n3920 & ~n3924 ) | ( n3920 & n3925 ) | ( ~n3924 & n3925 ) ;
  assign n3927 = ( ~n3774 & n3917 ) | ( ~n3774 & n3926 ) | ( n3917 & n3926 ) ;
  assign n3928 = ( n3774 & n3917 ) | ( n3774 & n3926 ) | ( n3917 & n3926 ) ;
  assign n3929 = ( n3774 & n3927 ) | ( n3774 & ~n3928 ) | ( n3927 & ~n3928 ) ;
  assign n3930 = ( n3808 & ~n3911 ) | ( n3808 & n3929 ) | ( ~n3911 & n3929 ) ;
  assign n3931 = ( n3808 & n3911 ) | ( n3808 & n3929 ) | ( n3911 & n3929 ) ;
  assign n3932 = ( n3911 & n3930 ) | ( n3911 & ~n3931 ) | ( n3930 & ~n3931 ) ;
  assign n3933 = ( ~n3798 & n3864 ) | ( ~n3798 & n3932 ) | ( n3864 & n3932 ) ;
  assign n3934 = ( n3798 & n3864 ) | ( n3798 & n3932 ) | ( n3864 & n3932 ) ;
  assign n3935 = ( n3798 & n3933 ) | ( n3798 & ~n3934 ) | ( n3933 & ~n3934 ) ;
  assign n3936 = ( n3810 & n3813 ) | ( n3810 & n3935 ) | ( n3813 & n3935 ) ;
  assign n3937 = ( n3810 & ~n3813 ) | ( n3810 & n3935 ) | ( ~n3813 & n3935 ) ;
  assign n3938 = ( n3813 & ~n3936 ) | ( n3813 & n3937 ) | ( ~n3936 & n3937 ) ;
  assign n3939 = ( n3883 & n3904 ) | ( n3883 & ~n3922 ) | ( n3904 & ~n3922 ) ;
  assign n3940 = ( n3883 & n3904 ) | ( n3883 & n3922 ) | ( n3904 & n3922 ) ;
  assign n3941 = ( n3922 & n3939 ) | ( n3922 & ~n3940 ) | ( n3939 & ~n3940 ) ;
  assign n3942 = ( n3830 & n3854 ) | ( n3830 & ~n3869 ) | ( n3854 & ~n3869 ) ;
  assign n3943 = ( n3830 & n3854 ) | ( n3830 & n3869 ) | ( n3854 & n3869 ) ;
  assign n3944 = ( n3869 & n3942 ) | ( n3869 & ~n3943 ) | ( n3942 & ~n3943 ) ;
  assign n3945 = x30 & x32 ;
  assign n3946 = x1 & x61 ;
  assign n3947 = n3945 & n3946 ;
  assign n3948 = n3945 | n3946 ;
  assign n3949 = ~n3947 & n3948 ;
  assign n3950 = ( ~n3889 & n3895 ) | ( ~n3889 & n3949 ) | ( n3895 & n3949 ) ;
  assign n3951 = ( n3889 & n3895 ) | ( n3889 & n3949 ) | ( n3895 & n3949 ) ;
  assign n3952 = ( n3889 & n3950 ) | ( n3889 & ~n3951 ) | ( n3950 & ~n3951 ) ;
  assign n3953 = ( n3842 & ~n3874 ) | ( n3842 & n3880 ) | ( ~n3874 & n3880 ) ;
  assign n3954 = ( n3842 & n3874 ) | ( n3842 & n3880 ) | ( n3874 & n3880 ) ;
  assign n3955 = ( n3874 & n3953 ) | ( n3874 & ~n3954 ) | ( n3953 & ~n3954 ) ;
  assign n3956 = ( n3944 & n3952 ) | ( n3944 & n3955 ) | ( n3952 & n3955 ) ;
  assign n3957 = ( ~n3944 & n3952 ) | ( ~n3944 & n3955 ) | ( n3952 & n3955 ) ;
  assign n3958 = ( n3944 & ~n3956 ) | ( n3944 & n3957 ) | ( ~n3956 & n3957 ) ;
  assign n3959 = ( n3859 & n3941 ) | ( n3859 & n3958 ) | ( n3941 & n3958 ) ;
  assign n3960 = ( ~n3859 & n3941 ) | ( ~n3859 & n3958 ) | ( n3941 & n3958 ) ;
  assign n3961 = ( n3859 & ~n3959 ) | ( n3859 & n3960 ) | ( ~n3959 & n3960 ) ;
  assign n3962 = ( n3824 & n3915 ) | ( n3824 & n3924 ) | ( n3915 & n3924 ) ;
  assign n3963 = ( n3824 & ~n3915 ) | ( n3824 & n3924 ) | ( ~n3915 & n3924 ) ;
  assign n3964 = ( n3915 & ~n3962 ) | ( n3915 & n3963 ) | ( ~n3962 & n3963 ) ;
  assign n3965 = ( n3909 & n3961 ) | ( n3909 & n3964 ) | ( n3961 & n3964 ) ;
  assign n3966 = ( ~n3909 & n3961 ) | ( ~n3909 & n3964 ) | ( n3961 & n3964 ) ;
  assign n3967 = ( n3909 & ~n3965 ) | ( n3909 & n3966 ) | ( ~n3965 & n3966 ) ;
  assign n3968 = x3 & x59 ;
  assign n3969 = x4 & x58 ;
  assign n3970 = x5 & x57 ;
  assign n3971 = ( ~n3968 & n3969 ) | ( ~n3968 & n3970 ) | ( n3969 & n3970 ) ;
  assign n3972 = ( n3968 & n3969 ) | ( n3968 & n3970 ) | ( n3969 & n3970 ) ;
  assign n3973 = ( n3968 & n3971 ) | ( n3968 & ~n3972 ) | ( n3971 & ~n3972 ) ;
  assign n3974 = ( n3848 & n3901 ) | ( n3848 & ~n3973 ) | ( n3901 & ~n3973 ) ;
  assign n3975 = ( n3848 & n3901 ) | ( n3848 & n3973 ) | ( n3901 & n3973 ) ;
  assign n3976 = ( n3973 & n3974 ) | ( n3973 & ~n3975 ) | ( n3974 & ~n3975 ) ;
  assign n3977 = ( n3833 & n3857 ) | ( n3833 & n3976 ) | ( n3857 & n3976 ) ;
  assign n3978 = ( n3833 & n3857 ) | ( n3833 & ~n3976 ) | ( n3857 & ~n3976 ) ;
  assign n3979 = ( n3976 & ~n3977 ) | ( n3976 & n3978 ) | ( ~n3977 & n3978 ) ;
  assign n3980 = ( ~n3820 & n3913 ) | ( ~n3820 & n3919 ) | ( n3913 & n3919 ) ;
  assign n3981 = ( n3820 & n3913 ) | ( n3820 & n3919 ) | ( n3913 & n3919 ) ;
  assign n3982 = ( n3820 & n3980 ) | ( n3820 & ~n3981 ) | ( n3980 & ~n3981 ) ;
  assign n3983 = ( ~n3906 & n3979 ) | ( ~n3906 & n3982 ) | ( n3979 & n3982 ) ;
  assign n3984 = ( n3906 & n3979 ) | ( n3906 & n3982 ) | ( n3979 & n3982 ) ;
  assign n3985 = ( n3906 & n3983 ) | ( n3906 & ~n3984 ) | ( n3983 & ~n3984 ) ;
  assign n3986 = ( x2 & ~x60 ) | ( x2 & n1098 ) | ( ~x60 & n1098 ) ;
  assign n3987 = x0 & x62 ;
  assign n3988 = x2 | n1098 ;
  assign n3989 = ( ~n3986 & n3987 ) | ( ~n3986 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3990 = ( n3986 & n3987 ) | ( n3986 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3991 = ( n3986 & n3989 ) | ( n3986 & ~n3990 ) | ( n3989 & ~n3990 ) ;
  assign n3992 = x9 & x53 ;
  assign n3993 = x17 & x45 ;
  assign n3994 = x10 & x52 ;
  assign n3995 = ( ~n3992 & n3993 ) | ( ~n3992 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3996 = ( n3992 & n3993 ) | ( n3992 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3997 = ( n3992 & n3995 ) | ( n3992 & ~n3996 ) | ( n3995 & ~n3996 ) ;
  assign n3998 = x25 & x37 ;
  assign n3999 = x21 & x41 ;
  assign n4000 = x26 & x36 ;
  assign n4001 = ( ~n3998 & n3999 ) | ( ~n3998 & n4000 ) | ( n3999 & n4000 ) ;
  assign n4002 = ( n3998 & n3999 ) | ( n3998 & n4000 ) | ( n3999 & n4000 ) ;
  assign n4003 = ( n3998 & n4001 ) | ( n3998 & ~n4002 ) | ( n4001 & ~n4002 ) ;
  assign n4004 = ( ~n3991 & n3997 ) | ( ~n3991 & n4003 ) | ( n3997 & n4003 ) ;
  assign n4005 = ( n3991 & n3997 ) | ( n3991 & n4003 ) | ( n3997 & n4003 ) ;
  assign n4006 = ( n3991 & n4004 ) | ( n3991 & ~n4005 ) | ( n4004 & ~n4005 ) ;
  assign n4007 = x27 & x35 ;
  assign n4008 = x28 & x34 ;
  assign n4009 = x29 & x33 ;
  assign n4010 = ( ~n4007 & n4008 ) | ( ~n4007 & n4009 ) | ( n4008 & n4009 ) ;
  assign n4011 = ( n4007 & n4008 ) | ( n4007 & n4009 ) | ( n4008 & n4009 ) ;
  assign n4012 = ( n4007 & n4010 ) | ( n4007 & ~n4011 ) | ( n4010 & ~n4011 ) ;
  assign n4013 = x8 & x54 ;
  assign n4014 = x18 & x44 ;
  assign n4015 = x19 & x43 ;
  assign n4016 = ( ~n4013 & n4014 ) | ( ~n4013 & n4015 ) | ( n4014 & n4015 ) ;
  assign n4017 = ( n4013 & n4014 ) | ( n4013 & n4015 ) | ( n4014 & n4015 ) ;
  assign n4018 = ( n4013 & n4016 ) | ( n4013 & ~n4017 ) | ( n4016 & ~n4017 ) ;
  assign n4019 = x23 & x39 ;
  assign n4020 = x22 & x40 ;
  assign n4021 = x24 & x38 ;
  assign n4022 = ( ~n4019 & n4020 ) | ( ~n4019 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4023 = ( n4019 & n4020 ) | ( n4019 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4024 = ( n4019 & n4022 ) | ( n4019 & ~n4023 ) | ( n4022 & ~n4023 ) ;
  assign n4025 = ( ~n4012 & n4018 ) | ( ~n4012 & n4024 ) | ( n4018 & n4024 ) ;
  assign n4026 = ( n4012 & n4018 ) | ( n4012 & n4024 ) | ( n4018 & n4024 ) ;
  assign n4027 = ( n4012 & n4025 ) | ( n4012 & ~n4026 ) | ( n4025 & ~n4026 ) ;
  assign n4028 = x15 & x47 ;
  assign n4029 = x11 & x51 ;
  assign n4030 = x16 & x46 ;
  assign n4031 = ( ~n4028 & n4029 ) | ( ~n4028 & n4030 ) | ( n4029 & n4030 ) ;
  assign n4032 = ( n4028 & n4029 ) | ( n4028 & n4030 ) | ( n4029 & n4030 ) ;
  assign n4033 = ( n4028 & n4031 ) | ( n4028 & ~n4032 ) | ( n4031 & ~n4032 ) ;
  assign n4034 = x12 & x50 ;
  assign n4035 = x13 & x49 ;
  assign n4036 = x14 & x48 ;
  assign n4037 = ( ~n4034 & n4035 ) | ( ~n4034 & n4036 ) | ( n4035 & n4036 ) ;
  assign n4038 = ( n4034 & n4035 ) | ( n4034 & n4036 ) | ( n4035 & n4036 ) ;
  assign n4039 = ( n4034 & n4037 ) | ( n4034 & ~n4038 ) | ( n4037 & ~n4038 ) ;
  assign n4040 = x7 & x55 ;
  assign n4041 = x20 & x42 ;
  assign n4042 = x6 & x56 ;
  assign n4043 = ( ~n4040 & n4041 ) | ( ~n4040 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4044 = ( n4040 & n4041 ) | ( n4040 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4045 = ( n4040 & n4043 ) | ( n4040 & ~n4044 ) | ( n4043 & ~n4044 ) ;
  assign n4046 = ( ~n4033 & n4039 ) | ( ~n4033 & n4045 ) | ( n4039 & n4045 ) ;
  assign n4047 = ( n4033 & n4039 ) | ( n4033 & n4045 ) | ( n4039 & n4045 ) ;
  assign n4048 = ( n4033 & n4046 ) | ( n4033 & ~n4047 ) | ( n4046 & ~n4047 ) ;
  assign n4049 = ( ~n4006 & n4027 ) | ( ~n4006 & n4048 ) | ( n4027 & n4048 ) ;
  assign n4050 = ( n4006 & n4027 ) | ( n4006 & n4048 ) | ( n4027 & n4048 ) ;
  assign n4051 = ( n4006 & n4049 ) | ( n4006 & ~n4050 ) | ( n4049 & ~n4050 ) ;
  assign n4052 = ( n3835 & ~n3928 ) | ( n3835 & n4051 ) | ( ~n3928 & n4051 ) ;
  assign n4053 = ( n3835 & n3928 ) | ( n3835 & n4051 ) | ( n3928 & n4051 ) ;
  assign n4054 = ( n3928 & n4052 ) | ( n3928 & ~n4053 ) | ( n4052 & ~n4053 ) ;
  assign n4055 = ( ~n3862 & n3985 ) | ( ~n3862 & n4054 ) | ( n3985 & n4054 ) ;
  assign n4056 = ( n3862 & n3985 ) | ( n3862 & n4054 ) | ( n3985 & n4054 ) ;
  assign n4057 = ( n3862 & n4055 ) | ( n3862 & ~n4056 ) | ( n4055 & ~n4056 ) ;
  assign n4058 = ( n3931 & n3967 ) | ( n3931 & n4057 ) | ( n3967 & n4057 ) ;
  assign n4059 = ( ~n3931 & n3967 ) | ( ~n3931 & n4057 ) | ( n3967 & n4057 ) ;
  assign n4060 = ( n3931 & ~n4058 ) | ( n3931 & n4059 ) | ( ~n4058 & n4059 ) ;
  assign n4061 = ( n3934 & n3936 ) | ( n3934 & n4060 ) | ( n3936 & n4060 ) ;
  assign n4062 = ( n3934 & ~n3936 ) | ( n3934 & n4060 ) | ( ~n3936 & n4060 ) ;
  assign n4063 = ( n3936 & ~n4061 ) | ( n3936 & n4062 ) | ( ~n4061 & n4062 ) ;
  assign n4064 = x3 & x60 ;
  assign n4065 = x2 & x61 ;
  assign n4066 = x4 & x59 ;
  assign n4067 = ( ~n4064 & n4065 ) | ( ~n4064 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4068 = ( n4064 & n4065 ) | ( n4064 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4069 = ( n4064 & n4067 ) | ( n4064 & ~n4068 ) | ( n4067 & ~n4068 ) ;
  assign n4070 = x5 & x58 ;
  assign n4071 = x21 & x42 ;
  assign n4072 = ( ~n1893 & n4070 ) | ( ~n1893 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4073 = ( n1893 & n4070 ) | ( n1893 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4074 = ( n1893 & n4072 ) | ( n1893 & ~n4073 ) | ( n4072 & ~n4073 ) ;
  assign n4075 = ( ~n4032 & n4069 ) | ( ~n4032 & n4074 ) | ( n4069 & n4074 ) ;
  assign n4076 = ( n4032 & n4069 ) | ( n4032 & n4074 ) | ( n4069 & n4074 ) ;
  assign n4077 = ( n4032 & n4075 ) | ( n4032 & ~n4076 ) | ( n4075 & ~n4076 ) ;
  assign n4078 = x30 & x33 ;
  assign n4079 = x31 & x32 ;
  assign n4080 = x14 & x49 ;
  assign n4081 = ( ~n4078 & n4079 ) | ( ~n4078 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4082 = ( n4078 & n4079 ) | ( n4078 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4083 = ( n4078 & n4081 ) | ( n4078 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  assign n4084 = x23 & x40 ;
  assign n4085 = x20 & x43 ;
  assign n4086 = x6 & x57 ;
  assign n4087 = ( ~n4084 & n4085 ) | ( ~n4084 & n4086 ) | ( n4085 & n4086 ) ;
  assign n4088 = ( n4084 & n4085 ) | ( n4084 & n4086 ) | ( n4085 & n4086 ) ;
  assign n4089 = ( n4084 & n4087 ) | ( n4084 & ~n4088 ) | ( n4087 & ~n4088 ) ;
  assign n4090 = x8 & x55 ;
  assign n4091 = x7 & x56 ;
  assign n4092 = x19 & x44 ;
  assign n4093 = ( ~n4090 & n4091 ) | ( ~n4090 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4094 = ( n4090 & n4091 ) | ( n4090 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4095 = ( n4090 & n4093 ) | ( n4090 & ~n4094 ) | ( n4093 & ~n4094 ) ;
  assign n4096 = ( ~n4083 & n4089 ) | ( ~n4083 & n4095 ) | ( n4089 & n4095 ) ;
  assign n4097 = ( n4083 & n4089 ) | ( n4083 & n4095 ) | ( n4089 & n4095 ) ;
  assign n4098 = ( n4083 & n4096 ) | ( n4083 & ~n4097 ) | ( n4096 & ~n4097 ) ;
  assign n4099 = x9 & x54 ;
  assign n4100 = x18 & x45 ;
  assign n4101 = x17 & x46 ;
  assign n4102 = ( ~n4099 & n4100 ) | ( ~n4099 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = ( n4099 & n4100 ) | ( n4099 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4104 = ( n4099 & n4102 ) | ( n4099 & ~n4103 ) | ( n4102 & ~n4103 ) ;
  assign n4105 = x11 & x52 ;
  assign n4106 = x10 & x53 ;
  assign n4107 = x16 & x47 ;
  assign n4108 = ( ~n4105 & n4106 ) | ( ~n4105 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = ( n4105 & n4106 ) | ( n4105 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4110 = ( n4105 & n4108 ) | ( n4105 & ~n4109 ) | ( n4108 & ~n4109 ) ;
  assign n4111 = x15 & x48 ;
  assign n4112 = x13 & x50 ;
  assign n4113 = x12 & x51 ;
  assign n4114 = ( ~n4111 & n4112 ) | ( ~n4111 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n4111 & n4112 ) | ( n4111 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4116 = ( n4111 & n4114 ) | ( n4111 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = ( ~n4104 & n4110 ) | ( ~n4104 & n4116 ) | ( n4110 & n4116 ) ;
  assign n4118 = ( n4104 & n4110 ) | ( n4104 & n4116 ) | ( n4110 & n4116 ) ;
  assign n4119 = ( n4104 & n4117 ) | ( n4104 & ~n4118 ) | ( n4117 & ~n4118 ) ;
  assign n4120 = ( ~n4077 & n4098 ) | ( ~n4077 & n4119 ) | ( n4098 & n4119 ) ;
  assign n4121 = ( n4077 & n4098 ) | ( n4077 & n4119 ) | ( n4098 & n4119 ) ;
  assign n4122 = ( n4077 & n4120 ) | ( n4077 & ~n4121 ) | ( n4120 & ~n4121 ) ;
  assign n4123 = ( n3959 & n3984 ) | ( n3959 & ~n4122 ) | ( n3984 & ~n4122 ) ;
  assign n4124 = ( n3959 & n3984 ) | ( n3959 & n4122 ) | ( n3984 & n4122 ) ;
  assign n4125 = ( n4122 & n4123 ) | ( n4122 & ~n4124 ) | ( n4123 & ~n4124 ) ;
  assign n4126 = x0 & x63 ;
  assign n4127 = ~x62 & n3947 ;
  assign n4128 = n4126 & n4127 ;
  assign n4129 = x1 & x62 ;
  assign n4130 = x32 & ~n4129 ;
  assign n4131 = x30 & x61 ;
  assign n4132 = x32 & ~n4131 ;
  assign n4133 = x32 | n4129 ;
  assign n4134 = ( n4130 & ~n4132 ) | ( n4130 & n4133 ) | ( ~n4132 & n4133 ) ;
  assign n4135 = ( n4126 & ~n4127 ) | ( n4126 & n4134 ) | ( ~n4127 & n4134 ) ;
  assign n4136 = n4126 & n4134 ;
  assign n4137 = ( n4128 & n4135 ) | ( n4128 & ~n4136 ) | ( n4135 & ~n4136 ) ;
  assign n4138 = x29 & x34 ;
  assign n4139 = x28 & x35 ;
  assign n4140 = x27 & x36 ;
  assign n4141 = ( ~n4138 & n4139 ) | ( ~n4138 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4142 = ( n4138 & n4139 ) | ( n4138 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4143 = ( n4138 & n4141 ) | ( n4138 & ~n4142 ) | ( n4141 & ~n4142 ) ;
  assign n4144 = x24 & x39 ;
  assign n4145 = x26 & x37 ;
  assign n4146 = x25 & x38 ;
  assign n4147 = ( ~n4144 & n4145 ) | ( ~n4144 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( n4144 & n4145 ) | ( n4144 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4149 = ( n4144 & n4147 ) | ( n4144 & ~n4148 ) | ( n4147 & ~n4148 ) ;
  assign n4150 = ( ~n4137 & n4143 ) | ( ~n4137 & n4149 ) | ( n4143 & n4149 ) ;
  assign n4151 = ( n4137 & n4143 ) | ( n4137 & n4149 ) | ( n4143 & n4149 ) ;
  assign n4152 = ( n4137 & n4150 ) | ( n4137 & ~n4151 ) | ( n4150 & ~n4151 ) ;
  assign n4153 = ( n3981 & n4005 ) | ( n3981 & n4152 ) | ( n4005 & n4152 ) ;
  assign n4154 = ( ~n3981 & n4005 ) | ( ~n3981 & n4152 ) | ( n4005 & n4152 ) ;
  assign n4155 = ( n3981 & ~n4153 ) | ( n3981 & n4154 ) | ( ~n4153 & n4154 ) ;
  assign n4156 = ( n3996 & ~n4011 ) | ( n3996 & n4017 ) | ( ~n4011 & n4017 ) ;
  assign n4157 = ( n3996 & n4011 ) | ( n3996 & n4017 ) | ( n4011 & n4017 ) ;
  assign n4158 = ( n4011 & n4156 ) | ( n4011 & ~n4157 ) | ( n4156 & ~n4157 ) ;
  assign n4159 = ( n4026 & n4047 ) | ( n4026 & n4158 ) | ( n4047 & n4158 ) ;
  assign n4160 = ( ~n4026 & n4047 ) | ( ~n4026 & n4158 ) | ( n4047 & n4158 ) ;
  assign n4161 = ( n4026 & ~n4159 ) | ( n4026 & n4160 ) | ( ~n4159 & n4160 ) ;
  assign n4162 = ( n3962 & n4155 ) | ( n3962 & n4161 ) | ( n4155 & n4161 ) ;
  assign n4163 = ( ~n3962 & n4155 ) | ( ~n3962 & n4161 ) | ( n4155 & n4161 ) ;
  assign n4164 = ( n3962 & ~n4162 ) | ( n3962 & n4163 ) | ( ~n4162 & n4163 ) ;
  assign n4165 = ( n3965 & n4125 ) | ( n3965 & n4164 ) | ( n4125 & n4164 ) ;
  assign n4166 = ( n3965 & ~n4125 ) | ( n3965 & n4164 ) | ( ~n4125 & n4164 ) ;
  assign n4167 = ( n4125 & ~n4165 ) | ( n4125 & n4166 ) | ( ~n4165 & n4166 ) ;
  assign n4168 = ( ~n4023 & n4038 ) | ( ~n4023 & n4044 ) | ( n4038 & n4044 ) ;
  assign n4169 = ( n4023 & n4038 ) | ( n4023 & n4044 ) | ( n4038 & n4044 ) ;
  assign n4170 = ( n4023 & n4168 ) | ( n4023 & ~n4169 ) | ( n4168 & ~n4169 ) ;
  assign n4171 = ( x2 & n1098 ) | ( x2 & n3987 ) | ( n1098 & n3987 ) ;
  assign n4172 = x60 & n4171 ;
  assign n4173 = ( n3972 & n4002 ) | ( n3972 & n4172 ) | ( n4002 & n4172 ) ;
  assign n4174 = ( n3972 & n4002 ) | ( n3972 & ~n4172 ) | ( n4002 & ~n4172 ) ;
  assign n4175 = ( n4172 & ~n4173 ) | ( n4172 & n4174 ) | ( ~n4173 & n4174 ) ;
  assign n4176 = ( n3954 & n4170 ) | ( n3954 & n4175 ) | ( n4170 & n4175 ) ;
  assign n4177 = ( n3954 & ~n4170 ) | ( n3954 & n4175 ) | ( ~n4170 & n4175 ) ;
  assign n4178 = ( n4170 & ~n4176 ) | ( n4170 & n4177 ) | ( ~n4176 & n4177 ) ;
  assign n4179 = ( n3943 & n3951 ) | ( n3943 & ~n3975 ) | ( n3951 & ~n3975 ) ;
  assign n4180 = ( n3943 & n3951 ) | ( n3943 & n3975 ) | ( n3951 & n3975 ) ;
  assign n4181 = ( n3975 & n4179 ) | ( n3975 & ~n4180 ) | ( n4179 & ~n4180 ) ;
  assign n4182 = ( n4050 & n4178 ) | ( n4050 & n4181 ) | ( n4178 & n4181 ) ;
  assign n4183 = ( ~n4050 & n4178 ) | ( ~n4050 & n4181 ) | ( n4178 & n4181 ) ;
  assign n4184 = ( n4050 & ~n4182 ) | ( n4050 & n4183 ) | ( ~n4182 & n4183 ) ;
  assign n4185 = ( n3940 & n3956 ) | ( n3940 & ~n3977 ) | ( n3956 & ~n3977 ) ;
  assign n4186 = ( n3940 & n3956 ) | ( n3940 & n3977 ) | ( n3956 & n3977 ) ;
  assign n4187 = ( n3977 & n4185 ) | ( n3977 & ~n4186 ) | ( n4185 & ~n4186 ) ;
  assign n4188 = ( n4053 & ~n4184 ) | ( n4053 & n4187 ) | ( ~n4184 & n4187 ) ;
  assign n4189 = ( n4053 & n4184 ) | ( n4053 & n4187 ) | ( n4184 & n4187 ) ;
  assign n4190 = ( n4184 & n4188 ) | ( n4184 & ~n4189 ) | ( n4188 & ~n4189 ) ;
  assign n4191 = ( ~n4056 & n4167 ) | ( ~n4056 & n4190 ) | ( n4167 & n4190 ) ;
  assign n4192 = ( n4056 & n4167 ) | ( n4056 & n4190 ) | ( n4167 & n4190 ) ;
  assign n4193 = ( n4056 & n4191 ) | ( n4056 & ~n4192 ) | ( n4191 & ~n4192 ) ;
  assign n4194 = ( n4058 & n4061 ) | ( n4058 & n4193 ) | ( n4061 & n4193 ) ;
  assign n4195 = ( n4058 & ~n4061 ) | ( n4058 & n4193 ) | ( ~n4061 & n4193 ) ;
  assign n4196 = ( n4061 & ~n4194 ) | ( n4061 & n4195 ) | ( ~n4194 & n4195 ) ;
  assign n4197 = x32 & x62 ;
  assign n4198 = ( ~x1 & x63 ) | ( ~x1 & n4197 ) | ( x63 & n4197 ) ;
  assign n4199 = ( x1 & x63 ) | ( x1 & n4197 ) | ( x63 & n4197 ) ;
  assign n4200 = ~n4198 & n4199 ;
  assign n4201 = n4082 & n4200 ;
  assign n4202 = n4082 | n4200 ;
  assign n4203 = ~n4201 & n4202 ;
  assign n4204 = x10 & x54 ;
  assign n4205 = x15 & x49 ;
  assign n4206 = x9 & x55 ;
  assign n4207 = ( ~n4204 & n4205 ) | ( ~n4204 & n4206 ) | ( n4205 & n4206 ) ;
  assign n4208 = ( n4204 & n4205 ) | ( n4204 & n4206 ) | ( n4205 & n4206 ) ;
  assign n4209 = ( n4204 & n4207 ) | ( n4204 & ~n4208 ) | ( n4207 & ~n4208 ) ;
  assign n4210 = x13 & x51 ;
  assign n4211 = x11 & x53 ;
  assign n4212 = x12 & x52 ;
  assign n4213 = ( ~n4210 & n4211 ) | ( ~n4210 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4214 = ( n4210 & n4211 ) | ( n4210 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4215 = ( n4210 & n4213 ) | ( n4210 & ~n4214 ) | ( n4213 & ~n4214 ) ;
  assign n4216 = ( n4203 & n4209 ) | ( n4203 & n4215 ) | ( n4209 & n4215 ) ;
  assign n4217 = ( ~n4203 & n4209 ) | ( ~n4203 & n4215 ) | ( n4209 & n4215 ) ;
  assign n4218 = ( n4203 & ~n4216 ) | ( n4203 & n4217 ) | ( ~n4216 & n4217 ) ;
  assign n4219 = ( n4076 & n4180 ) | ( n4076 & ~n4218 ) | ( n4180 & ~n4218 ) ;
  assign n4220 = ( n4076 & n4180 ) | ( n4076 & n4218 ) | ( n4180 & n4218 ) ;
  assign n4221 = ( n4218 & n4219 ) | ( n4218 & ~n4220 ) | ( n4219 & ~n4220 ) ;
  assign n4222 = ( n4109 & n4115 ) | ( n4109 & ~n4148 ) | ( n4115 & ~n4148 ) ;
  assign n4223 = ( n4109 & n4115 ) | ( n4109 & n4148 ) | ( n4115 & n4148 ) ;
  assign n4224 = ( n4148 & n4222 ) | ( n4148 & ~n4223 ) | ( n4222 & ~n4223 ) ;
  assign n4225 = ( n4097 & n4118 ) | ( n4097 & n4224 ) | ( n4118 & n4224 ) ;
  assign n4226 = ( n4097 & n4118 ) | ( n4097 & ~n4224 ) | ( n4118 & ~n4224 ) ;
  assign n4227 = ( n4224 & ~n4225 ) | ( n4224 & n4226 ) | ( ~n4225 & n4226 ) ;
  assign n4228 = ( n4186 & n4221 ) | ( n4186 & n4227 ) | ( n4221 & n4227 ) ;
  assign n4229 = ( ~n4186 & n4221 ) | ( ~n4186 & n4227 ) | ( n4221 & n4227 ) ;
  assign n4230 = ( n4186 & ~n4228 ) | ( n4186 & n4229 ) | ( ~n4228 & n4229 ) ;
  assign n4231 = x22 & x42 ;
  assign n4232 = x21 & x43 ;
  assign n4233 = x20 & x44 ;
  assign n4234 = ( ~n4231 & n4232 ) | ( ~n4231 & n4233 ) | ( n4232 & n4233 ) ;
  assign n4235 = ( n4231 & n4232 ) | ( n4231 & n4233 ) | ( n4232 & n4233 ) ;
  assign n4236 = ( n4231 & n4234 ) | ( n4231 & ~n4235 ) | ( n4234 & ~n4235 ) ;
  assign n4237 = x7 & x57 ;
  assign n4238 = x17 & x47 ;
  assign n4239 = x6 & x58 ;
  assign n4240 = ( ~n4237 & n4238 ) | ( ~n4237 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4241 = ( n4237 & n4238 ) | ( n4237 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4242 = ( n4237 & n4240 ) | ( n4237 & ~n4241 ) | ( n4240 & ~n4241 ) ;
  assign n4243 = x24 & x40 ;
  assign n4244 = x23 & x41 ;
  assign n4245 = x25 & x39 ;
  assign n4246 = ( ~n4243 & n4244 ) | ( ~n4243 & n4245 ) | ( n4244 & n4245 ) ;
  assign n4247 = ( n4243 & n4244 ) | ( n4243 & n4245 ) | ( n4244 & n4245 ) ;
  assign n4248 = ( n4243 & n4246 ) | ( n4243 & ~n4247 ) | ( n4246 & ~n4247 ) ;
  assign n4249 = ( ~n4236 & n4242 ) | ( ~n4236 & n4248 ) | ( n4242 & n4248 ) ;
  assign n4250 = ( n4236 & n4242 ) | ( n4236 & n4248 ) | ( n4242 & n4248 ) ;
  assign n4251 = ( n4236 & n4249 ) | ( n4236 & ~n4250 ) | ( n4249 & ~n4250 ) ;
  assign n4252 = n4127 | n4136 ;
  assign n4253 = x18 & x46 ;
  assign n4254 = x5 & x59 ;
  assign n4255 = x19 & x45 ;
  assign n4256 = ( ~n4253 & n4254 ) | ( ~n4253 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4257 = ( n4253 & n4254 ) | ( n4253 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4258 = ( n4253 & n4256 ) | ( n4253 & ~n4257 ) | ( n4256 & ~n4257 ) ;
  assign n4259 = x3 & x61 ;
  assign n4260 = x2 & x62 ;
  assign n4261 = x4 & x60 ;
  assign n4262 = ( ~n4259 & n4260 ) | ( ~n4259 & n4261 ) | ( n4260 & n4261 ) ;
  assign n4263 = ( n4259 & n4260 ) | ( n4259 & n4261 ) | ( n4260 & n4261 ) ;
  assign n4264 = ( n4259 & n4262 ) | ( n4259 & ~n4263 ) | ( n4262 & ~n4263 ) ;
  assign n4265 = ( n4252 & n4258 ) | ( n4252 & n4264 ) | ( n4258 & n4264 ) ;
  assign n4266 = ( ~n4252 & n4258 ) | ( ~n4252 & n4264 ) | ( n4258 & n4264 ) ;
  assign n4267 = ( n4252 & ~n4265 ) | ( n4252 & n4266 ) | ( ~n4265 & n4266 ) ;
  assign n4268 = x26 & x38 ;
  assign n4269 = x16 & x48 ;
  assign n4270 = x8 & x56 ;
  assign n4271 = ( ~n4268 & n4269 ) | ( ~n4268 & n4270 ) | ( n4269 & n4270 ) ;
  assign n4272 = ( n4268 & n4269 ) | ( n4268 & n4270 ) | ( n4269 & n4270 ) ;
  assign n4273 = ( n4268 & n4271 ) | ( n4268 & ~n4272 ) | ( n4271 & ~n4272 ) ;
  assign n4274 = x27 & x37 ;
  assign n4275 = x28 & x36 ;
  assign n4276 = x29 & x35 ;
  assign n4277 = ( ~n4274 & n4275 ) | ( ~n4274 & n4276 ) | ( n4275 & n4276 ) ;
  assign n4278 = ( n4274 & n4275 ) | ( n4274 & n4276 ) | ( n4275 & n4276 ) ;
  assign n4279 = ( n4274 & n4277 ) | ( n4274 & ~n4278 ) | ( n4277 & ~n4278 ) ;
  assign n4280 = x31 & x33 ;
  assign n4281 = x14 & x50 ;
  assign n4282 = x30 & x34 ;
  assign n4283 = ( ~n4280 & n4281 ) | ( ~n4280 & n4282 ) | ( n4281 & n4282 ) ;
  assign n4284 = ( n4280 & n4281 ) | ( n4280 & n4282 ) | ( n4281 & n4282 ) ;
  assign n4285 = ( n4280 & n4283 ) | ( n4280 & ~n4284 ) | ( n4283 & ~n4284 ) ;
  assign n4286 = ( ~n4273 & n4279 ) | ( ~n4273 & n4285 ) | ( n4279 & n4285 ) ;
  assign n4287 = ( n4273 & n4279 ) | ( n4273 & n4285 ) | ( n4279 & n4285 ) ;
  assign n4288 = ( n4273 & n4286 ) | ( n4273 & ~n4287 ) | ( n4286 & ~n4287 ) ;
  assign n4289 = ( ~n4251 & n4267 ) | ( ~n4251 & n4288 ) | ( n4267 & n4288 ) ;
  assign n4290 = ( n4251 & n4267 ) | ( n4251 & n4288 ) | ( n4267 & n4288 ) ;
  assign n4291 = ( n4251 & n4289 ) | ( n4251 & ~n4290 ) | ( n4289 & ~n4290 ) ;
  assign n4292 = ( n4157 & ~n4169 ) | ( n4157 & n4173 ) | ( ~n4169 & n4173 ) ;
  assign n4293 = ( n4157 & n4169 ) | ( n4157 & n4173 ) | ( n4169 & n4173 ) ;
  assign n4294 = ( n4169 & n4292 ) | ( n4169 & ~n4293 ) | ( n4292 & ~n4293 ) ;
  assign n4295 = ( n4159 & n4176 ) | ( n4159 & n4294 ) | ( n4176 & n4294 ) ;
  assign n4296 = ( n4159 & n4176 ) | ( n4159 & ~n4294 ) | ( n4176 & ~n4294 ) ;
  assign n4297 = ( n4294 & ~n4295 ) | ( n4294 & n4296 ) | ( ~n4295 & n4296 ) ;
  assign n4298 = ( n4182 & n4291 ) | ( n4182 & n4297 ) | ( n4291 & n4297 ) ;
  assign n4299 = ( ~n4182 & n4291 ) | ( ~n4182 & n4297 ) | ( n4291 & n4297 ) ;
  assign n4300 = ( n4182 & ~n4298 ) | ( n4182 & n4299 ) | ( ~n4298 & n4299 ) ;
  assign n4301 = ( n4189 & n4230 ) | ( n4189 & n4300 ) | ( n4230 & n4300 ) ;
  assign n4302 = ( ~n4189 & n4230 ) | ( ~n4189 & n4300 ) | ( n4230 & n4300 ) ;
  assign n4303 = ( n4189 & ~n4301 ) | ( n4189 & n4302 ) | ( ~n4301 & n4302 ) ;
  assign n4304 = ( n4088 & n4103 ) | ( n4088 & ~n4142 ) | ( n4103 & ~n4142 ) ;
  assign n4305 = ( n4088 & n4103 ) | ( n4088 & n4142 ) | ( n4103 & n4142 ) ;
  assign n4306 = ( n4142 & n4304 ) | ( n4142 & ~n4305 ) | ( n4304 & ~n4305 ) ;
  assign n4307 = ( n4068 & n4073 ) | ( n4068 & ~n4094 ) | ( n4073 & ~n4094 ) ;
  assign n4308 = ( n4068 & n4073 ) | ( n4068 & n4094 ) | ( n4073 & n4094 ) ;
  assign n4309 = ( n4094 & n4307 ) | ( n4094 & ~n4308 ) | ( n4307 & ~n4308 ) ;
  assign n4310 = ( ~n4151 & n4306 ) | ( ~n4151 & n4309 ) | ( n4306 & n4309 ) ;
  assign n4311 = ( n4151 & n4306 ) | ( n4151 & n4309 ) | ( n4306 & n4309 ) ;
  assign n4312 = ( n4151 & n4310 ) | ( n4151 & ~n4311 ) | ( n4310 & ~n4311 ) ;
  assign n4313 = ( n4121 & n4153 ) | ( n4121 & n4312 ) | ( n4153 & n4312 ) ;
  assign n4314 = ( n4121 & ~n4153 ) | ( n4121 & n4312 ) | ( ~n4153 & n4312 ) ;
  assign n4315 = ( n4153 & ~n4313 ) | ( n4153 & n4314 ) | ( ~n4313 & n4314 ) ;
  assign n4316 = ( n4124 & n4162 ) | ( n4124 & n4315 ) | ( n4162 & n4315 ) ;
  assign n4317 = ( ~n4124 & n4162 ) | ( ~n4124 & n4315 ) | ( n4162 & n4315 ) ;
  assign n4318 = ( n4124 & ~n4316 ) | ( n4124 & n4317 ) | ( ~n4316 & n4317 ) ;
  assign n4319 = ( n4165 & ~n4303 ) | ( n4165 & n4318 ) | ( ~n4303 & n4318 ) ;
  assign n4320 = ( n4165 & n4303 ) | ( n4165 & n4318 ) | ( n4303 & n4318 ) ;
  assign n4321 = ( n4303 & n4319 ) | ( n4303 & ~n4320 ) | ( n4319 & ~n4320 ) ;
  assign n4322 = ( n4192 & n4194 ) | ( n4192 & n4321 ) | ( n4194 & n4321 ) ;
  assign n4323 = ( n4192 & ~n4194 ) | ( n4192 & n4321 ) | ( ~n4194 & n4321 ) ;
  assign n4324 = ( n4194 & ~n4322 ) | ( n4194 & n4323 ) | ( ~n4322 & n4323 ) ;
  assign n4325 = x32 & x63 ;
  assign n4326 = n4129 & n4325 ;
  assign n4327 = n4201 | n4326 ;
  assign n4328 = x8 & x57 ;
  assign n4329 = x22 & x43 ;
  assign n4330 = x21 & x44 ;
  assign n4331 = ( ~n4328 & n4329 ) | ( ~n4328 & n4330 ) | ( n4329 & n4330 ) ;
  assign n4332 = ( n4328 & n4329 ) | ( n4328 & n4330 ) | ( n4329 & n4330 ) ;
  assign n4333 = ( n4328 & n4331 ) | ( n4328 & ~n4332 ) | ( n4331 & ~n4332 ) ;
  assign n4334 = x5 & x60 ;
  assign n4335 = x7 & x58 ;
  assign n4336 = x6 & x59 ;
  assign n4337 = ( ~n4334 & n4335 ) | ( ~n4334 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4338 = ( n4334 & n4335 ) | ( n4334 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4339 = ( n4334 & n4337 ) | ( n4334 & ~n4338 ) | ( n4337 & ~n4338 ) ;
  assign n4340 = ( ~n4327 & n4333 ) | ( ~n4327 & n4339 ) | ( n4333 & n4339 ) ;
  assign n4341 = ( n4327 & n4333 ) | ( n4327 & n4339 ) | ( n4333 & n4339 ) ;
  assign n4342 = ( n4327 & n4340 ) | ( n4327 & ~n4341 ) | ( n4340 & ~n4341 ) ;
  assign n4343 = x17 & x48 ;
  assign n4344 = x3 & x62 ;
  assign n4345 = ( ~x33 & n4343 ) | ( ~x33 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = ( x33 & n4343 ) | ( x33 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4347 = ( x33 & n4345 ) | ( x33 & ~n4346 ) | ( n4345 & ~n4346 ) ;
  assign n4348 = x11 & x54 ;
  assign n4349 = x19 & x46 ;
  assign n4350 = x29 & x36 ;
  assign n4351 = ( ~n4348 & n4349 ) | ( ~n4348 & n4350 ) | ( n4349 & n4350 ) ;
  assign n4352 = ( n4348 & n4349 ) | ( n4348 & n4350 ) | ( n4349 & n4350 ) ;
  assign n4353 = ( n4348 & n4351 ) | ( n4348 & ~n4352 ) | ( n4351 & ~n4352 ) ;
  assign n4354 = x31 & x34 ;
  assign n4355 = x32 & x33 ;
  assign n4356 = x30 & x35 ;
  assign n4357 = ( ~n4354 & n4355 ) | ( ~n4354 & n4356 ) | ( n4355 & n4356 ) ;
  assign n4358 = ( n4354 & n4355 ) | ( n4354 & n4356 ) | ( n4355 & n4356 ) ;
  assign n4359 = ( n4354 & n4357 ) | ( n4354 & ~n4358 ) | ( n4357 & ~n4358 ) ;
  assign n4360 = ( ~n4347 & n4353 ) | ( ~n4347 & n4359 ) | ( n4353 & n4359 ) ;
  assign n4361 = ( n4347 & n4353 ) | ( n4347 & n4359 ) | ( n4353 & n4359 ) ;
  assign n4362 = ( n4347 & n4360 ) | ( n4347 & ~n4361 ) | ( n4360 & ~n4361 ) ;
  assign n4363 = x23 & x42 ;
  assign n4364 = x25 & x40 ;
  assign n4365 = x24 & x41 ;
  assign n4366 = ( ~n4363 & n4364 ) | ( ~n4363 & n4365 ) | ( n4364 & n4365 ) ;
  assign n4367 = ( n4363 & n4364 ) | ( n4363 & n4365 ) | ( n4364 & n4365 ) ;
  assign n4368 = ( n4363 & n4366 ) | ( n4363 & ~n4367 ) | ( n4366 & ~n4367 ) ;
  assign n4369 = x9 & x56 ;
  assign n4370 = x10 & x55 ;
  assign n4371 = x20 & x45 ;
  assign n4372 = ( ~n4369 & n4370 ) | ( ~n4369 & n4371 ) | ( n4370 & n4371 ) ;
  assign n4373 = ( n4369 & n4370 ) | ( n4369 & n4371 ) | ( n4370 & n4371 ) ;
  assign n4374 = ( n4369 & n4372 ) | ( n4369 & ~n4373 ) | ( n4372 & ~n4373 ) ;
  assign n4375 = x27 & x38 ;
  assign n4376 = x28 & x37 ;
  assign n4377 = x26 & x39 ;
  assign n4378 = ( ~n4375 & n4376 ) | ( ~n4375 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4379 = ( n4375 & n4376 ) | ( n4375 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4380 = ( n4375 & n4378 ) | ( n4375 & ~n4379 ) | ( n4378 & ~n4379 ) ;
  assign n4381 = ( ~n4368 & n4374 ) | ( ~n4368 & n4380 ) | ( n4374 & n4380 ) ;
  assign n4382 = ( n4368 & n4374 ) | ( n4368 & n4380 ) | ( n4374 & n4380 ) ;
  assign n4383 = ( n4368 & n4381 ) | ( n4368 & ~n4382 ) | ( n4381 & ~n4382 ) ;
  assign n4384 = ( ~n4342 & n4362 ) | ( ~n4342 & n4383 ) | ( n4362 & n4383 ) ;
  assign n4385 = ( n4342 & n4362 ) | ( n4342 & n4383 ) | ( n4362 & n4383 ) ;
  assign n4386 = ( n4342 & n4384 ) | ( n4342 & ~n4385 ) | ( n4384 & ~n4385 ) ;
  assign n4387 = ( ~n4223 & n4305 ) | ( ~n4223 & n4308 ) | ( n4305 & n4308 ) ;
  assign n4388 = ( n4223 & n4305 ) | ( n4223 & n4308 ) | ( n4305 & n4308 ) ;
  assign n4389 = ( n4223 & n4387 ) | ( n4223 & ~n4388 ) | ( n4387 & ~n4388 ) ;
  assign n4390 = ( n4225 & n4311 ) | ( n4225 & ~n4389 ) | ( n4311 & ~n4389 ) ;
  assign n4391 = ( n4225 & n4311 ) | ( n4225 & n4389 ) | ( n4311 & n4389 ) ;
  assign n4392 = ( n4389 & n4390 ) | ( n4389 & ~n4391 ) | ( n4390 & ~n4391 ) ;
  assign n4393 = ( n4313 & n4386 ) | ( n4313 & n4392 ) | ( n4386 & n4392 ) ;
  assign n4394 = ( ~n4313 & n4386 ) | ( ~n4313 & n4392 ) | ( n4386 & n4392 ) ;
  assign n4395 = ( n4313 & ~n4393 ) | ( n4313 & n4394 ) | ( ~n4393 & n4394 ) ;
  assign n4396 = x4 & x61 ;
  assign n4397 = x2 & x63 ;
  assign n4398 = ( n4284 & n4396 ) | ( n4284 & n4397 ) | ( n4396 & n4397 ) ;
  assign n4399 = ( ~n4284 & n4396 ) | ( ~n4284 & n4397 ) | ( n4396 & n4397 ) ;
  assign n4400 = ( n4284 & ~n4398 ) | ( n4284 & n4399 ) | ( ~n4398 & n4399 ) ;
  assign n4401 = x16 & x49 ;
  assign n4402 = x15 & x50 ;
  assign n4403 = x14 & x51 ;
  assign n4404 = ( ~n4401 & n4402 ) | ( ~n4401 & n4403 ) | ( n4402 & n4403 ) ;
  assign n4405 = ( n4401 & n4402 ) | ( n4401 & n4403 ) | ( n4402 & n4403 ) ;
  assign n4406 = ( n4401 & n4404 ) | ( n4401 & ~n4405 ) | ( n4404 & ~n4405 ) ;
  assign n4407 = x12 & x53 ;
  assign n4408 = x13 & x52 ;
  assign n4409 = x18 & x47 ;
  assign n4410 = ( ~n4407 & n4408 ) | ( ~n4407 & n4409 ) | ( n4408 & n4409 ) ;
  assign n4411 = ( n4407 & n4408 ) | ( n4407 & n4409 ) | ( n4408 & n4409 ) ;
  assign n4412 = ( n4407 & n4410 ) | ( n4407 & ~n4411 ) | ( n4410 & ~n4411 ) ;
  assign n4413 = ( n4400 & n4406 ) | ( n4400 & n4412 ) | ( n4406 & n4412 ) ;
  assign n4414 = ( ~n4400 & n4406 ) | ( ~n4400 & n4412 ) | ( n4406 & n4412 ) ;
  assign n4415 = ( n4400 & ~n4413 ) | ( n4400 & n4414 ) | ( ~n4413 & n4414 ) ;
  assign n4416 = ( n4265 & n4293 ) | ( n4265 & ~n4415 ) | ( n4293 & ~n4415 ) ;
  assign n4417 = ( n4265 & n4293 ) | ( n4265 & n4415 ) | ( n4293 & n4415 ) ;
  assign n4418 = ( n4415 & n4416 ) | ( n4415 & ~n4417 ) | ( n4416 & ~n4417 ) ;
  assign n4419 = ( n4214 & ~n4235 ) | ( n4214 & n4278 ) | ( ~n4235 & n4278 ) ;
  assign n4420 = ( n4214 & n4235 ) | ( n4214 & n4278 ) | ( n4235 & n4278 ) ;
  assign n4421 = ( n4235 & n4419 ) | ( n4235 & ~n4420 ) | ( n4419 & ~n4420 ) ;
  assign n4422 = ( n4250 & n4287 ) | ( n4250 & n4421 ) | ( n4287 & n4421 ) ;
  assign n4423 = ( n4250 & n4287 ) | ( n4250 & ~n4421 ) | ( n4287 & ~n4421 ) ;
  assign n4424 = ( n4421 & ~n4422 ) | ( n4421 & n4423 ) | ( ~n4422 & n4423 ) ;
  assign n4425 = ( n4295 & n4418 ) | ( n4295 & n4424 ) | ( n4418 & n4424 ) ;
  assign n4426 = ( n4295 & ~n4418 ) | ( n4295 & n4424 ) | ( ~n4418 & n4424 ) ;
  assign n4427 = ( n4418 & ~n4425 ) | ( n4418 & n4426 ) | ( ~n4425 & n4426 ) ;
  assign n4428 = ( n4316 & ~n4395 ) | ( n4316 & n4427 ) | ( ~n4395 & n4427 ) ;
  assign n4429 = ( n4316 & n4395 ) | ( n4316 & n4427 ) | ( n4395 & n4427 ) ;
  assign n4430 = ( n4395 & n4428 ) | ( n4395 & ~n4429 ) | ( n4428 & ~n4429 ) ;
  assign n4431 = ( n4257 & n4263 ) | ( n4257 & ~n4272 ) | ( n4263 & ~n4272 ) ;
  assign n4432 = ( n4257 & n4263 ) | ( n4257 & n4272 ) | ( n4263 & n4272 ) ;
  assign n4433 = ( n4272 & n4431 ) | ( n4272 & ~n4432 ) | ( n4431 & ~n4432 ) ;
  assign n4434 = ( n4208 & ~n4241 ) | ( n4208 & n4247 ) | ( ~n4241 & n4247 ) ;
  assign n4435 = ( n4208 & n4241 ) | ( n4208 & n4247 ) | ( n4241 & n4247 ) ;
  assign n4436 = ( n4241 & n4434 ) | ( n4241 & ~n4435 ) | ( n4434 & ~n4435 ) ;
  assign n4437 = ( n4216 & n4433 ) | ( n4216 & n4436 ) | ( n4433 & n4436 ) ;
  assign n4438 = ( ~n4216 & n4433 ) | ( ~n4216 & n4436 ) | ( n4433 & n4436 ) ;
  assign n4439 = ( n4216 & ~n4437 ) | ( n4216 & n4438 ) | ( ~n4437 & n4438 ) ;
  assign n4440 = ( n4220 & n4290 ) | ( n4220 & n4439 ) | ( n4290 & n4439 ) ;
  assign n4441 = ( ~n4220 & n4290 ) | ( ~n4220 & n4439 ) | ( n4290 & n4439 ) ;
  assign n4442 = ( n4220 & ~n4440 ) | ( n4220 & n4441 ) | ( ~n4440 & n4441 ) ;
  assign n4443 = ( n4228 & n4298 ) | ( n4228 & n4442 ) | ( n4298 & n4442 ) ;
  assign n4444 = ( ~n4228 & n4298 ) | ( ~n4228 & n4442 ) | ( n4298 & n4442 ) ;
  assign n4445 = ( n4228 & ~n4443 ) | ( n4228 & n4444 ) | ( ~n4443 & n4444 ) ;
  assign n4446 = ( ~n4301 & n4430 ) | ( ~n4301 & n4445 ) | ( n4430 & n4445 ) ;
  assign n4447 = ( n4301 & n4430 ) | ( n4301 & n4445 ) | ( n4430 & n4445 ) ;
  assign n4448 = ( n4301 & n4446 ) | ( n4301 & ~n4447 ) | ( n4446 & ~n4447 ) ;
  assign n4449 = ( n4320 & ~n4322 ) | ( n4320 & n4448 ) | ( ~n4322 & n4448 ) ;
  assign n4450 = ( n4320 & n4322 ) | ( n4320 & n4448 ) | ( n4322 & n4448 ) ;
  assign n4451 = ( n4322 & n4449 ) | ( n4322 & ~n4450 ) | ( n4449 & ~n4450 ) ;
  assign n4452 = ( ~n4420 & n4432 ) | ( ~n4420 & n4435 ) | ( n4432 & n4435 ) ;
  assign n4453 = ( n4420 & n4432 ) | ( n4420 & n4435 ) | ( n4432 & n4435 ) ;
  assign n4454 = ( n4420 & n4452 ) | ( n4420 & ~n4453 ) | ( n4452 & ~n4453 ) ;
  assign n4455 = ( n4422 & n4437 ) | ( n4422 & ~n4454 ) | ( n4437 & ~n4454 ) ;
  assign n4456 = ( n4422 & n4437 ) | ( n4422 & n4454 ) | ( n4437 & n4454 ) ;
  assign n4457 = ( n4454 & n4455 ) | ( n4454 & ~n4456 ) | ( n4455 & ~n4456 ) ;
  assign n4458 = x29 & x37 ;
  assign n4459 = x28 & x38 ;
  assign n4460 = x27 & x39 ;
  assign n4461 = ( ~n4458 & n4459 ) | ( ~n4458 & n4460 ) | ( n4459 & n4460 ) ;
  assign n4462 = ( n4458 & n4459 ) | ( n4458 & n4460 ) | ( n4459 & n4460 ) ;
  assign n4463 = ( n4458 & n4461 ) | ( n4458 & ~n4462 ) | ( n4461 & ~n4462 ) ;
  assign n4464 = x3 & x63 ;
  assign n4465 = x4 & x62 ;
  assign n4466 = x5 & x61 ;
  assign n4467 = ( ~n4464 & n4465 ) | ( ~n4464 & n4466 ) | ( n4465 & n4466 ) ;
  assign n4468 = ( n4464 & n4465 ) | ( n4464 & n4466 ) | ( n4465 & n4466 ) ;
  assign n4469 = ( n4464 & n4467 ) | ( n4464 & ~n4468 ) | ( n4467 & ~n4468 ) ;
  assign n4470 = x19 & x47 ;
  assign n4471 = x11 & x55 ;
  assign n4472 = x12 & x54 ;
  assign n4473 = ( ~n4470 & n4471 ) | ( ~n4470 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4474 = ( n4470 & n4471 ) | ( n4470 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4475 = ( n4470 & n4473 ) | ( n4470 & ~n4474 ) | ( n4473 & ~n4474 ) ;
  assign n4476 = ( ~n4463 & n4469 ) | ( ~n4463 & n4475 ) | ( n4469 & n4475 ) ;
  assign n4477 = ( n4463 & n4469 ) | ( n4463 & n4475 ) | ( n4469 & n4475 ) ;
  assign n4478 = ( n4463 & n4476 ) | ( n4463 & ~n4477 ) | ( n4476 & ~n4477 ) ;
  assign n4479 = x32 & x34 ;
  assign n4480 = x17 & x49 ;
  assign n4481 = x16 & x50 ;
  assign n4482 = ( ~n4479 & n4480 ) | ( ~n4479 & n4481 ) | ( n4480 & n4481 ) ;
  assign n4483 = ( n4479 & n4480 ) | ( n4479 & n4481 ) | ( n4480 & n4481 ) ;
  assign n4484 = ( n4479 & n4482 ) | ( n4479 & ~n4483 ) | ( n4482 & ~n4483 ) ;
  assign n4485 = x30 & x36 ;
  assign n4486 = x31 & x35 ;
  assign n4487 = x14 & x52 ;
  assign n4488 = ( ~n4485 & n4486 ) | ( ~n4485 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4489 = ( n4485 & n4486 ) | ( n4485 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4490 = ( n4485 & n4488 ) | ( n4485 & ~n4489 ) | ( n4488 & ~n4489 ) ;
  assign n4491 = x15 & x51 ;
  assign n4492 = x18 & x48 ;
  assign n4493 = x13 & x53 ;
  assign n4494 = ( ~n4491 & n4492 ) | ( ~n4491 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4495 = ( n4491 & n4492 ) | ( n4491 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4496 = ( n4491 & n4494 ) | ( n4491 & ~n4495 ) | ( n4494 & ~n4495 ) ;
  assign n4497 = ( ~n4484 & n4490 ) | ( ~n4484 & n4496 ) | ( n4490 & n4496 ) ;
  assign n4498 = ( n4484 & n4490 ) | ( n4484 & n4496 ) | ( n4490 & n4496 ) ;
  assign n4499 = ( n4484 & n4497 ) | ( n4484 & ~n4498 ) | ( n4497 & ~n4498 ) ;
  assign n4500 = x26 & x40 ;
  assign n4501 = x25 & x41 ;
  assign n4502 = x10 & x56 ;
  assign n4503 = ( ~n4500 & n4501 ) | ( ~n4500 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4504 = ( n4500 & n4501 ) | ( n4500 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4505 = ( n4500 & n4503 ) | ( n4500 & ~n4504 ) | ( n4503 & ~n4504 ) ;
  assign n4506 = x22 & x44 ;
  assign n4507 = x21 & x45 ;
  assign n4508 = x20 & x46 ;
  assign n4509 = ( ~n4506 & n4507 ) | ( ~n4506 & n4508 ) | ( n4507 & n4508 ) ;
  assign n4510 = ( n4506 & n4507 ) | ( n4506 & n4508 ) | ( n4507 & n4508 ) ;
  assign n4511 = ( n4506 & n4509 ) | ( n4506 & ~n4510 ) | ( n4509 & ~n4510 ) ;
  assign n4512 = x9 & x57 ;
  assign n4513 = x24 & x42 ;
  assign n4514 = ( ~n2074 & n4512 ) | ( ~n2074 & n4513 ) | ( n4512 & n4513 ) ;
  assign n4515 = ( n2074 & n4512 ) | ( n2074 & n4513 ) | ( n4512 & n4513 ) ;
  assign n4516 = ( n2074 & n4514 ) | ( n2074 & ~n4515 ) | ( n4514 & ~n4515 ) ;
  assign n4517 = ( ~n4505 & n4511 ) | ( ~n4505 & n4516 ) | ( n4511 & n4516 ) ;
  assign n4518 = ( n4505 & n4511 ) | ( n4505 & n4516 ) | ( n4511 & n4516 ) ;
  assign n4519 = ( n4505 & n4517 ) | ( n4505 & ~n4518 ) | ( n4517 & ~n4518 ) ;
  assign n4520 = ( ~n4478 & n4499 ) | ( ~n4478 & n4519 ) | ( n4499 & n4519 ) ;
  assign n4521 = ( n4478 & n4499 ) | ( n4478 & n4519 ) | ( n4499 & n4519 ) ;
  assign n4522 = ( n4478 & n4520 ) | ( n4478 & ~n4521 ) | ( n4520 & ~n4521 ) ;
  assign n4523 = ( n4440 & n4457 ) | ( n4440 & n4522 ) | ( n4457 & n4522 ) ;
  assign n4524 = ( ~n4440 & n4457 ) | ( ~n4440 & n4522 ) | ( n4457 & n4522 ) ;
  assign n4525 = ( n4440 & ~n4523 ) | ( n4440 & n4524 ) | ( ~n4523 & n4524 ) ;
  assign n4526 = ( n4393 & ~n4443 ) | ( n4393 & n4525 ) | ( ~n4443 & n4525 ) ;
  assign n4527 = ( n4393 & n4443 ) | ( n4393 & n4525 ) | ( n4443 & n4525 ) ;
  assign n4528 = ( n4443 & n4526 ) | ( n4443 & ~n4527 ) | ( n4526 & ~n4527 ) ;
  assign n4529 = x7 & x59 ;
  assign n4530 = x6 & x60 ;
  assign n4531 = x8 & x58 ;
  assign n4532 = ( ~n4529 & n4530 ) | ( ~n4529 & n4531 ) | ( n4530 & n4531 ) ;
  assign n4533 = ( n4529 & n4530 ) | ( n4529 & n4531 ) | ( n4530 & n4531 ) ;
  assign n4534 = ( n4529 & n4532 ) | ( n4529 & ~n4533 ) | ( n4532 & ~n4533 ) ;
  assign n4535 = ( n4379 & ~n4398 ) | ( n4379 & n4534 ) | ( ~n4398 & n4534 ) ;
  assign n4536 = ( n4379 & n4398 ) | ( n4379 & n4534 ) | ( n4398 & n4534 ) ;
  assign n4537 = ( n4398 & n4535 ) | ( n4398 & ~n4536 ) | ( n4535 & ~n4536 ) ;
  assign n4538 = ( ~n4388 & n4413 ) | ( ~n4388 & n4537 ) | ( n4413 & n4537 ) ;
  assign n4539 = ( n4388 & n4413 ) | ( n4388 & n4537 ) | ( n4413 & n4537 ) ;
  assign n4540 = ( n4388 & n4538 ) | ( n4388 & ~n4539 ) | ( n4538 & ~n4539 ) ;
  assign n4541 = ( n4332 & n4338 ) | ( n4332 & ~n4352 ) | ( n4338 & ~n4352 ) ;
  assign n4542 = ( n4332 & n4338 ) | ( n4332 & n4352 ) | ( n4338 & n4352 ) ;
  assign n4543 = ( n4352 & n4541 ) | ( n4352 & ~n4542 ) | ( n4541 & ~n4542 ) ;
  assign n4544 = ( n4346 & n4358 ) | ( n4346 & ~n4405 ) | ( n4358 & ~n4405 ) ;
  assign n4545 = ( n4346 & n4358 ) | ( n4346 & n4405 ) | ( n4358 & n4405 ) ;
  assign n4546 = ( n4405 & n4544 ) | ( n4405 & ~n4545 ) | ( n4544 & ~n4545 ) ;
  assign n4547 = ( n4361 & n4543 ) | ( n4361 & n4546 ) | ( n4543 & n4546 ) ;
  assign n4548 = ( n4361 & ~n4543 ) | ( n4361 & n4546 ) | ( ~n4543 & n4546 ) ;
  assign n4549 = ( n4543 & ~n4547 ) | ( n4543 & n4548 ) | ( ~n4547 & n4548 ) ;
  assign n4550 = ( n4391 & n4540 ) | ( n4391 & n4549 ) | ( n4540 & n4549 ) ;
  assign n4551 = ( ~n4391 & n4540 ) | ( ~n4391 & n4549 ) | ( n4540 & n4549 ) ;
  assign n4552 = ( n4391 & ~n4550 ) | ( n4391 & n4551 ) | ( ~n4550 & n4551 ) ;
  assign n4553 = ( n4367 & n4373 ) | ( n4367 & ~n4411 ) | ( n4373 & ~n4411 ) ;
  assign n4554 = ( n4367 & n4373 ) | ( n4367 & n4411 ) | ( n4373 & n4411 ) ;
  assign n4555 = ( n4411 & n4553 ) | ( n4411 & ~n4554 ) | ( n4553 & ~n4554 ) ;
  assign n4556 = ( n4341 & n4382 ) | ( n4341 & n4555 ) | ( n4382 & n4555 ) ;
  assign n4557 = ( ~n4341 & n4382 ) | ( ~n4341 & n4555 ) | ( n4382 & n4555 ) ;
  assign n4558 = ( n4341 & ~n4556 ) | ( n4341 & n4557 ) | ( ~n4556 & n4557 ) ;
  assign n4559 = ( n4385 & n4417 ) | ( n4385 & n4558 ) | ( n4417 & n4558 ) ;
  assign n4560 = ( n4385 & n4417 ) | ( n4385 & ~n4558 ) | ( n4417 & ~n4558 ) ;
  assign n4561 = ( n4558 & ~n4559 ) | ( n4558 & n4560 ) | ( ~n4559 & n4560 ) ;
  assign n4562 = ( n4425 & n4552 ) | ( n4425 & n4561 ) | ( n4552 & n4561 ) ;
  assign n4563 = ( n4425 & ~n4552 ) | ( n4425 & n4561 ) | ( ~n4552 & n4561 ) ;
  assign n4564 = ( n4552 & ~n4562 ) | ( n4552 & n4563 ) | ( ~n4562 & n4563 ) ;
  assign n4565 = ( n4429 & n4528 ) | ( n4429 & n4564 ) | ( n4528 & n4564 ) ;
  assign n4566 = ( ~n4429 & n4528 ) | ( ~n4429 & n4564 ) | ( n4528 & n4564 ) ;
  assign n4567 = ( n4429 & ~n4565 ) | ( n4429 & n4566 ) | ( ~n4565 & n4566 ) ;
  assign n4568 = ( n4447 & ~n4450 ) | ( n4447 & n4567 ) | ( ~n4450 & n4567 ) ;
  assign n4569 = ( n4447 & n4450 ) | ( n4447 & n4567 ) | ( n4450 & n4567 ) ;
  assign n4570 = ( n4450 & n4568 ) | ( n4450 & ~n4569 ) | ( n4568 & ~n4569 ) ;
  assign n4571 = ( n4542 & n4545 ) | ( n4542 & n4554 ) | ( n4545 & n4554 ) ;
  assign n4572 = ( n4542 & n4545 ) | ( n4542 & ~n4554 ) | ( n4545 & ~n4554 ) ;
  assign n4573 = ( n4554 & ~n4571 ) | ( n4554 & n4572 ) | ( ~n4571 & n4572 ) ;
  assign n4574 = ( n4547 & n4556 ) | ( n4547 & n4573 ) | ( n4556 & n4573 ) ;
  assign n4575 = ( n4547 & n4556 ) | ( n4547 & ~n4573 ) | ( n4556 & ~n4573 ) ;
  assign n4576 = ( n4573 & ~n4574 ) | ( n4573 & n4575 ) | ( ~n4574 & n4575 ) ;
  assign n4577 = x4 & x63 ;
  assign n4578 = x28 & x39 ;
  assign n4579 = x27 & x40 ;
  assign n4580 = ( ~n4577 & n4578 ) | ( ~n4577 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4581 = ( n4577 & n4578 ) | ( n4577 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4582 = ( n4577 & n4580 ) | ( n4577 & ~n4581 ) | ( n4580 & ~n4581 ) ;
  assign n4583 = x21 & x46 ;
  assign n4584 = x26 & x41 ;
  assign n4585 = x25 & x42 ;
  assign n4586 = ( ~n4583 & n4584 ) | ( ~n4583 & n4585 ) | ( n4584 & n4585 ) ;
  assign n4587 = ( n4583 & n4584 ) | ( n4583 & n4585 ) | ( n4584 & n4585 ) ;
  assign n4588 = ( n4583 & n4586 ) | ( n4583 & ~n4587 ) | ( n4586 & ~n4587 ) ;
  assign n4589 = x17 & x50 ;
  assign n4590 = x19 & x48 ;
  assign n4591 = x14 & x53 ;
  assign n4592 = ( ~n4589 & n4590 ) | ( ~n4589 & n4591 ) | ( n4590 & n4591 ) ;
  assign n4593 = ( n4589 & n4590 ) | ( n4589 & n4591 ) | ( n4590 & n4591 ) ;
  assign n4594 = ( n4589 & n4592 ) | ( n4589 & ~n4593 ) | ( n4592 & ~n4593 ) ;
  assign n4595 = ( ~n4582 & n4588 ) | ( ~n4582 & n4594 ) | ( n4588 & n4594 ) ;
  assign n4596 = ( n4582 & n4588 ) | ( n4582 & n4594 ) | ( n4588 & n4594 ) ;
  assign n4597 = ( n4582 & n4595 ) | ( n4582 & ~n4596 ) | ( n4595 & ~n4596 ) ;
  assign n4598 = x24 & x43 ;
  assign n4599 = x23 & x44 ;
  assign n4600 = x22 & x45 ;
  assign n4601 = ( ~n4598 & n4599 ) | ( ~n4598 & n4600 ) | ( n4599 & n4600 ) ;
  assign n4602 = ( n4598 & n4599 ) | ( n4598 & n4600 ) | ( n4599 & n4600 ) ;
  assign n4603 = ( n4598 & n4601 ) | ( n4598 & ~n4602 ) | ( n4601 & ~n4602 ) ;
  assign n4604 = x15 & x52 ;
  assign n4605 = x16 & x51 ;
  assign n4606 = x30 & x37 ;
  assign n4607 = ( ~n4604 & n4605 ) | ( ~n4604 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4608 = ( n4604 & n4605 ) | ( n4604 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4609 = ( n4604 & n4607 ) | ( n4604 & ~n4608 ) | ( n4607 & ~n4608 ) ;
  assign n4610 = x8 & x59 ;
  assign n4611 = x7 & x60 ;
  assign n4612 = x9 & x58 ;
  assign n4613 = ( ~n4610 & n4611 ) | ( ~n4610 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4614 = ( n4610 & n4611 ) | ( n4610 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4615 = ( n4610 & n4613 ) | ( n4610 & ~n4614 ) | ( n4613 & ~n4614 ) ;
  assign n4616 = ( ~n4603 & n4609 ) | ( ~n4603 & n4615 ) | ( n4609 & n4615 ) ;
  assign n4617 = ( n4603 & n4609 ) | ( n4603 & n4615 ) | ( n4609 & n4615 ) ;
  assign n4618 = ( n4603 & n4616 ) | ( n4603 & ~n4617 ) | ( n4616 & ~n4617 ) ;
  assign n4619 = x18 & x49 ;
  assign n4620 = x5 & x62 ;
  assign n4621 = ( ~x34 & n4619 ) | ( ~x34 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4622 = ( x34 & n4619 ) | ( x34 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4623 = ( x34 & n4621 ) | ( x34 & ~n4622 ) | ( n4621 & ~n4622 ) ;
  assign n4624 = x32 & x35 ;
  assign n4625 = x33 & x34 ;
  assign n4626 = x31 & x36 ;
  assign n4627 = ( ~n4624 & n4625 ) | ( ~n4624 & n4626 ) | ( n4625 & n4626 ) ;
  assign n4628 = ( n4624 & n4625 ) | ( n4624 & n4626 ) | ( n4625 & n4626 ) ;
  assign n4629 = ( n4624 & n4627 ) | ( n4624 & ~n4628 ) | ( n4627 & ~n4628 ) ;
  assign n4630 = x12 & x55 ;
  assign n4631 = x13 & x54 ;
  assign n4632 = x29 & x38 ;
  assign n4633 = ( ~n4630 & n4631 ) | ( ~n4630 & n4632 ) | ( n4631 & n4632 ) ;
  assign n4634 = ( n4630 & n4631 ) | ( n4630 & n4632 ) | ( n4631 & n4632 ) ;
  assign n4635 = ( n4630 & n4633 ) | ( n4630 & ~n4634 ) | ( n4633 & ~n4634 ) ;
  assign n4636 = ( ~n4623 & n4629 ) | ( ~n4623 & n4635 ) | ( n4629 & n4635 ) ;
  assign n4637 = ( n4623 & n4629 ) | ( n4623 & n4635 ) | ( n4629 & n4635 ) ;
  assign n4638 = ( n4623 & n4636 ) | ( n4623 & ~n4637 ) | ( n4636 & ~n4637 ) ;
  assign n4639 = ( ~n4597 & n4618 ) | ( ~n4597 & n4638 ) | ( n4618 & n4638 ) ;
  assign n4640 = ( n4597 & n4618 ) | ( n4597 & n4638 ) | ( n4618 & n4638 ) ;
  assign n4641 = ( n4597 & n4639 ) | ( n4597 & ~n4640 ) | ( n4639 & ~n4640 ) ;
  assign n4642 = ( n4559 & n4576 ) | ( n4559 & n4641 ) | ( n4576 & n4641 ) ;
  assign n4643 = ( ~n4559 & n4576 ) | ( ~n4559 & n4641 ) | ( n4576 & n4641 ) ;
  assign n4644 = ( n4559 & ~n4642 ) | ( n4559 & n4643 ) | ( ~n4642 & n4643 ) ;
  assign n4645 = ( n4523 & n4562 ) | ( n4523 & n4644 ) | ( n4562 & n4644 ) ;
  assign n4646 = ( n4523 & ~n4562 ) | ( n4523 & n4644 ) | ( ~n4562 & n4644 ) ;
  assign n4647 = ( n4562 & ~n4645 ) | ( n4562 & n4646 ) | ( ~n4645 & n4646 ) ;
  assign n4648 = ( n4462 & n4468 ) | ( n4462 & ~n4533 ) | ( n4468 & ~n4533 ) ;
  assign n4649 = ( n4462 & n4468 ) | ( n4462 & n4533 ) | ( n4468 & n4533 ) ;
  assign n4650 = ( n4533 & n4648 ) | ( n4533 & ~n4649 ) | ( n4648 & ~n4649 ) ;
  assign n4651 = ( ~n4504 & n4510 ) | ( ~n4504 & n4515 ) | ( n4510 & n4515 ) ;
  assign n4652 = ( n4504 & n4510 ) | ( n4504 & n4515 ) | ( n4510 & n4515 ) ;
  assign n4653 = ( n4504 & n4651 ) | ( n4504 & ~n4652 ) | ( n4651 & ~n4652 ) ;
  assign n4654 = x6 & x61 ;
  assign n4655 = ( n4483 & n4489 ) | ( n4483 & n4654 ) | ( n4489 & n4654 ) ;
  assign n4656 = ( ~n4483 & n4489 ) | ( ~n4483 & n4654 ) | ( n4489 & n4654 ) ;
  assign n4657 = ( n4483 & ~n4655 ) | ( n4483 & n4656 ) | ( ~n4655 & n4656 ) ;
  assign n4658 = ( ~n4650 & n4653 ) | ( ~n4650 & n4657 ) | ( n4653 & n4657 ) ;
  assign n4659 = ( n4650 & n4653 ) | ( n4650 & n4657 ) | ( n4653 & n4657 ) ;
  assign n4660 = ( n4650 & n4658 ) | ( n4650 & ~n4659 ) | ( n4658 & ~n4659 ) ;
  assign n4661 = ( n4477 & n4518 ) | ( n4477 & ~n4536 ) | ( n4518 & ~n4536 ) ;
  assign n4662 = ( n4477 & n4518 ) | ( n4477 & n4536 ) | ( n4518 & n4536 ) ;
  assign n4663 = ( n4536 & n4661 ) | ( n4536 & ~n4662 ) | ( n4661 & ~n4662 ) ;
  assign n4664 = ( n4456 & n4660 ) | ( n4456 & n4663 ) | ( n4660 & n4663 ) ;
  assign n4665 = ( ~n4456 & n4660 ) | ( ~n4456 & n4663 ) | ( n4660 & n4663 ) ;
  assign n4666 = ( n4456 & ~n4664 ) | ( n4456 & n4665 ) | ( ~n4664 & n4665 ) ;
  assign n4667 = x20 & x47 ;
  assign n4668 = x10 & x57 ;
  assign n4669 = x11 & x56 ;
  assign n4670 = ( ~n4667 & n4668 ) | ( ~n4667 & n4669 ) | ( n4668 & n4669 ) ;
  assign n4671 = ( n4667 & n4668 ) | ( n4667 & n4669 ) | ( n4668 & n4669 ) ;
  assign n4672 = ( n4667 & n4670 ) | ( n4667 & ~n4671 ) | ( n4670 & ~n4671 ) ;
  assign n4673 = ( n4474 & n4495 ) | ( n4474 & ~n4672 ) | ( n4495 & ~n4672 ) ;
  assign n4674 = ( n4474 & n4495 ) | ( n4474 & n4672 ) | ( n4495 & n4672 ) ;
  assign n4675 = ( n4672 & n4673 ) | ( n4672 & ~n4674 ) | ( n4673 & ~n4674 ) ;
  assign n4676 = ( n4453 & n4498 ) | ( n4453 & n4675 ) | ( n4498 & n4675 ) ;
  assign n4677 = ( n4453 & n4498 ) | ( n4453 & ~n4675 ) | ( n4498 & ~n4675 ) ;
  assign n4678 = ( n4675 & ~n4676 ) | ( n4675 & n4677 ) | ( ~n4676 & n4677 ) ;
  assign n4679 = ( n4521 & n4539 ) | ( n4521 & ~n4678 ) | ( n4539 & ~n4678 ) ;
  assign n4680 = ( n4521 & n4539 ) | ( n4521 & n4678 ) | ( n4539 & n4678 ) ;
  assign n4681 = ( n4678 & n4679 ) | ( n4678 & ~n4680 ) | ( n4679 & ~n4680 ) ;
  assign n4682 = ( n4550 & n4666 ) | ( n4550 & n4681 ) | ( n4666 & n4681 ) ;
  assign n4683 = ( n4550 & ~n4666 ) | ( n4550 & n4681 ) | ( ~n4666 & n4681 ) ;
  assign n4684 = ( n4666 & ~n4682 ) | ( n4666 & n4683 ) | ( ~n4682 & n4683 ) ;
  assign n4685 = ( n4527 & n4647 ) | ( n4527 & n4684 ) | ( n4647 & n4684 ) ;
  assign n4686 = ( n4527 & ~n4647 ) | ( n4527 & n4684 ) | ( ~n4647 & n4684 ) ;
  assign n4687 = ( n4647 & ~n4685 ) | ( n4647 & n4686 ) | ( ~n4685 & n4686 ) ;
  assign n4688 = ( n4565 & n4569 ) | ( n4565 & n4687 ) | ( n4569 & n4687 ) ;
  assign n4689 = ( n4565 & ~n4569 ) | ( n4565 & n4687 ) | ( ~n4569 & n4687 ) ;
  assign n4690 = ( n4569 & ~n4688 ) | ( n4569 & n4689 ) | ( ~n4688 & n4689 ) ;
  assign n4691 = ( n4659 & n4662 ) | ( n4659 & ~n4676 ) | ( n4662 & ~n4676 ) ;
  assign n4692 = ( n4659 & n4662 ) | ( n4659 & n4676 ) | ( n4662 & n4676 ) ;
  assign n4693 = ( n4676 & n4691 ) | ( n4676 & ~n4692 ) | ( n4691 & ~n4692 ) ;
  assign n4694 = x26 & x42 ;
  assign n4695 = x24 & x44 ;
  assign n4696 = x25 & x43 ;
  assign n4697 = ( ~n4694 & n4695 ) | ( ~n4694 & n4696 ) | ( n4695 & n4696 ) ;
  assign n4698 = ( n4694 & n4695 ) | ( n4694 & n4696 ) | ( n4695 & n4696 ) ;
  assign n4699 = ( n4694 & n4697 ) | ( n4694 & ~n4698 ) | ( n4697 & ~n4698 ) ;
  assign n4700 = x22 & x46 ;
  assign n4701 = x23 & x45 ;
  assign n4702 = x20 & x48 ;
  assign n4703 = ( ~n4700 & n4701 ) | ( ~n4700 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4704 = ( n4700 & n4701 ) | ( n4700 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4705 = ( n4700 & n4703 ) | ( n4700 & ~n4704 ) | ( n4703 & ~n4704 ) ;
  assign n4706 = x14 & x54 ;
  assign n4707 = x15 & x53 ;
  assign n4708 = x16 & x52 ;
  assign n4709 = ( ~n4706 & n4707 ) | ( ~n4706 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4710 = ( n4706 & n4707 ) | ( n4706 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4711 = ( n4706 & n4709 ) | ( n4706 & ~n4710 ) | ( n4709 & ~n4710 ) ;
  assign n4712 = ( ~n4699 & n4705 ) | ( ~n4699 & n4711 ) | ( n4705 & n4711 ) ;
  assign n4713 = ( n4699 & n4705 ) | ( n4699 & n4711 ) | ( n4705 & n4711 ) ;
  assign n4714 = ( n4699 & n4712 ) | ( n4699 & ~n4713 ) | ( n4712 & ~n4713 ) ;
  assign n4715 = x33 & x35 ;
  assign n4716 = x19 & x49 ;
  assign n4717 = x18 & x50 ;
  assign n4718 = ( ~n4715 & n4716 ) | ( ~n4715 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4719 = ( n4715 & n4716 ) | ( n4715 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4720 = ( n4715 & n4718 ) | ( n4715 & ~n4719 ) | ( n4718 & ~n4719 ) ;
  assign n4721 = x32 & x36 ;
  assign n4722 = x31 & x37 ;
  assign n4723 = x30 & x38 ;
  assign n4724 = ( ~n4721 & n4722 ) | ( ~n4721 & n4723 ) | ( n4722 & n4723 ) ;
  assign n4725 = ( n4721 & n4722 ) | ( n4721 & n4723 ) | ( n4722 & n4723 ) ;
  assign n4726 = ( n4721 & n4724 ) | ( n4721 & ~n4725 ) | ( n4724 & ~n4725 ) ;
  assign n4727 = x17 & x51 ;
  assign n4728 = x13 & x55 ;
  assign n4729 = x12 & x56 ;
  assign n4730 = ( ~n4727 & n4728 ) | ( ~n4727 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = ( n4727 & n4728 ) | ( n4727 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4732 = ( n4727 & n4730 ) | ( n4727 & ~n4731 ) | ( n4730 & ~n4731 ) ;
  assign n4733 = ( ~n4720 & n4726 ) | ( ~n4720 & n4732 ) | ( n4726 & n4732 ) ;
  assign n4734 = ( n4720 & n4726 ) | ( n4720 & n4732 ) | ( n4726 & n4732 ) ;
  assign n4735 = ( n4720 & n4733 ) | ( n4720 & ~n4734 ) | ( n4733 & ~n4734 ) ;
  assign n4736 = x21 & x47 ;
  assign n4737 = x5 & x63 ;
  assign n4738 = x6 & x62 ;
  assign n4739 = ( ~n4736 & n4737 ) | ( ~n4736 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4740 = ( n4736 & n4737 ) | ( n4736 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4741 = ( n4736 & n4739 ) | ( n4736 & ~n4740 ) | ( n4739 & ~n4740 ) ;
  assign n4742 = x11 & x57 ;
  assign n4743 = x9 & x59 ;
  assign n4744 = x10 & x58 ;
  assign n4745 = ( ~n4742 & n4743 ) | ( ~n4742 & n4744 ) | ( n4743 & n4744 ) ;
  assign n4746 = ( n4742 & n4743 ) | ( n4742 & n4744 ) | ( n4743 & n4744 ) ;
  assign n4747 = ( n4742 & n4745 ) | ( n4742 & ~n4746 ) | ( n4745 & ~n4746 ) ;
  assign n4748 = x29 & x39 ;
  assign n4749 = x27 & x41 ;
  assign n4750 = x28 & x40 ;
  assign n4751 = ( ~n4748 & n4749 ) | ( ~n4748 & n4750 ) | ( n4749 & n4750 ) ;
  assign n4752 = ( n4748 & n4749 ) | ( n4748 & n4750 ) | ( n4749 & n4750 ) ;
  assign n4753 = ( n4748 & n4751 ) | ( n4748 & ~n4752 ) | ( n4751 & ~n4752 ) ;
  assign n4754 = ( ~n4741 & n4747 ) | ( ~n4741 & n4753 ) | ( n4747 & n4753 ) ;
  assign n4755 = ( n4741 & n4747 ) | ( n4741 & n4753 ) | ( n4747 & n4753 ) ;
  assign n4756 = ( n4741 & n4754 ) | ( n4741 & ~n4755 ) | ( n4754 & ~n4755 ) ;
  assign n4757 = ( ~n4714 & n4735 ) | ( ~n4714 & n4756 ) | ( n4735 & n4756 ) ;
  assign n4758 = ( n4714 & n4735 ) | ( n4714 & n4756 ) | ( n4735 & n4756 ) ;
  assign n4759 = ( n4714 & n4757 ) | ( n4714 & ~n4758 ) | ( n4757 & ~n4758 ) ;
  assign n4760 = ( ~n4680 & n4693 ) | ( ~n4680 & n4759 ) | ( n4693 & n4759 ) ;
  assign n4761 = ( n4680 & n4693 ) | ( n4680 & n4759 ) | ( n4693 & n4759 ) ;
  assign n4762 = ( n4680 & n4760 ) | ( n4680 & ~n4761 ) | ( n4760 & ~n4761 ) ;
  assign n4763 = ( n4642 & n4682 ) | ( n4642 & n4762 ) | ( n4682 & n4762 ) ;
  assign n4764 = ( n4642 & n4682 ) | ( n4642 & ~n4762 ) | ( n4682 & ~n4762 ) ;
  assign n4765 = ( n4762 & ~n4763 ) | ( n4762 & n4764 ) | ( ~n4763 & n4764 ) ;
  assign n4766 = ( ~n4581 & n4608 ) | ( ~n4581 & n4628 ) | ( n4608 & n4628 ) ;
  assign n4767 = ( n4581 & n4608 ) | ( n4581 & n4628 ) | ( n4608 & n4628 ) ;
  assign n4768 = ( n4581 & n4766 ) | ( n4581 & ~n4767 ) | ( n4766 & ~n4767 ) ;
  assign n4769 = ( n4602 & ~n4614 ) | ( n4602 & n4671 ) | ( ~n4614 & n4671 ) ;
  assign n4770 = ( n4602 & n4614 ) | ( n4602 & n4671 ) | ( n4614 & n4671 ) ;
  assign n4771 = ( n4614 & n4769 ) | ( n4614 & ~n4770 ) | ( n4769 & ~n4770 ) ;
  assign n4772 = ( n4571 & n4768 ) | ( n4571 & n4771 ) | ( n4768 & n4771 ) ;
  assign n4773 = ( ~n4571 & n4768 ) | ( ~n4571 & n4771 ) | ( n4768 & n4771 ) ;
  assign n4774 = ( n4571 & ~n4772 ) | ( n4571 & n4773 ) | ( ~n4772 & n4773 ) ;
  assign n4775 = ( ~n4587 & n4593 ) | ( ~n4587 & n4634 ) | ( n4593 & n4634 ) ;
  assign n4776 = ( n4587 & n4593 ) | ( n4587 & n4634 ) | ( n4593 & n4634 ) ;
  assign n4777 = ( n4587 & n4775 ) | ( n4587 & ~n4776 ) | ( n4775 & ~n4776 ) ;
  assign n4778 = ( n4596 & n4637 ) | ( n4596 & n4777 ) | ( n4637 & n4777 ) ;
  assign n4779 = ( ~n4596 & n4637 ) | ( ~n4596 & n4777 ) | ( n4637 & n4777 ) ;
  assign n4780 = ( n4596 & ~n4778 ) | ( n4596 & n4779 ) | ( ~n4778 & n4779 ) ;
  assign n4781 = ( n4574 & n4774 ) | ( n4574 & n4780 ) | ( n4774 & n4780 ) ;
  assign n4782 = ( ~n4574 & n4774 ) | ( ~n4574 & n4780 ) | ( n4774 & n4780 ) ;
  assign n4783 = ( n4574 & ~n4781 ) | ( n4574 & n4782 ) | ( ~n4781 & n4782 ) ;
  assign n4784 = x7 & x61 ;
  assign n4785 = x8 & x60 ;
  assign n4786 = ( n4622 & n4784 ) | ( n4622 & n4785 ) | ( n4784 & n4785 ) ;
  assign n4787 = ( ~n4622 & n4784 ) | ( ~n4622 & n4785 ) | ( n4784 & n4785 ) ;
  assign n4788 = ( n4622 & ~n4786 ) | ( n4622 & n4787 ) | ( ~n4786 & n4787 ) ;
  assign n4789 = ( n4649 & n4655 ) | ( n4649 & n4788 ) | ( n4655 & n4788 ) ;
  assign n4790 = ( n4649 & n4655 ) | ( n4649 & ~n4788 ) | ( n4655 & ~n4788 ) ;
  assign n4791 = ( n4788 & ~n4789 ) | ( n4788 & n4790 ) | ( ~n4789 & n4790 ) ;
  assign n4792 = ( n4617 & n4652 ) | ( n4617 & n4674 ) | ( n4652 & n4674 ) ;
  assign n4793 = ( ~n4617 & n4652 ) | ( ~n4617 & n4674 ) | ( n4652 & n4674 ) ;
  assign n4794 = ( n4617 & ~n4792 ) | ( n4617 & n4793 ) | ( ~n4792 & n4793 ) ;
  assign n4795 = ( n4640 & n4791 ) | ( n4640 & n4794 ) | ( n4791 & n4794 ) ;
  assign n4796 = ( n4640 & ~n4791 ) | ( n4640 & n4794 ) | ( ~n4791 & n4794 ) ;
  assign n4797 = ( n4791 & ~n4795 ) | ( n4791 & n4796 ) | ( ~n4795 & n4796 ) ;
  assign n4798 = ( n4664 & n4783 ) | ( n4664 & n4797 ) | ( n4783 & n4797 ) ;
  assign n4799 = ( n4664 & ~n4783 ) | ( n4664 & n4797 ) | ( ~n4783 & n4797 ) ;
  assign n4800 = ( n4783 & ~n4798 ) | ( n4783 & n4799 ) | ( ~n4798 & n4799 ) ;
  assign n4801 = ( n4645 & ~n4765 ) | ( n4645 & n4800 ) | ( ~n4765 & n4800 ) ;
  assign n4802 = ( n4645 & n4765 ) | ( n4645 & n4800 ) | ( n4765 & n4800 ) ;
  assign n4803 = ( n4765 & n4801 ) | ( n4765 & ~n4802 ) | ( n4801 & ~n4802 ) ;
  assign n4804 = ( n4685 & n4688 ) | ( n4685 & n4803 ) | ( n4688 & n4803 ) ;
  assign n4805 = ( n4685 & ~n4688 ) | ( n4685 & n4803 ) | ( ~n4688 & n4803 ) ;
  assign n4806 = ( n4688 & ~n4804 ) | ( n4688 & n4805 ) | ( ~n4804 & n4805 ) ;
  assign n4807 = x21 & x48 ;
  assign n4808 = x22 & x47 ;
  assign n4809 = x14 & x55 ;
  assign n4810 = ( ~n4807 & n4808 ) | ( ~n4807 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4811 = ( n4807 & n4808 ) | ( n4807 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4812 = ( n4807 & n4810 ) | ( n4807 & ~n4811 ) | ( n4810 & ~n4811 ) ;
  assign n4813 = x13 & x56 ;
  assign n4814 = x11 & x58 ;
  assign n4815 = x12 & x57 ;
  assign n4816 = ( ~n4813 & n4814 ) | ( ~n4813 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4817 = ( n4813 & n4814 ) | ( n4813 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4818 = ( n4813 & n4816 ) | ( n4813 & ~n4817 ) | ( n4816 & ~n4817 ) ;
  assign n4819 = ( ~n4786 & n4812 ) | ( ~n4786 & n4818 ) | ( n4812 & n4818 ) ;
  assign n4820 = ( n4786 & n4812 ) | ( n4786 & n4818 ) | ( n4812 & n4818 ) ;
  assign n4821 = ( n4786 & n4819 ) | ( n4786 & ~n4820 ) | ( n4819 & ~n4820 ) ;
  assign n4822 = x27 & x42 ;
  assign n4823 = x26 & x43 ;
  assign n4824 = x6 & x63 ;
  assign n4825 = ( ~n4822 & n4823 ) | ( ~n4822 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4826 = ( n4822 & n4823 ) | ( n4822 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4827 = ( n4822 & n4825 ) | ( n4822 & ~n4826 ) | ( n4825 & ~n4826 ) ;
  assign n4828 = x10 & x59 ;
  assign n4829 = x9 & x60 ;
  assign n4830 = x8 & x61 ;
  assign n4831 = ( ~n4828 & n4829 ) | ( ~n4828 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4832 = ( n4828 & n4829 ) | ( n4828 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4833 = ( n4828 & n4831 ) | ( n4828 & ~n4832 ) | ( n4831 & ~n4832 ) ;
  assign n4834 = x24 & x45 ;
  assign n4835 = x25 & x44 ;
  assign n4836 = x23 & x46 ;
  assign n4837 = ( ~n4834 & n4835 ) | ( ~n4834 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4838 = ( n4834 & n4835 ) | ( n4834 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4839 = ( n4834 & n4837 ) | ( n4834 & ~n4838 ) | ( n4837 & ~n4838 ) ;
  assign n4840 = ( ~n4827 & n4833 ) | ( ~n4827 & n4839 ) | ( n4833 & n4839 ) ;
  assign n4841 = ( n4827 & n4833 ) | ( n4827 & n4839 ) | ( n4833 & n4839 ) ;
  assign n4842 = ( n4827 & n4840 ) | ( n4827 & ~n4841 ) | ( n4840 & ~n4841 ) ;
  assign n4843 = ( n4792 & n4821 ) | ( n4792 & n4842 ) | ( n4821 & n4842 ) ;
  assign n4844 = ( ~n4792 & n4821 ) | ( ~n4792 & n4842 ) | ( n4821 & n4842 ) ;
  assign n4845 = ( n4792 & ~n4843 ) | ( n4792 & n4844 ) | ( ~n4843 & n4844 ) ;
  assign n4846 = x19 & x50 ;
  assign n4847 = x17 & x52 ;
  assign n4848 = x18 & x51 ;
  assign n4849 = ( ~n4846 & n4847 ) | ( ~n4846 & n4848 ) | ( n4847 & n4848 ) ;
  assign n4850 = ( n4846 & n4847 ) | ( n4846 & n4848 ) | ( n4847 & n4848 ) ;
  assign n4851 = ( n4846 & n4849 ) | ( n4846 & ~n4850 ) | ( n4849 & ~n4850 ) ;
  assign n4852 = x28 & x41 ;
  assign n4853 = x30 & x39 ;
  assign n4854 = x29 & x40 ;
  assign n4855 = ( ~n4852 & n4853 ) | ( ~n4852 & n4854 ) | ( n4853 & n4854 ) ;
  assign n4856 = ( n4852 & n4853 ) | ( n4852 & n4854 ) | ( n4853 & n4854 ) ;
  assign n4857 = ( n4852 & n4855 ) | ( n4852 & ~n4856 ) | ( n4855 & ~n4856 ) ;
  assign n4858 = ( ~n4770 & n4851 ) | ( ~n4770 & n4857 ) | ( n4851 & n4857 ) ;
  assign n4859 = ( n4770 & n4851 ) | ( n4770 & n4857 ) | ( n4851 & n4857 ) ;
  assign n4860 = ( n4770 & n4858 ) | ( n4770 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  assign n4861 = x7 & x62 ;
  assign n4862 = x34 & x35 ;
  assign n4863 = ( x35 & n4861 ) | ( x35 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4864 = ( x35 & ~n4861 ) | ( x35 & n4862 ) | ( ~n4861 & n4862 ) ;
  assign n4865 = ( n4861 & ~n4863 ) | ( n4861 & n4864 ) | ( ~n4863 & n4864 ) ;
  assign n4866 = x16 & x53 ;
  assign n4867 = x15 & x54 ;
  assign n4868 = x20 & x49 ;
  assign n4869 = ( ~n4866 & n4867 ) | ( ~n4866 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4870 = ( n4866 & n4867 ) | ( n4866 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4871 = ( n4866 & n4869 ) | ( n4866 & ~n4870 ) | ( n4869 & ~n4870 ) ;
  assign n4872 = x33 & x36 ;
  assign n4873 = x31 & x38 ;
  assign n4874 = x32 & x37 ;
  assign n4875 = ( ~n4872 & n4873 ) | ( ~n4872 & n4874 ) | ( n4873 & n4874 ) ;
  assign n4876 = ( n4872 & n4873 ) | ( n4872 & n4874 ) | ( n4873 & n4874 ) ;
  assign n4877 = ( n4872 & n4875 ) | ( n4872 & ~n4876 ) | ( n4875 & ~n4876 ) ;
  assign n4878 = ( ~n4865 & n4871 ) | ( ~n4865 & n4877 ) | ( n4871 & n4877 ) ;
  assign n4879 = ( n4865 & n4871 ) | ( n4865 & n4877 ) | ( n4871 & n4877 ) ;
  assign n4880 = ( n4865 & n4878 ) | ( n4865 & ~n4879 ) | ( n4878 & ~n4879 ) ;
  assign n4881 = ( n4778 & n4860 ) | ( n4778 & n4880 ) | ( n4860 & n4880 ) ;
  assign n4882 = ( ~n4778 & n4860 ) | ( ~n4778 & n4880 ) | ( n4860 & n4880 ) ;
  assign n4883 = ( n4778 & ~n4881 ) | ( n4778 & n4882 ) | ( ~n4881 & n4882 ) ;
  assign n4884 = ( n4795 & n4845 ) | ( n4795 & n4883 ) | ( n4845 & n4883 ) ;
  assign n4885 = ( ~n4795 & n4845 ) | ( ~n4795 & n4883 ) | ( n4845 & n4883 ) ;
  assign n4886 = ( n4795 & ~n4884 ) | ( n4795 & n4885 ) | ( ~n4884 & n4885 ) ;
  assign n4887 = ( n4761 & n4798 ) | ( n4761 & ~n4886 ) | ( n4798 & ~n4886 ) ;
  assign n4888 = ( n4761 & n4798 ) | ( n4761 & n4886 ) | ( n4798 & n4886 ) ;
  assign n4889 = ( n4886 & n4887 ) | ( n4886 & ~n4888 ) | ( n4887 & ~n4888 ) ;
  assign n4890 = ( n4713 & n4734 ) | ( n4713 & ~n4789 ) | ( n4734 & ~n4789 ) ;
  assign n4891 = ( n4713 & n4734 ) | ( n4713 & n4789 ) | ( n4734 & n4789 ) ;
  assign n4892 = ( n4789 & n4890 ) | ( n4789 & ~n4891 ) | ( n4890 & ~n4891 ) ;
  assign n4893 = ( ~n4710 & n4719 ) | ( ~n4710 & n4725 ) | ( n4719 & n4725 ) ;
  assign n4894 = ( n4710 & n4719 ) | ( n4710 & n4725 ) | ( n4719 & n4725 ) ;
  assign n4895 = ( n4710 & n4893 ) | ( n4710 & ~n4894 ) | ( n4893 & ~n4894 ) ;
  assign n4896 = ( ~n4704 & n4740 ) | ( ~n4704 & n4746 ) | ( n4740 & n4746 ) ;
  assign n4897 = ( n4704 & n4740 ) | ( n4704 & n4746 ) | ( n4740 & n4746 ) ;
  assign n4898 = ( n4704 & n4896 ) | ( n4704 & ~n4897 ) | ( n4896 & ~n4897 ) ;
  assign n4899 = ( n4755 & n4895 ) | ( n4755 & n4898 ) | ( n4895 & n4898 ) ;
  assign n4900 = ( ~n4755 & n4895 ) | ( ~n4755 & n4898 ) | ( n4895 & n4898 ) ;
  assign n4901 = ( n4755 & ~n4899 ) | ( n4755 & n4900 ) | ( ~n4899 & n4900 ) ;
  assign n4902 = ( n4692 & n4892 ) | ( n4692 & n4901 ) | ( n4892 & n4901 ) ;
  assign n4903 = ( ~n4692 & n4892 ) | ( ~n4692 & n4901 ) | ( n4892 & n4901 ) ;
  assign n4904 = ( n4692 & ~n4902 ) | ( n4692 & n4903 ) | ( ~n4902 & n4903 ) ;
  assign n4905 = ( ~n4698 & n4731 ) | ( ~n4698 & n4752 ) | ( n4731 & n4752 ) ;
  assign n4906 = ( n4698 & n4731 ) | ( n4698 & n4752 ) | ( n4731 & n4752 ) ;
  assign n4907 = ( n4698 & n4905 ) | ( n4698 & ~n4906 ) | ( n4905 & ~n4906 ) ;
  assign n4908 = ( n4767 & n4776 ) | ( n4767 & n4907 ) | ( n4776 & n4907 ) ;
  assign n4909 = ( n4767 & n4776 ) | ( n4767 & ~n4907 ) | ( n4776 & ~n4907 ) ;
  assign n4910 = ( n4907 & ~n4908 ) | ( n4907 & n4909 ) | ( ~n4908 & n4909 ) ;
  assign n4911 = ( n4758 & ~n4772 ) | ( n4758 & n4910 ) | ( ~n4772 & n4910 ) ;
  assign n4912 = ( n4758 & n4772 ) | ( n4758 & n4910 ) | ( n4772 & n4910 ) ;
  assign n4913 = ( n4772 & n4911 ) | ( n4772 & ~n4912 ) | ( n4911 & ~n4912 ) ;
  assign n4914 = ( n4781 & n4904 ) | ( n4781 & n4913 ) | ( n4904 & n4913 ) ;
  assign n4915 = ( n4781 & ~n4904 ) | ( n4781 & n4913 ) | ( ~n4904 & n4913 ) ;
  assign n4916 = ( n4904 & ~n4914 ) | ( n4904 & n4915 ) | ( ~n4914 & n4915 ) ;
  assign n4917 = ( n4763 & n4889 ) | ( n4763 & n4916 ) | ( n4889 & n4916 ) ;
  assign n4918 = ( n4763 & ~n4889 ) | ( n4763 & n4916 ) | ( ~n4889 & n4916 ) ;
  assign n4919 = ( n4889 & ~n4917 ) | ( n4889 & n4918 ) | ( ~n4917 & n4918 ) ;
  assign n4920 = ( n4802 & ~n4804 ) | ( n4802 & n4919 ) | ( ~n4804 & n4919 ) ;
  assign n4921 = ( n4802 & n4804 ) | ( n4802 & n4919 ) | ( n4804 & n4919 ) ;
  assign n4922 = ( n4804 & n4920 ) | ( n4804 & ~n4921 ) | ( n4920 & ~n4921 ) ;
  assign n4923 = x34 & x36 ;
  assign n4924 = x32 & x38 ;
  assign n4925 = x33 & x37 ;
  assign n4926 = ( ~n4923 & n4924 ) | ( ~n4923 & n4925 ) | ( n4924 & n4925 ) ;
  assign n4927 = ( n4923 & n4924 ) | ( n4923 & n4925 ) | ( n4924 & n4925 ) ;
  assign n4928 = ( n4923 & n4926 ) | ( n4923 & ~n4927 ) | ( n4926 & ~n4927 ) ;
  assign n4929 = ( n4850 & n4870 ) | ( n4850 & ~n4928 ) | ( n4870 & ~n4928 ) ;
  assign n4930 = ( n4850 & n4870 ) | ( n4850 & n4928 ) | ( n4870 & n4928 ) ;
  assign n4931 = ( n4928 & n4929 ) | ( n4928 & ~n4930 ) | ( n4929 & ~n4930 ) ;
  assign n4932 = x18 & x52 ;
  assign n4933 = x16 & x54 ;
  assign n4934 = x17 & x53 ;
  assign n4935 = ( ~n4932 & n4933 ) | ( ~n4932 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4936 = ( n4932 & n4933 ) | ( n4932 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4937 = ( n4932 & n4935 ) | ( n4932 & ~n4936 ) | ( n4935 & ~n4936 ) ;
  assign n4938 = x11 & x59 ;
  assign n4939 = x9 & x61 ;
  assign n4940 = x10 & x60 ;
  assign n4941 = ( ~n4938 & n4939 ) | ( ~n4938 & n4940 ) | ( n4939 & n4940 ) ;
  assign n4942 = ( n4938 & n4939 ) | ( n4938 & n4940 ) | ( n4939 & n4940 ) ;
  assign n4943 = ( n4938 & n4941 ) | ( n4938 & ~n4942 ) | ( n4941 & ~n4942 ) ;
  assign n4944 = x12 & x58 ;
  assign n4945 = x13 & x57 ;
  assign n4946 = ( ~n2308 & n4944 ) | ( ~n2308 & n4945 ) | ( n4944 & n4945 ) ;
  assign n4947 = ( n2308 & n4944 ) | ( n2308 & n4945 ) | ( n4944 & n4945 ) ;
  assign n4948 = ( n2308 & n4946 ) | ( n2308 & ~n4947 ) | ( n4946 & ~n4947 ) ;
  assign n4949 = ( ~n4937 & n4943 ) | ( ~n4937 & n4948 ) | ( n4943 & n4948 ) ;
  assign n4950 = ( n4937 & n4943 ) | ( n4937 & n4948 ) | ( n4943 & n4948 ) ;
  assign n4951 = ( n4937 & n4949 ) | ( n4937 & ~n4950 ) | ( n4949 & ~n4950 ) ;
  assign n4952 = ( n4908 & n4931 ) | ( n4908 & n4951 ) | ( n4931 & n4951 ) ;
  assign n4953 = ( ~n4908 & n4931 ) | ( ~n4908 & n4951 ) | ( n4931 & n4951 ) ;
  assign n4954 = ( n4908 & ~n4952 ) | ( n4908 & n4953 ) | ( ~n4952 & n4953 ) ;
  assign n4955 = x30 & x40 ;
  assign n4956 = x31 & x39 ;
  assign n4957 = x29 & x41 ;
  assign n4958 = ( ~n4955 & n4956 ) | ( ~n4955 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4959 = ( n4955 & n4956 ) | ( n4955 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4960 = ( n4955 & n4958 ) | ( n4955 & ~n4959 ) | ( n4958 & ~n4959 ) ;
  assign n4961 = x23 & x47 ;
  assign n4962 = x7 & x63 ;
  assign n4963 = x28 & x42 ;
  assign n4964 = ( ~n4961 & n4962 ) | ( ~n4961 & n4963 ) | ( n4962 & n4963 ) ;
  assign n4965 = ( n4961 & n4962 ) | ( n4961 & n4963 ) | ( n4962 & n4963 ) ;
  assign n4966 = ( n4961 & n4964 ) | ( n4961 & ~n4965 ) | ( n4964 & ~n4965 ) ;
  assign n4967 = ( ~n4894 & n4960 ) | ( ~n4894 & n4966 ) | ( n4960 & n4966 ) ;
  assign n4968 = ( n4894 & n4960 ) | ( n4894 & n4966 ) | ( n4960 & n4966 ) ;
  assign n4969 = ( n4894 & n4967 ) | ( n4894 & ~n4968 ) | ( n4967 & ~n4968 ) ;
  assign n4970 = x15 & x55 ;
  assign n4971 = x14 & x56 ;
  assign n4972 = x22 & x48 ;
  assign n4973 = ( ~n4970 & n4971 ) | ( ~n4970 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = ( n4970 & n4971 ) | ( n4970 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4975 = ( n4970 & n4973 ) | ( n4970 & ~n4974 ) | ( n4973 & ~n4974 ) ;
  assign n4976 = x26 & x44 ;
  assign n4977 = x25 & x45 ;
  assign n4978 = x27 & x43 ;
  assign n4979 = ( ~n4976 & n4977 ) | ( ~n4976 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4980 = ( n4976 & n4977 ) | ( n4976 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4981 = ( n4976 & n4979 ) | ( n4976 & ~n4980 ) | ( n4979 & ~n4980 ) ;
  assign n4982 = x21 & x49 ;
  assign n4983 = x19 & x51 ;
  assign n4984 = x20 & x50 ;
  assign n4985 = ( ~n4982 & n4983 ) | ( ~n4982 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4986 = ( n4982 & n4983 ) | ( n4982 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4987 = ( n4982 & n4985 ) | ( n4982 & ~n4986 ) | ( n4985 & ~n4986 ) ;
  assign n4988 = ( ~n4975 & n4981 ) | ( ~n4975 & n4987 ) | ( n4981 & n4987 ) ;
  assign n4989 = ( n4975 & n4981 ) | ( n4975 & n4987 ) | ( n4981 & n4987 ) ;
  assign n4990 = ( n4975 & n4988 ) | ( n4975 & ~n4989 ) | ( n4988 & ~n4989 ) ;
  assign n4991 = ( n4899 & n4969 ) | ( n4899 & n4990 ) | ( n4969 & n4990 ) ;
  assign n4992 = ( ~n4899 & n4969 ) | ( ~n4899 & n4990 ) | ( n4969 & n4990 ) ;
  assign n4993 = ( n4899 & ~n4991 ) | ( n4899 & n4992 ) | ( ~n4991 & n4992 ) ;
  assign n4994 = ( n4912 & ~n4954 ) | ( n4912 & n4993 ) | ( ~n4954 & n4993 ) ;
  assign n4995 = ( n4912 & n4954 ) | ( n4912 & n4993 ) | ( n4954 & n4993 ) ;
  assign n4996 = ( n4954 & n4994 ) | ( n4954 & ~n4995 ) | ( n4994 & ~n4995 ) ;
  assign n4997 = ( n4826 & n4838 ) | ( n4826 & ~n4856 ) | ( n4838 & ~n4856 ) ;
  assign n4998 = ( n4826 & n4838 ) | ( n4826 & n4856 ) | ( n4838 & n4856 ) ;
  assign n4999 = ( n4856 & n4997 ) | ( n4856 & ~n4998 ) | ( n4997 & ~n4998 ) ;
  assign n5000 = x8 & x62 ;
  assign n5001 = ( n4863 & n4876 ) | ( n4863 & n5000 ) | ( n4876 & n5000 ) ;
  assign n5002 = ( n4863 & ~n4876 ) | ( n4863 & n5000 ) | ( ~n4876 & n5000 ) ;
  assign n5003 = ( n4876 & ~n5001 ) | ( n4876 & n5002 ) | ( ~n5001 & n5002 ) ;
  assign n5004 = ( n4859 & n4999 ) | ( n4859 & n5003 ) | ( n4999 & n5003 ) ;
  assign n5005 = ( ~n4859 & n4999 ) | ( ~n4859 & n5003 ) | ( n4999 & n5003 ) ;
  assign n5006 = ( n4859 & ~n5004 ) | ( n4859 & n5005 ) | ( ~n5004 & n5005 ) ;
  assign n5007 = ( ~n4820 & n4841 ) | ( ~n4820 & n4879 ) | ( n4841 & n4879 ) ;
  assign n5008 = ( n4820 & n4841 ) | ( n4820 & n4879 ) | ( n4841 & n4879 ) ;
  assign n5009 = ( n4820 & n5007 ) | ( n4820 & ~n5008 ) | ( n5007 & ~n5008 ) ;
  assign n5010 = ( n4881 & n5006 ) | ( n4881 & n5009 ) | ( n5006 & n5009 ) ;
  assign n5011 = ( n4881 & ~n5006 ) | ( n4881 & n5009 ) | ( ~n5006 & n5009 ) ;
  assign n5012 = ( n5006 & ~n5010 ) | ( n5006 & n5011 ) | ( ~n5010 & n5011 ) ;
  assign n5013 = ( ~n4914 & n4996 ) | ( ~n4914 & n5012 ) | ( n4996 & n5012 ) ;
  assign n5014 = ( n4914 & n4996 ) | ( n4914 & n5012 ) | ( n4996 & n5012 ) ;
  assign n5015 = ( n4914 & n5013 ) | ( n4914 & ~n5014 ) | ( n5013 & ~n5014 ) ;
  assign n5016 = ( n4811 & n4817 ) | ( n4811 & ~n4832 ) | ( n4817 & ~n4832 ) ;
  assign n5017 = ( n4811 & n4817 ) | ( n4811 & n4832 ) | ( n4817 & n4832 ) ;
  assign n5018 = ( n4832 & n5016 ) | ( n4832 & ~n5017 ) | ( n5016 & ~n5017 ) ;
  assign n5019 = ( n4897 & n4906 ) | ( n4897 & n5018 ) | ( n4906 & n5018 ) ;
  assign n5020 = ( n4897 & n4906 ) | ( n4897 & ~n5018 ) | ( n4906 & ~n5018 ) ;
  assign n5021 = ( n5018 & ~n5019 ) | ( n5018 & n5020 ) | ( ~n5019 & n5020 ) ;
  assign n5022 = ( ~n4843 & n4891 ) | ( ~n4843 & n5021 ) | ( n4891 & n5021 ) ;
  assign n5023 = ( n4843 & n4891 ) | ( n4843 & n5021 ) | ( n4891 & n5021 ) ;
  assign n5024 = ( n4843 & n5022 ) | ( n4843 & ~n5023 ) | ( n5022 & ~n5023 ) ;
  assign n5025 = ( n4884 & n4902 ) | ( n4884 & n5024 ) | ( n4902 & n5024 ) ;
  assign n5026 = ( n4884 & ~n4902 ) | ( n4884 & n5024 ) | ( ~n4902 & n5024 ) ;
  assign n5027 = ( n4902 & ~n5025 ) | ( n4902 & n5026 ) | ( ~n5025 & n5026 ) ;
  assign n5028 = ( n4888 & n5015 ) | ( n4888 & n5027 ) | ( n5015 & n5027 ) ;
  assign n5029 = ( n4888 & ~n5015 ) | ( n4888 & n5027 ) | ( ~n5015 & n5027 ) ;
  assign n5030 = ( n5015 & ~n5028 ) | ( n5015 & n5029 ) | ( ~n5028 & n5029 ) ;
  assign n5031 = ( n4917 & n4921 ) | ( n4917 & n5030 ) | ( n4921 & n5030 ) ;
  assign n5032 = ( n4917 & ~n4921 ) | ( n4917 & n5030 ) | ( ~n4921 & n5030 ) ;
  assign n5033 = ( n4921 & ~n5031 ) | ( n4921 & n5032 ) | ( ~n5031 & n5032 ) ;
  assign n5034 = x22 & x49 ;
  assign n5035 = x9 & x62 ;
  assign n5036 = ( ~x36 & n5034 ) | ( ~x36 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5037 = ( x36 & n5034 ) | ( x36 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5038 = ( x36 & n5036 ) | ( x36 & ~n5037 ) | ( n5036 & ~n5037 ) ;
  assign n5039 = x35 & x36 ;
  assign n5040 = x33 & x38 ;
  assign n5041 = x34 & x37 ;
  assign n5042 = ( ~n5039 & n5040 ) | ( ~n5039 & n5041 ) | ( n5040 & n5041 ) ;
  assign n5043 = ( n5039 & n5040 ) | ( n5039 & n5041 ) | ( n5040 & n5041 ) ;
  assign n5044 = ( n5039 & n5042 ) | ( n5039 & ~n5043 ) | ( n5042 & ~n5043 ) ;
  assign n5045 = x20 & x51 ;
  assign n5046 = x21 & x50 ;
  assign n5047 = x19 & x52 ;
  assign n5048 = ( ~n5045 & n5046 ) | ( ~n5045 & n5047 ) | ( n5046 & n5047 ) ;
  assign n5049 = ( n5045 & n5046 ) | ( n5045 & n5047 ) | ( n5046 & n5047 ) ;
  assign n5050 = ( n5045 & n5048 ) | ( n5045 & ~n5049 ) | ( n5048 & ~n5049 ) ;
  assign n5051 = ( ~n5038 & n5044 ) | ( ~n5038 & n5050 ) | ( n5044 & n5050 ) ;
  assign n5052 = ( n5038 & n5044 ) | ( n5038 & n5050 ) | ( n5044 & n5050 ) ;
  assign n5053 = ( n5038 & n5051 ) | ( n5038 & ~n5052 ) | ( n5051 & ~n5052 ) ;
  assign n5054 = x10 & x61 ;
  assign n5055 = x11 & x60 ;
  assign n5056 = x8 & x63 ;
  assign n5057 = ( ~n5054 & n5055 ) | ( ~n5054 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5058 = ( n5054 & n5055 ) | ( n5054 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5059 = ( n5054 & n5057 ) | ( n5054 & ~n5058 ) | ( n5057 & ~n5058 ) ;
  assign n5060 = ( n4927 & n4936 ) | ( n4927 & ~n5059 ) | ( n4936 & ~n5059 ) ;
  assign n5061 = ( n4927 & n4936 ) | ( n4927 & n5059 ) | ( n4936 & n5059 ) ;
  assign n5062 = ( n5059 & n5060 ) | ( n5059 & ~n5061 ) | ( n5060 & ~n5061 ) ;
  assign n5063 = ( n5019 & n5053 ) | ( n5019 & n5062 ) | ( n5053 & n5062 ) ;
  assign n5064 = ( ~n5019 & n5053 ) | ( ~n5019 & n5062 ) | ( n5053 & n5062 ) ;
  assign n5065 = ( n5019 & ~n5063 ) | ( n5019 & n5064 ) | ( ~n5063 & n5064 ) ;
  assign n5066 = x13 & x58 ;
  assign n5067 = x12 & x59 ;
  assign n5068 = ( n4986 & n5066 ) | ( n4986 & n5067 ) | ( n5066 & n5067 ) ;
  assign n5069 = ( ~n4986 & n5066 ) | ( ~n4986 & n5067 ) | ( n5066 & n5067 ) ;
  assign n5070 = ( n4986 & ~n5068 ) | ( n4986 & n5069 ) | ( ~n5068 & n5069 ) ;
  assign n5071 = x16 & x55 ;
  assign n5072 = x14 & x57 ;
  assign n5073 = x15 & x56 ;
  assign n5074 = ( ~n5071 & n5072 ) | ( ~n5071 & n5073 ) | ( n5072 & n5073 ) ;
  assign n5075 = ( n5071 & n5072 ) | ( n5071 & n5073 ) | ( n5072 & n5073 ) ;
  assign n5076 = ( n5071 & n5074 ) | ( n5071 & ~n5075 ) | ( n5074 & ~n5075 ) ;
  assign n5077 = x26 & x45 ;
  assign n5078 = x24 & x47 ;
  assign n5079 = x25 & x46 ;
  assign n5080 = ( ~n5077 & n5078 ) | ( ~n5077 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5081 = ( n5077 & n5078 ) | ( n5077 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5082 = ( n5077 & n5080 ) | ( n5077 & ~n5081 ) | ( n5080 & ~n5081 ) ;
  assign n5083 = ( n5070 & n5076 ) | ( n5070 & n5082 ) | ( n5076 & n5082 ) ;
  assign n5084 = ( ~n5070 & n5076 ) | ( ~n5070 & n5082 ) | ( n5076 & n5082 ) ;
  assign n5085 = ( n5070 & ~n5083 ) | ( n5070 & n5084 ) | ( ~n5083 & n5084 ) ;
  assign n5086 = x31 & x40 ;
  assign n5087 = x30 & x41 ;
  assign n5088 = x32 & x39 ;
  assign n5089 = ( ~n5086 & n5087 ) | ( ~n5086 & n5088 ) | ( n5087 & n5088 ) ;
  assign n5090 = ( n5086 & n5087 ) | ( n5086 & n5088 ) | ( n5087 & n5088 ) ;
  assign n5091 = ( n5086 & n5089 ) | ( n5086 & ~n5090 ) | ( n5089 & ~n5090 ) ;
  assign n5092 = x28 & x43 ;
  assign n5093 = x29 & x42 ;
  assign n5094 = x27 & x44 ;
  assign n5095 = ( ~n5092 & n5093 ) | ( ~n5092 & n5094 ) | ( n5093 & n5094 ) ;
  assign n5096 = ( n5092 & n5093 ) | ( n5092 & n5094 ) | ( n5093 & n5094 ) ;
  assign n5097 = ( n5092 & n5095 ) | ( n5092 & ~n5096 ) | ( n5095 & ~n5096 ) ;
  assign n5098 = x17 & x54 ;
  assign n5099 = x18 & x53 ;
  assign n5100 = x23 & x48 ;
  assign n5101 = ( ~n5098 & n5099 ) | ( ~n5098 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ( n5098 & n5099 ) | ( n5098 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5103 = ( n5098 & n5101 ) | ( n5098 & ~n5102 ) | ( n5101 & ~n5102 ) ;
  assign n5104 = ( ~n5091 & n5097 ) | ( ~n5091 & n5103 ) | ( n5097 & n5103 ) ;
  assign n5105 = ( n5091 & n5097 ) | ( n5091 & n5103 ) | ( n5097 & n5103 ) ;
  assign n5106 = ( n5091 & n5104 ) | ( n5091 & ~n5105 ) | ( n5104 & ~n5105 ) ;
  assign n5107 = ( n5008 & n5085 ) | ( n5008 & n5106 ) | ( n5085 & n5106 ) ;
  assign n5108 = ( ~n5008 & n5085 ) | ( ~n5008 & n5106 ) | ( n5085 & n5106 ) ;
  assign n5109 = ( n5008 & ~n5107 ) | ( n5008 & n5108 ) | ( ~n5107 & n5108 ) ;
  assign n5110 = ( n5023 & n5065 ) | ( n5023 & n5109 ) | ( n5065 & n5109 ) ;
  assign n5111 = ( ~n5023 & n5065 ) | ( ~n5023 & n5109 ) | ( n5065 & n5109 ) ;
  assign n5112 = ( n5023 & ~n5110 ) | ( n5023 & n5111 ) | ( ~n5110 & n5111 ) ;
  assign n5113 = ( n4959 & n4965 ) | ( n4959 & ~n4974 ) | ( n4965 & ~n4974 ) ;
  assign n5114 = ( n4959 & n4965 ) | ( n4959 & n4974 ) | ( n4965 & n4974 ) ;
  assign n5115 = ( n4974 & n5113 ) | ( n4974 & ~n5114 ) | ( n5113 & ~n5114 ) ;
  assign n5116 = ( ~n4942 & n4947 ) | ( ~n4942 & n4980 ) | ( n4947 & n4980 ) ;
  assign n5117 = ( n4942 & n4947 ) | ( n4942 & n4980 ) | ( n4947 & n4980 ) ;
  assign n5118 = ( n4942 & n5116 ) | ( n4942 & ~n5117 ) | ( n5116 & ~n5117 ) ;
  assign n5119 = ( n4968 & n5115 ) | ( n4968 & n5118 ) | ( n5115 & n5118 ) ;
  assign n5120 = ( ~n4968 & n5115 ) | ( ~n4968 & n5118 ) | ( n5115 & n5118 ) ;
  assign n5121 = ( n4968 & ~n5119 ) | ( n4968 & n5120 ) | ( ~n5119 & n5120 ) ;
  assign n5122 = ( n4950 & n4989 ) | ( n4950 & ~n5017 ) | ( n4989 & ~n5017 ) ;
  assign n5123 = ( n4950 & n4989 ) | ( n4950 & n5017 ) | ( n4989 & n5017 ) ;
  assign n5124 = ( n5017 & n5122 ) | ( n5017 & ~n5123 ) | ( n5122 & ~n5123 ) ;
  assign n5125 = ( n4991 & n5121 ) | ( n4991 & n5124 ) | ( n5121 & n5124 ) ;
  assign n5126 = ( n4991 & ~n5121 ) | ( n4991 & n5124 ) | ( ~n5121 & n5124 ) ;
  assign n5127 = ( n5121 & ~n5125 ) | ( n5121 & n5126 ) | ( ~n5125 & n5126 ) ;
  assign n5128 = ( n5025 & n5112 ) | ( n5025 & n5127 ) | ( n5112 & n5127 ) ;
  assign n5129 = ( ~n5025 & n5112 ) | ( ~n5025 & n5127 ) | ( n5112 & n5127 ) ;
  assign n5130 = ( n5025 & ~n5128 ) | ( n5025 & n5129 ) | ( ~n5128 & n5129 ) ;
  assign n5131 = ( n4930 & n4998 ) | ( n4930 & n5001 ) | ( n4998 & n5001 ) ;
  assign n5132 = ( ~n4930 & n4998 ) | ( ~n4930 & n5001 ) | ( n4998 & n5001 ) ;
  assign n5133 = ( n4930 & ~n5131 ) | ( n4930 & n5132 ) | ( ~n5131 & n5132 ) ;
  assign n5134 = ( n4952 & n5004 ) | ( n4952 & n5133 ) | ( n5004 & n5133 ) ;
  assign n5135 = ( n4952 & n5004 ) | ( n4952 & ~n5133 ) | ( n5004 & ~n5133 ) ;
  assign n5136 = ( n5133 & ~n5134 ) | ( n5133 & n5135 ) | ( ~n5134 & n5135 ) ;
  assign n5137 = ( ~n4995 & n5010 ) | ( ~n4995 & n5136 ) | ( n5010 & n5136 ) ;
  assign n5138 = ( n4995 & n5010 ) | ( n4995 & n5136 ) | ( n5010 & n5136 ) ;
  assign n5139 = ( n4995 & n5137 ) | ( n4995 & ~n5138 ) | ( n5137 & ~n5138 ) ;
  assign n5140 = ( ~n5014 & n5130 ) | ( ~n5014 & n5139 ) | ( n5130 & n5139 ) ;
  assign n5141 = ( n5014 & n5130 ) | ( n5014 & n5139 ) | ( n5130 & n5139 ) ;
  assign n5142 = ( n5014 & n5140 ) | ( n5014 & ~n5141 ) | ( n5140 & ~n5141 ) ;
  assign n5143 = ( n5028 & ~n5031 ) | ( n5028 & n5142 ) | ( ~n5031 & n5142 ) ;
  assign n5144 = ( n5028 & n5031 ) | ( n5028 & n5142 ) | ( n5031 & n5142 ) ;
  assign n5145 = ( n5031 & n5143 ) | ( n5031 & ~n5144 ) | ( n5143 & ~n5144 ) ;
  assign n5146 = ( n5058 & ~n5075 ) | ( n5058 & n5081 ) | ( ~n5075 & n5081 ) ;
  assign n5147 = ( n5058 & n5075 ) | ( n5058 & n5081 ) | ( n5075 & n5081 ) ;
  assign n5148 = ( n5075 & n5146 ) | ( n5075 & ~n5147 ) | ( n5146 & ~n5147 ) ;
  assign n5149 = x19 & x53 ;
  assign n5150 = x33 & x39 ;
  assign n5151 = x34 & x38 ;
  assign n5152 = ( ~n5149 & n5150 ) | ( ~n5149 & n5151 ) | ( n5150 & n5151 ) ;
  assign n5153 = ( n5149 & n5150 ) | ( n5149 & n5151 ) | ( n5150 & n5151 ) ;
  assign n5154 = ( n5149 & n5152 ) | ( n5149 & ~n5153 ) | ( n5152 & ~n5153 ) ;
  assign n5155 = x15 & x57 ;
  assign n5156 = x13 & x59 ;
  assign n5157 = x14 & x58 ;
  assign n5158 = ( ~n5155 & n5156 ) | ( ~n5155 & n5157 ) | ( n5156 & n5157 ) ;
  assign n5159 = ( n5155 & n5156 ) | ( n5155 & n5157 ) | ( n5156 & n5157 ) ;
  assign n5160 = ( n5155 & n5158 ) | ( n5155 & ~n5159 ) | ( n5158 & ~n5159 ) ;
  assign n5161 = x28 & x44 ;
  assign n5162 = x27 & x45 ;
  assign n5163 = x26 & x46 ;
  assign n5164 = ( ~n5161 & n5162 ) | ( ~n5161 & n5163 ) | ( n5162 & n5163 ) ;
  assign n5165 = ( n5161 & n5162 ) | ( n5161 & n5163 ) | ( n5162 & n5163 ) ;
  assign n5166 = ( n5161 & n5164 ) | ( n5161 & ~n5165 ) | ( n5164 & ~n5165 ) ;
  assign n5167 = ( ~n5154 & n5160 ) | ( ~n5154 & n5166 ) | ( n5160 & n5166 ) ;
  assign n5168 = ( n5154 & n5160 ) | ( n5154 & n5166 ) | ( n5160 & n5166 ) ;
  assign n5169 = ( n5154 & n5167 ) | ( n5154 & ~n5168 ) | ( n5167 & ~n5168 ) ;
  assign n5170 = ( n5131 & n5148 ) | ( n5131 & n5169 ) | ( n5148 & n5169 ) ;
  assign n5171 = ( ~n5131 & n5148 ) | ( ~n5131 & n5169 ) | ( n5148 & n5169 ) ;
  assign n5172 = ( n5131 & ~n5170 ) | ( n5131 & n5171 ) | ( ~n5170 & n5171 ) ;
  assign n5173 = x24 & x48 ;
  assign n5174 = x12 & x60 ;
  assign n5175 = ( ~n2393 & n5173 ) | ( ~n2393 & n5174 ) | ( n5173 & n5174 ) ;
  assign n5176 = ( n2393 & n5173 ) | ( n2393 & n5174 ) | ( n5173 & n5174 ) ;
  assign n5177 = ( n2393 & n5175 ) | ( n2393 & ~n5176 ) | ( n5175 & ~n5176 ) ;
  assign n5178 = x10 & x62 ;
  assign n5179 = x11 & x61 ;
  assign n5180 = x9 & x63 ;
  assign n5181 = ( ~n5178 & n5179 ) | ( ~n5178 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5182 = ( n5178 & n5179 ) | ( n5178 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5183 = ( n5178 & n5181 ) | ( n5178 & ~n5182 ) | ( n5181 & ~n5182 ) ;
  assign n5184 = ( ~n5068 & n5177 ) | ( ~n5068 & n5183 ) | ( n5177 & n5183 ) ;
  assign n5185 = ( n5068 & n5177 ) | ( n5068 & n5183 ) | ( n5177 & n5183 ) ;
  assign n5186 = ( n5068 & n5184 ) | ( n5068 & ~n5185 ) | ( n5184 & ~n5185 ) ;
  assign n5187 = x32 & x40 ;
  assign n5188 = x23 & x49 ;
  assign n5189 = x16 & x56 ;
  assign n5190 = ( ~n5187 & n5188 ) | ( ~n5187 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = ( n5187 & n5188 ) | ( n5187 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5192 = ( n5187 & n5190 ) | ( n5187 & ~n5191 ) | ( n5190 & ~n5191 ) ;
  assign n5193 = x17 & x55 ;
  assign n5194 = x18 & x54 ;
  assign n5195 = x20 & x52 ;
  assign n5196 = ( ~n5193 & n5194 ) | ( ~n5193 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5197 = ( n5193 & n5194 ) | ( n5193 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5198 = ( n5193 & n5196 ) | ( n5193 & ~n5197 ) | ( n5196 & ~n5197 ) ;
  assign n5199 = x35 & x37 ;
  assign n5200 = x21 & x51 ;
  assign n5201 = x22 & x50 ;
  assign n5202 = ( ~n5199 & n5200 ) | ( ~n5199 & n5201 ) | ( n5200 & n5201 ) ;
  assign n5203 = ( n5199 & n5200 ) | ( n5199 & n5201 ) | ( n5200 & n5201 ) ;
  assign n5204 = ( n5199 & n5202 ) | ( n5199 & ~n5203 ) | ( n5202 & ~n5203 ) ;
  assign n5205 = ( ~n5192 & n5198 ) | ( ~n5192 & n5204 ) | ( n5198 & n5204 ) ;
  assign n5206 = ( n5192 & n5198 ) | ( n5192 & n5204 ) | ( n5198 & n5204 ) ;
  assign n5207 = ( n5192 & n5205 ) | ( n5192 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = ( n5123 & n5186 ) | ( n5123 & n5207 ) | ( n5186 & n5207 ) ;
  assign n5209 = ( ~n5123 & n5186 ) | ( ~n5123 & n5207 ) | ( n5186 & n5207 ) ;
  assign n5210 = ( n5123 & ~n5208 ) | ( n5123 & n5209 ) | ( ~n5208 & n5209 ) ;
  assign n5211 = ( n5134 & ~n5172 ) | ( n5134 & n5210 ) | ( ~n5172 & n5210 ) ;
  assign n5212 = ( n5134 & n5172 ) | ( n5134 & n5210 ) | ( n5172 & n5210 ) ;
  assign n5213 = ( n5172 & n5211 ) | ( n5172 & ~n5212 ) | ( n5211 & ~n5212 ) ;
  assign n5214 = ( n5037 & n5043 ) | ( n5037 & ~n5049 ) | ( n5043 & ~n5049 ) ;
  assign n5215 = ( n5037 & n5043 ) | ( n5037 & n5049 ) | ( n5043 & n5049 ) ;
  assign n5216 = ( n5049 & n5214 ) | ( n5049 & ~n5215 ) | ( n5214 & ~n5215 ) ;
  assign n5217 = ( ~n5090 & n5096 ) | ( ~n5090 & n5102 ) | ( n5096 & n5102 ) ;
  assign n5218 = ( n5090 & n5096 ) | ( n5090 & n5102 ) | ( n5096 & n5102 ) ;
  assign n5219 = ( n5090 & n5217 ) | ( n5090 & ~n5218 ) | ( n5217 & ~n5218 ) ;
  assign n5220 = ( n5083 & n5216 ) | ( n5083 & n5219 ) | ( n5216 & n5219 ) ;
  assign n5221 = ( ~n5083 & n5216 ) | ( ~n5083 & n5219 ) | ( n5216 & n5219 ) ;
  assign n5222 = ( n5083 & ~n5220 ) | ( n5083 & n5221 ) | ( ~n5220 & n5221 ) ;
  assign n5223 = ( n5052 & n5105 ) | ( n5052 & ~n5117 ) | ( n5105 & ~n5117 ) ;
  assign n5224 = ( n5052 & n5105 ) | ( n5052 & n5117 ) | ( n5105 & n5117 ) ;
  assign n5225 = ( n5117 & n5223 ) | ( n5117 & ~n5224 ) | ( n5223 & ~n5224 ) ;
  assign n5226 = ( n5107 & ~n5222 ) | ( n5107 & n5225 ) | ( ~n5222 & n5225 ) ;
  assign n5227 = ( n5107 & n5222 ) | ( n5107 & n5225 ) | ( n5222 & n5225 ) ;
  assign n5228 = ( n5222 & n5226 ) | ( n5222 & ~n5227 ) | ( n5226 & ~n5227 ) ;
  assign n5229 = ( n5138 & n5213 ) | ( n5138 & n5228 ) | ( n5213 & n5228 ) ;
  assign n5230 = ( ~n5138 & n5213 ) | ( ~n5138 & n5228 ) | ( n5213 & n5228 ) ;
  assign n5231 = ( n5138 & ~n5229 ) | ( n5138 & n5230 ) | ( ~n5229 & n5230 ) ;
  assign n5232 = x30 & x42 ;
  assign n5233 = x31 & x41 ;
  assign n5234 = x29 & x43 ;
  assign n5235 = ( ~n5232 & n5233 ) | ( ~n5232 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5236 = ( n5232 & n5233 ) | ( n5232 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5237 = ( n5232 & n5235 ) | ( n5232 & ~n5236 ) | ( n5235 & ~n5236 ) ;
  assign n5238 = ( n5061 & n5114 ) | ( n5061 & n5237 ) | ( n5114 & n5237 ) ;
  assign n5239 = ( ~n5061 & n5114 ) | ( ~n5061 & n5237 ) | ( n5114 & n5237 ) ;
  assign n5240 = ( n5061 & ~n5238 ) | ( n5061 & n5239 ) | ( ~n5238 & n5239 ) ;
  assign n5241 = ( n5063 & n5119 ) | ( n5063 & n5240 ) | ( n5119 & n5240 ) ;
  assign n5242 = ( n5063 & n5119 ) | ( n5063 & ~n5240 ) | ( n5119 & ~n5240 ) ;
  assign n5243 = ( n5240 & ~n5241 ) | ( n5240 & n5242 ) | ( ~n5241 & n5242 ) ;
  assign n5244 = ( n5110 & n5125 ) | ( n5110 & n5243 ) | ( n5125 & n5243 ) ;
  assign n5245 = ( ~n5110 & n5125 ) | ( ~n5110 & n5243 ) | ( n5125 & n5243 ) ;
  assign n5246 = ( n5110 & ~n5244 ) | ( n5110 & n5245 ) | ( ~n5244 & n5245 ) ;
  assign n5247 = ( n5128 & n5231 ) | ( n5128 & n5246 ) | ( n5231 & n5246 ) ;
  assign n5248 = ( n5128 & ~n5231 ) | ( n5128 & n5246 ) | ( ~n5231 & n5246 ) ;
  assign n5249 = ( n5231 & ~n5247 ) | ( n5231 & n5248 ) | ( ~n5247 & n5248 ) ;
  assign n5250 = ( n5141 & n5144 ) | ( n5141 & n5249 ) | ( n5144 & n5249 ) ;
  assign n5251 = ( n5141 & ~n5144 ) | ( n5141 & n5249 ) | ( ~n5144 & n5249 ) ;
  assign n5252 = ( n5144 & ~n5250 ) | ( n5144 & n5251 ) | ( ~n5250 & n5251 ) ;
  assign n5253 = x10 & x63 ;
  assign n5254 = x25 & x48 ;
  assign n5255 = x12 & x61 ;
  assign n5256 = ( ~n5253 & n5254 ) | ( ~n5253 & n5255 ) | ( n5254 & n5255 ) ;
  assign n5257 = ( n5253 & n5254 ) | ( n5253 & n5255 ) | ( n5254 & n5255 ) ;
  assign n5258 = ( n5253 & n5256 ) | ( n5253 & ~n5257 ) | ( n5256 & ~n5257 ) ;
  assign n5259 = x36 & x37 ;
  assign n5260 = x34 & x39 ;
  assign n5261 = x35 & x38 ;
  assign n5262 = ( ~n5259 & n5260 ) | ( ~n5259 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = ( n5259 & n5260 ) | ( n5259 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5264 = ( n5259 & n5262 ) | ( n5259 & ~n5263 ) | ( n5262 & ~n5263 ) ;
  assign n5265 = x29 & x44 ;
  assign n5266 = x30 & x43 ;
  assign n5267 = x28 & x45 ;
  assign n5268 = ( ~n5265 & n5266 ) | ( ~n5265 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = ( n5265 & n5266 ) | ( n5265 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5270 = ( n5265 & n5268 ) | ( n5265 & ~n5269 ) | ( n5268 & ~n5269 ) ;
  assign n5271 = ( ~n5258 & n5264 ) | ( ~n5258 & n5270 ) | ( n5264 & n5270 ) ;
  assign n5272 = ( n5258 & n5264 ) | ( n5258 & n5270 ) | ( n5264 & n5270 ) ;
  assign n5273 = ( n5258 & n5271 ) | ( n5258 & ~n5272 ) | ( n5271 & ~n5272 ) ;
  assign n5274 = ( ~n5159 & n5165 ) | ( ~n5159 & n5236 ) | ( n5165 & n5236 ) ;
  assign n5275 = ( n5159 & n5165 ) | ( n5159 & n5236 ) | ( n5165 & n5236 ) ;
  assign n5276 = ( n5159 & n5274 ) | ( n5159 & ~n5275 ) | ( n5274 & ~n5275 ) ;
  assign n5277 = ( n5238 & n5273 ) | ( n5238 & n5276 ) | ( n5273 & n5276 ) ;
  assign n5278 = ( ~n5238 & n5273 ) | ( ~n5238 & n5276 ) | ( n5273 & n5276 ) ;
  assign n5279 = ( n5238 & ~n5277 ) | ( n5238 & n5278 ) | ( ~n5277 & n5278 ) ;
  assign n5280 = x24 & x49 ;
  assign n5281 = x18 & x55 ;
  assign n5282 = x19 & x54 ;
  assign n5283 = ( ~n5280 & n5281 ) | ( ~n5280 & n5282 ) | ( n5281 & n5282 ) ;
  assign n5284 = ( n5280 & n5281 ) | ( n5280 & n5282 ) | ( n5281 & n5282 ) ;
  assign n5285 = ( n5280 & n5283 ) | ( n5280 & ~n5284 ) | ( n5283 & ~n5284 ) ;
  assign n5286 = x20 & x53 ;
  assign n5287 = x22 & x51 ;
  assign n5288 = x21 & x52 ;
  assign n5289 = ( ~n5286 & n5287 ) | ( ~n5286 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5290 = ( n5286 & n5287 ) | ( n5286 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5291 = ( n5286 & n5289 ) | ( n5286 & ~n5290 ) | ( n5289 & ~n5290 ) ;
  assign n5292 = x23 & x50 ;
  assign n5293 = x11 & x62 ;
  assign n5294 = ( ~x37 & n5292 ) | ( ~x37 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5295 = ( x37 & n5292 ) | ( x37 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5296 = ( x37 & n5294 ) | ( x37 & ~n5295 ) | ( n5294 & ~n5295 ) ;
  assign n5297 = ( ~n5285 & n5291 ) | ( ~n5285 & n5296 ) | ( n5291 & n5296 ) ;
  assign n5298 = ( n5285 & n5291 ) | ( n5285 & n5296 ) | ( n5291 & n5296 ) ;
  assign n5299 = ( n5285 & n5297 ) | ( n5285 & ~n5298 ) | ( n5297 & ~n5298 ) ;
  assign n5300 = x14 & x59 ;
  assign n5301 = x15 & x58 ;
  assign n5302 = x16 & x57 ;
  assign n5303 = ( ~n5300 & n5301 ) | ( ~n5300 & n5302 ) | ( n5301 & n5302 ) ;
  assign n5304 = ( n5300 & n5301 ) | ( n5300 & n5302 ) | ( n5301 & n5302 ) ;
  assign n5305 = ( n5300 & n5303 ) | ( n5300 & ~n5304 ) | ( n5303 & ~n5304 ) ;
  assign n5306 = x27 & x46 ;
  assign n5307 = x17 & x56 ;
  assign n5308 = x26 & x47 ;
  assign n5309 = ( ~n5306 & n5307 ) | ( ~n5306 & n5308 ) | ( n5307 & n5308 ) ;
  assign n5310 = ( n5306 & n5307 ) | ( n5306 & n5308 ) | ( n5307 & n5308 ) ;
  assign n5311 = ( n5306 & n5309 ) | ( n5306 & ~n5310 ) | ( n5309 & ~n5310 ) ;
  assign n5312 = ( ~n5191 & n5305 ) | ( ~n5191 & n5311 ) | ( n5305 & n5311 ) ;
  assign n5313 = ( n5191 & n5305 ) | ( n5191 & n5311 ) | ( n5305 & n5311 ) ;
  assign n5314 = ( n5191 & n5312 ) | ( n5191 & ~n5313 ) | ( n5312 & ~n5313 ) ;
  assign n5315 = ( n5224 & n5299 ) | ( n5224 & n5314 ) | ( n5299 & n5314 ) ;
  assign n5316 = ( ~n5224 & n5299 ) | ( ~n5224 & n5314 ) | ( n5299 & n5314 ) ;
  assign n5317 = ( n5224 & ~n5315 ) | ( n5224 & n5316 ) | ( ~n5315 & n5316 ) ;
  assign n5318 = ( n5241 & ~n5279 ) | ( n5241 & n5317 ) | ( ~n5279 & n5317 ) ;
  assign n5319 = ( n5241 & n5279 ) | ( n5241 & n5317 ) | ( n5279 & n5317 ) ;
  assign n5320 = ( n5279 & n5318 ) | ( n5279 & ~n5319 ) | ( n5318 & ~n5319 ) ;
  assign n5321 = ( n5168 & ~n5185 ) | ( n5168 & n5215 ) | ( ~n5185 & n5215 ) ;
  assign n5322 = ( n5168 & n5185 ) | ( n5168 & n5215 ) | ( n5185 & n5215 ) ;
  assign n5323 = ( n5185 & n5321 ) | ( n5185 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5324 = ( n5176 & n5182 ) | ( n5176 & ~n5197 ) | ( n5182 & ~n5197 ) ;
  assign n5325 = ( n5176 & n5182 ) | ( n5176 & n5197 ) | ( n5182 & n5197 ) ;
  assign n5326 = ( n5197 & n5324 ) | ( n5197 & ~n5325 ) | ( n5324 & ~n5325 ) ;
  assign n5327 = x13 & x60 ;
  assign n5328 = ( n5153 & n5203 ) | ( n5153 & n5327 ) | ( n5203 & n5327 ) ;
  assign n5329 = ( ~n5153 & n5203 ) | ( ~n5153 & n5327 ) | ( n5203 & n5327 ) ;
  assign n5330 = ( n5153 & ~n5328 ) | ( n5153 & n5329 ) | ( ~n5328 & n5329 ) ;
  assign n5331 = ( n5206 & n5326 ) | ( n5206 & n5330 ) | ( n5326 & n5330 ) ;
  assign n5332 = ( n5206 & ~n5326 ) | ( n5206 & n5330 ) | ( ~n5326 & n5330 ) ;
  assign n5333 = ( n5326 & ~n5331 ) | ( n5326 & n5332 ) | ( ~n5331 & n5332 ) ;
  assign n5334 = ( n5208 & ~n5323 ) | ( n5208 & n5333 ) | ( ~n5323 & n5333 ) ;
  assign n5335 = ( n5208 & n5323 ) | ( n5208 & n5333 ) | ( n5323 & n5333 ) ;
  assign n5336 = ( n5323 & n5334 ) | ( n5323 & ~n5335 ) | ( n5334 & ~n5335 ) ;
  assign n5337 = ( n5244 & n5320 ) | ( n5244 & n5336 ) | ( n5320 & n5336 ) ;
  assign n5338 = ( ~n5244 & n5320 ) | ( ~n5244 & n5336 ) | ( n5320 & n5336 ) ;
  assign n5339 = ( n5244 & ~n5337 ) | ( n5244 & n5338 ) | ( ~n5337 & n5338 ) ;
  assign n5340 = x31 & x42 ;
  assign n5341 = x33 & x40 ;
  assign n5342 = x32 & x41 ;
  assign n5343 = ( ~n5340 & n5341 ) | ( ~n5340 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = ( n5340 & n5341 ) | ( n5340 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5345 = ( n5340 & n5343 ) | ( n5340 & ~n5344 ) | ( n5343 & ~n5344 ) ;
  assign n5346 = ( ~n5147 & n5218 ) | ( ~n5147 & n5345 ) | ( n5218 & n5345 ) ;
  assign n5347 = ( n5147 & n5218 ) | ( n5147 & n5345 ) | ( n5218 & n5345 ) ;
  assign n5348 = ( n5147 & n5346 ) | ( n5147 & ~n5347 ) | ( n5346 & ~n5347 ) ;
  assign n5349 = ( n5170 & ~n5220 ) | ( n5170 & n5348 ) | ( ~n5220 & n5348 ) ;
  assign n5350 = ( n5170 & n5220 ) | ( n5170 & n5348 ) | ( n5220 & n5348 ) ;
  assign n5351 = ( n5220 & n5349 ) | ( n5220 & ~n5350 ) | ( n5349 & ~n5350 ) ;
  assign n5352 = ( n5212 & n5227 ) | ( n5212 & n5351 ) | ( n5227 & n5351 ) ;
  assign n5353 = ( ~n5212 & n5227 ) | ( ~n5212 & n5351 ) | ( n5227 & n5351 ) ;
  assign n5354 = ( n5212 & ~n5352 ) | ( n5212 & n5353 ) | ( ~n5352 & n5353 ) ;
  assign n5355 = ( n5229 & n5339 ) | ( n5229 & n5354 ) | ( n5339 & n5354 ) ;
  assign n5356 = ( n5229 & ~n5339 ) | ( n5229 & n5354 ) | ( ~n5339 & n5354 ) ;
  assign n5357 = ( n5339 & ~n5355 ) | ( n5339 & n5356 ) | ( ~n5355 & n5356 ) ;
  assign n5358 = ( n5247 & ~n5250 ) | ( n5247 & n5357 ) | ( ~n5250 & n5357 ) ;
  assign n5359 = ( n5247 & n5250 ) | ( n5247 & n5357 ) | ( n5250 & n5357 ) ;
  assign n5360 = ( n5250 & n5358 ) | ( n5250 & ~n5359 ) | ( n5358 & ~n5359 ) ;
  assign n5361 = x12 & x62 ;
  assign n5362 = x13 & x61 ;
  assign n5363 = ( n5295 & n5361 ) | ( n5295 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = ( ~n5295 & n5361 ) | ( ~n5295 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5365 = ( n5295 & ~n5363 ) | ( n5295 & n5364 ) | ( ~n5363 & n5364 ) ;
  assign n5366 = x30 & x44 ;
  assign n5367 = x29 & x45 ;
  assign n5368 = x17 & x57 ;
  assign n5369 = ( ~n5366 & n5367 ) | ( ~n5366 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5370 = ( n5366 & n5367 ) | ( n5366 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5371 = ( n5366 & n5369 ) | ( n5366 & ~n5370 ) | ( n5369 & ~n5370 ) ;
  assign n5372 = ( n5275 & n5365 ) | ( n5275 & n5371 ) | ( n5365 & n5371 ) ;
  assign n5373 = ( n5275 & ~n5365 ) | ( n5275 & n5371 ) | ( ~n5365 & n5371 ) ;
  assign n5374 = ( n5365 & ~n5372 ) | ( n5365 & n5373 ) | ( ~n5372 & n5373 ) ;
  assign n5375 = x19 & x55 ;
  assign n5376 = x22 & x52 ;
  assign n5377 = x21 & x53 ;
  assign n5378 = ( ~n5375 & n5376 ) | ( ~n5375 & n5377 ) | ( n5376 & n5377 ) ;
  assign n5379 = ( n5375 & n5376 ) | ( n5375 & n5377 ) | ( n5376 & n5377 ) ;
  assign n5380 = ( n5375 & n5378 ) | ( n5375 & ~n5379 ) | ( n5378 & ~n5379 ) ;
  assign n5381 = x20 & x54 ;
  assign n5382 = x35 & x39 ;
  assign n5383 = x34 & x40 ;
  assign n5384 = ( ~n5381 & n5382 ) | ( ~n5381 & n5383 ) | ( n5382 & n5383 ) ;
  assign n5385 = ( n5381 & n5382 ) | ( n5381 & n5383 ) | ( n5382 & n5383 ) ;
  assign n5386 = ( n5381 & n5384 ) | ( n5381 & ~n5385 ) | ( n5384 & ~n5385 ) ;
  assign n5387 = x36 & x38 ;
  assign n5388 = x24 & x50 ;
  assign n5389 = x23 & x51 ;
  assign n5390 = ( ~n5387 & n5388 ) | ( ~n5387 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5391 = ( n5387 & n5388 ) | ( n5387 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5392 = ( n5387 & n5390 ) | ( n5387 & ~n5391 ) | ( n5390 & ~n5391 ) ;
  assign n5393 = ( ~n5380 & n5386 ) | ( ~n5380 & n5392 ) | ( n5386 & n5392 ) ;
  assign n5394 = ( n5380 & n5386 ) | ( n5380 & n5392 ) | ( n5386 & n5392 ) ;
  assign n5395 = ( n5380 & n5393 ) | ( n5380 & ~n5394 ) | ( n5393 & ~n5394 ) ;
  assign n5396 = x33 & x41 ;
  assign n5397 = x25 & x49 ;
  assign n5398 = x18 & x56 ;
  assign n5399 = ( ~n5396 & n5397 ) | ( ~n5396 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5400 = ( n5396 & n5397 ) | ( n5396 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5401 = ( n5396 & n5399 ) | ( n5396 & ~n5400 ) | ( n5399 & ~n5400 ) ;
  assign n5402 = x27 & x47 ;
  assign n5403 = x28 & x46 ;
  assign n5404 = x26 & x48 ;
  assign n5405 = ( ~n5402 & n5403 ) | ( ~n5402 & n5404 ) | ( n5403 & n5404 ) ;
  assign n5406 = ( n5402 & n5403 ) | ( n5402 & n5404 ) | ( n5403 & n5404 ) ;
  assign n5407 = ( n5402 & n5405 ) | ( n5402 & ~n5406 ) | ( n5405 & ~n5406 ) ;
  assign n5408 = x11 & x63 ;
  assign n5409 = x32 & x42 ;
  assign n5410 = x31 & x43 ;
  assign n5411 = ( ~n5408 & n5409 ) | ( ~n5408 & n5410 ) | ( n5409 & n5410 ) ;
  assign n5412 = ( n5408 & n5409 ) | ( n5408 & n5410 ) | ( n5409 & n5410 ) ;
  assign n5413 = ( n5408 & n5411 ) | ( n5408 & ~n5412 ) | ( n5411 & ~n5412 ) ;
  assign n5414 = ( ~n5401 & n5407 ) | ( ~n5401 & n5413 ) | ( n5407 & n5413 ) ;
  assign n5415 = ( n5401 & n5407 ) | ( n5401 & n5413 ) | ( n5407 & n5413 ) ;
  assign n5416 = ( n5401 & n5414 ) | ( n5401 & ~n5415 ) | ( n5414 & ~n5415 ) ;
  assign n5417 = ( ~n5374 & n5395 ) | ( ~n5374 & n5416 ) | ( n5395 & n5416 ) ;
  assign n5418 = ( n5374 & n5395 ) | ( n5374 & n5416 ) | ( n5395 & n5416 ) ;
  assign n5419 = ( n5374 & n5417 ) | ( n5374 & ~n5418 ) | ( n5417 & ~n5418 ) ;
  assign n5420 = ( n5257 & n5284 ) | ( n5257 & ~n5290 ) | ( n5284 & ~n5290 ) ;
  assign n5421 = ( n5257 & n5284 ) | ( n5257 & n5290 ) | ( n5284 & n5290 ) ;
  assign n5422 = ( n5290 & n5420 ) | ( n5290 & ~n5421 ) | ( n5420 & ~n5421 ) ;
  assign n5423 = ( n5269 & ~n5304 ) | ( n5269 & n5310 ) | ( ~n5304 & n5310 ) ;
  assign n5424 = ( n5269 & n5304 ) | ( n5269 & n5310 ) | ( n5304 & n5310 ) ;
  assign n5425 = ( n5304 & n5423 ) | ( n5304 & ~n5424 ) | ( n5423 & ~n5424 ) ;
  assign n5426 = ( n5272 & n5422 ) | ( n5272 & n5425 ) | ( n5422 & n5425 ) ;
  assign n5427 = ( n5272 & ~n5422 ) | ( n5272 & n5425 ) | ( ~n5422 & n5425 ) ;
  assign n5428 = ( n5422 & ~n5426 ) | ( n5422 & n5427 ) | ( ~n5426 & n5427 ) ;
  assign n5429 = ( n5350 & n5419 ) | ( n5350 & n5428 ) | ( n5419 & n5428 ) ;
  assign n5430 = ( ~n5350 & n5419 ) | ( ~n5350 & n5428 ) | ( n5419 & n5428 ) ;
  assign n5431 = ( n5350 & ~n5429 ) | ( n5350 & n5430 ) | ( ~n5429 & n5430 ) ;
  assign n5432 = x16 & x58 ;
  assign n5433 = x14 & x60 ;
  assign n5434 = x15 & x59 ;
  assign n5435 = ( ~n5432 & n5433 ) | ( ~n5432 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = ( n5432 & n5433 ) | ( n5432 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5437 = ( n5432 & n5435 ) | ( n5432 & ~n5436 ) | ( n5435 & ~n5436 ) ;
  assign n5438 = ( n5263 & n5344 ) | ( n5263 & ~n5437 ) | ( n5344 & ~n5437 ) ;
  assign n5439 = ( n5263 & n5344 ) | ( n5263 & n5437 ) | ( n5344 & n5437 ) ;
  assign n5440 = ( n5437 & n5438 ) | ( n5437 & ~n5439 ) | ( n5438 & ~n5439 ) ;
  assign n5441 = ( n5298 & n5347 ) | ( n5298 & n5440 ) | ( n5347 & n5440 ) ;
  assign n5442 = ( n5298 & ~n5347 ) | ( n5298 & n5440 ) | ( ~n5347 & n5440 ) ;
  assign n5443 = ( n5347 & ~n5441 ) | ( n5347 & n5442 ) | ( ~n5441 & n5442 ) ;
  assign n5444 = ( n5277 & n5315 ) | ( n5277 & n5443 ) | ( n5315 & n5443 ) ;
  assign n5445 = ( n5277 & ~n5315 ) | ( n5277 & n5443 ) | ( ~n5315 & n5443 ) ;
  assign n5446 = ( n5315 & ~n5444 ) | ( n5315 & n5445 ) | ( ~n5444 & n5445 ) ;
  assign n5447 = ( n5352 & n5431 ) | ( n5352 & n5446 ) | ( n5431 & n5446 ) ;
  assign n5448 = ( ~n5352 & n5431 ) | ( ~n5352 & n5446 ) | ( n5431 & n5446 ) ;
  assign n5449 = ( n5352 & ~n5447 ) | ( n5352 & n5448 ) | ( ~n5447 & n5448 ) ;
  assign n5450 = ( ~n5313 & n5325 ) | ( ~n5313 & n5328 ) | ( n5325 & n5328 ) ;
  assign n5451 = ( n5313 & n5325 ) | ( n5313 & n5328 ) | ( n5325 & n5328 ) ;
  assign n5452 = ( n5313 & n5450 ) | ( n5313 & ~n5451 ) | ( n5450 & ~n5451 ) ;
  assign n5453 = ( n5322 & n5331 ) | ( n5322 & n5452 ) | ( n5331 & n5452 ) ;
  assign n5454 = ( n5322 & n5331 ) | ( n5322 & ~n5452 ) | ( n5331 & ~n5452 ) ;
  assign n5455 = ( n5452 & ~n5453 ) | ( n5452 & n5454 ) | ( ~n5453 & n5454 ) ;
  assign n5456 = ( n5319 & n5335 ) | ( n5319 & n5455 ) | ( n5335 & n5455 ) ;
  assign n5457 = ( ~n5319 & n5335 ) | ( ~n5319 & n5455 ) | ( n5335 & n5455 ) ;
  assign n5458 = ( n5319 & ~n5456 ) | ( n5319 & n5457 ) | ( ~n5456 & n5457 ) ;
  assign n5459 = ( n5337 & n5449 ) | ( n5337 & n5458 ) | ( n5449 & n5458 ) ;
  assign n5460 = ( n5337 & ~n5449 ) | ( n5337 & n5458 ) | ( ~n5449 & n5458 ) ;
  assign n5461 = ( n5449 & ~n5459 ) | ( n5449 & n5460 ) | ( ~n5459 & n5460 ) ;
  assign n5462 = ( n5355 & n5359 ) | ( n5355 & n5461 ) | ( n5359 & n5461 ) ;
  assign n5463 = ( n5355 & n5359 ) | ( n5355 & ~n5461 ) | ( n5359 & ~n5461 ) ;
  assign n5464 = ( n5461 & ~n5462 ) | ( n5461 & n5463 ) | ( ~n5462 & n5463 ) ;
  assign n5465 = x16 & x59 ;
  assign n5466 = x14 & x61 ;
  assign n5467 = x15 & x60 ;
  assign n5468 = ( ~n5465 & n5466 ) | ( ~n5465 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5469 = ( n5465 & n5466 ) | ( n5465 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5470 = ( n5465 & n5468 ) | ( n5465 & ~n5469 ) | ( n5468 & ~n5469 ) ;
  assign n5471 = x27 & x48 ;
  assign n5472 = x28 & x47 ;
  assign n5473 = x29 & x46 ;
  assign n5474 = ( ~n5471 & n5472 ) | ( ~n5471 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5475 = ( n5471 & n5472 ) | ( n5471 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5476 = ( n5471 & n5474 ) | ( n5471 & ~n5475 ) | ( n5474 & ~n5475 ) ;
  assign n5477 = x17 & x58 ;
  assign n5478 = x18 & x57 ;
  assign n5479 = ( ~n2598 & n5477 ) | ( ~n2598 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5480 = ( n2598 & n5477 ) | ( n2598 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5481 = ( n2598 & n5479 ) | ( n2598 & ~n5480 ) | ( n5479 & ~n5480 ) ;
  assign n5482 = ( ~n5470 & n5476 ) | ( ~n5470 & n5481 ) | ( n5476 & n5481 ) ;
  assign n5483 = ( n5470 & n5476 ) | ( n5470 & n5481 ) | ( n5476 & n5481 ) ;
  assign n5484 = ( n5470 & n5482 ) | ( n5470 & ~n5483 ) | ( n5482 & ~n5483 ) ;
  assign n5485 = x12 & x63 ;
  assign n5486 = x30 & x45 ;
  assign n5487 = x19 & x56 ;
  assign n5488 = ( ~n5485 & n5486 ) | ( ~n5485 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5489 = ( n5485 & n5486 ) | ( n5485 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5490 = ( n5485 & n5488 ) | ( n5485 & ~n5489 ) | ( n5488 & ~n5489 ) ;
  assign n5491 = x35 & x40 ;
  assign n5492 = x36 & x39 ;
  assign n5493 = x23 & x52 ;
  assign n5494 = ( ~n5491 & n5492 ) | ( ~n5491 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5495 = ( n5491 & n5492 ) | ( n5491 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5496 = ( n5491 & n5494 ) | ( n5491 & ~n5495 ) | ( n5494 & ~n5495 ) ;
  assign n5497 = x13 & x62 ;
  assign n5498 = x37 & x38 ;
  assign n5499 = ( x38 & n5497 ) | ( x38 & n5498 ) | ( n5497 & n5498 ) ;
  assign n5500 = ( x38 & ~n5497 ) | ( x38 & n5498 ) | ( ~n5497 & n5498 ) ;
  assign n5501 = ( n5497 & ~n5499 ) | ( n5497 & n5500 ) | ( ~n5499 & n5500 ) ;
  assign n5502 = ( ~n5490 & n5496 ) | ( ~n5490 & n5501 ) | ( n5496 & n5501 ) ;
  assign n5503 = ( n5490 & n5496 ) | ( n5490 & n5501 ) | ( n5496 & n5501 ) ;
  assign n5504 = ( n5490 & n5502 ) | ( n5490 & ~n5503 ) | ( n5502 & ~n5503 ) ;
  assign n5505 = ( ~n5451 & n5484 ) | ( ~n5451 & n5504 ) | ( n5484 & n5504 ) ;
  assign n5506 = ( n5451 & n5484 ) | ( n5451 & n5504 ) | ( n5484 & n5504 ) ;
  assign n5507 = ( n5451 & n5505 ) | ( n5451 & ~n5506 ) | ( n5505 & ~n5506 ) ;
  assign n5508 = ( n5370 & n5406 ) | ( n5370 & ~n5436 ) | ( n5406 & ~n5436 ) ;
  assign n5509 = ( n5370 & n5406 ) | ( n5370 & n5436 ) | ( n5406 & n5436 ) ;
  assign n5510 = ( n5436 & n5508 ) | ( n5436 & ~n5509 ) | ( n5508 & ~n5509 ) ;
  assign n5511 = ( n5394 & n5415 ) | ( n5394 & n5510 ) | ( n5415 & n5510 ) ;
  assign n5512 = ( n5394 & n5415 ) | ( n5394 & ~n5510 ) | ( n5415 & ~n5510 ) ;
  assign n5513 = ( n5510 & ~n5511 ) | ( n5510 & n5512 ) | ( ~n5511 & n5512 ) ;
  assign n5514 = ( n5453 & n5507 ) | ( n5453 & n5513 ) | ( n5507 & n5513 ) ;
  assign n5515 = ( ~n5453 & n5507 ) | ( ~n5453 & n5513 ) | ( n5507 & n5513 ) ;
  assign n5516 = ( n5453 & ~n5514 ) | ( n5453 & n5515 ) | ( ~n5514 & n5515 ) ;
  assign n5517 = ( n5421 & n5424 ) | ( n5421 & ~n5439 ) | ( n5424 & ~n5439 ) ;
  assign n5518 = ( n5421 & n5424 ) | ( n5421 & n5439 ) | ( n5424 & n5439 ) ;
  assign n5519 = ( n5439 & n5517 ) | ( n5439 & ~n5518 ) | ( n5517 & ~n5518 ) ;
  assign n5520 = ( ~n5363 & n5400 ) | ( ~n5363 & n5412 ) | ( n5400 & n5412 ) ;
  assign n5521 = ( n5363 & n5400 ) | ( n5363 & n5412 ) | ( n5400 & n5412 ) ;
  assign n5522 = ( n5363 & n5520 ) | ( n5363 & ~n5521 ) | ( n5520 & ~n5521 ) ;
  assign n5523 = ( n5379 & ~n5385 ) | ( n5379 & n5391 ) | ( ~n5385 & n5391 ) ;
  assign n5524 = ( n5379 & n5385 ) | ( n5379 & n5391 ) | ( n5385 & n5391 ) ;
  assign n5525 = ( n5385 & n5523 ) | ( n5385 & ~n5524 ) | ( n5523 & ~n5524 ) ;
  assign n5526 = ( n5372 & n5522 ) | ( n5372 & n5525 ) | ( n5522 & n5525 ) ;
  assign n5527 = ( ~n5372 & n5522 ) | ( ~n5372 & n5525 ) | ( n5522 & n5525 ) ;
  assign n5528 = ( n5372 & ~n5526 ) | ( n5372 & n5527 ) | ( ~n5526 & n5527 ) ;
  assign n5529 = ( n5418 & n5519 ) | ( n5418 & n5528 ) | ( n5519 & n5528 ) ;
  assign n5530 = ( ~n5418 & n5519 ) | ( ~n5418 & n5528 ) | ( n5519 & n5528 ) ;
  assign n5531 = ( n5418 & ~n5529 ) | ( n5418 & n5530 ) | ( ~n5529 & n5530 ) ;
  assign n5532 = ( n5456 & ~n5516 ) | ( n5456 & n5531 ) | ( ~n5516 & n5531 ) ;
  assign n5533 = ( n5456 & n5516 ) | ( n5456 & n5531 ) | ( n5516 & n5531 ) ;
  assign n5534 = ( n5516 & n5532 ) | ( n5516 & ~n5533 ) | ( n5532 & ~n5533 ) ;
  assign n5535 = x21 & x54 ;
  assign n5536 = x24 & x51 ;
  assign n5537 = x22 & x53 ;
  assign n5538 = ( ~n5535 & n5536 ) | ( ~n5535 & n5537 ) | ( n5536 & n5537 ) ;
  assign n5539 = ( n5535 & n5536 ) | ( n5535 & n5537 ) | ( n5536 & n5537 ) ;
  assign n5540 = ( n5535 & n5538 ) | ( n5535 & ~n5539 ) | ( n5538 & ~n5539 ) ;
  assign n5541 = x31 & x44 ;
  assign n5542 = x32 & x43 ;
  assign n5543 = x33 & x42 ;
  assign n5544 = ( ~n5541 & n5542 ) | ( ~n5541 & n5543 ) | ( n5542 & n5543 ) ;
  assign n5545 = ( n5541 & n5542 ) | ( n5541 & n5543 ) | ( n5542 & n5543 ) ;
  assign n5546 = ( n5541 & n5544 ) | ( n5541 & ~n5545 ) | ( n5544 & ~n5545 ) ;
  assign n5547 = x34 & x41 ;
  assign n5548 = x25 & x50 ;
  assign n5549 = x20 & x55 ;
  assign n5550 = ( ~n5547 & n5548 ) | ( ~n5547 & n5549 ) | ( n5548 & n5549 ) ;
  assign n5551 = ( n5547 & n5548 ) | ( n5547 & n5549 ) | ( n5548 & n5549 ) ;
  assign n5552 = ( n5547 & n5550 ) | ( n5547 & ~n5551 ) | ( n5550 & ~n5551 ) ;
  assign n5553 = ( ~n5540 & n5546 ) | ( ~n5540 & n5552 ) | ( n5546 & n5552 ) ;
  assign n5554 = ( n5540 & n5546 ) | ( n5540 & n5552 ) | ( n5546 & n5552 ) ;
  assign n5555 = ( n5540 & n5553 ) | ( n5540 & ~n5554 ) | ( n5553 & ~n5554 ) ;
  assign n5556 = ( n5426 & n5441 ) | ( n5426 & n5555 ) | ( n5441 & n5555 ) ;
  assign n5557 = ( n5426 & ~n5441 ) | ( n5426 & n5555 ) | ( ~n5441 & n5555 ) ;
  assign n5558 = ( n5441 & ~n5556 ) | ( n5441 & n5557 ) | ( ~n5556 & n5557 ) ;
  assign n5559 = ( n5429 & n5444 ) | ( n5429 & n5558 ) | ( n5444 & n5558 ) ;
  assign n5560 = ( ~n5429 & n5444 ) | ( ~n5429 & n5558 ) | ( n5444 & n5558 ) ;
  assign n5561 = ( n5429 & ~n5559 ) | ( n5429 & n5560 ) | ( ~n5559 & n5560 ) ;
  assign n5562 = ( ~n5447 & n5534 ) | ( ~n5447 & n5561 ) | ( n5534 & n5561 ) ;
  assign n5563 = ( n5447 & n5534 ) | ( n5447 & n5561 ) | ( n5534 & n5561 ) ;
  assign n5564 = ( n5447 & n5562 ) | ( n5447 & ~n5563 ) | ( n5562 & ~n5563 ) ;
  assign n5565 = ( n5459 & ~n5462 ) | ( n5459 & n5564 ) | ( ~n5462 & n5564 ) ;
  assign n5566 = ( n5459 & n5462 ) | ( n5459 & n5564 ) | ( n5462 & n5564 ) ;
  assign n5567 = ( n5462 & n5565 ) | ( n5462 & ~n5566 ) | ( n5565 & ~n5566 ) ;
  assign n5568 = ( n5475 & n5489 ) | ( n5475 & ~n5551 ) | ( n5489 & ~n5551 ) ;
  assign n5569 = ( n5475 & n5489 ) | ( n5475 & n5551 ) | ( n5489 & n5551 ) ;
  assign n5570 = ( n5551 & n5568 ) | ( n5551 & ~n5569 ) | ( n5568 & ~n5569 ) ;
  assign n5571 = x14 & x62 ;
  assign n5572 = ( n5495 & n5499 ) | ( n5495 & n5571 ) | ( n5499 & n5571 ) ;
  assign n5573 = ( ~n5495 & n5499 ) | ( ~n5495 & n5571 ) | ( n5499 & n5571 ) ;
  assign n5574 = ( n5495 & ~n5572 ) | ( n5495 & n5573 ) | ( ~n5572 & n5573 ) ;
  assign n5575 = ( n5554 & n5570 ) | ( n5554 & n5574 ) | ( n5570 & n5574 ) ;
  assign n5576 = ( n5554 & ~n5570 ) | ( n5554 & n5574 ) | ( ~n5570 & n5574 ) ;
  assign n5577 = ( n5570 & ~n5575 ) | ( n5570 & n5576 ) | ( ~n5575 & n5576 ) ;
  assign n5578 = ( n5509 & ~n5521 ) | ( n5509 & n5524 ) | ( ~n5521 & n5524 ) ;
  assign n5579 = ( n5509 & n5521 ) | ( n5509 & n5524 ) | ( n5521 & n5524 ) ;
  assign n5580 = ( n5521 & n5578 ) | ( n5521 & ~n5579 ) | ( n5578 & ~n5579 ) ;
  assign n5581 = ( n5506 & ~n5577 ) | ( n5506 & n5580 ) | ( ~n5577 & n5580 ) ;
  assign n5582 = ( n5506 & n5577 ) | ( n5506 & n5580 ) | ( n5577 & n5580 ) ;
  assign n5583 = ( n5577 & n5581 ) | ( n5577 & ~n5582 ) | ( n5581 & ~n5582 ) ;
  assign n5584 = x15 & x61 ;
  assign n5585 = x16 & x60 ;
  assign n5586 = x17 & x59 ;
  assign n5587 = ( ~n5584 & n5585 ) | ( ~n5584 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5588 = ( n5584 & n5585 ) | ( n5584 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5589 = ( n5584 & n5587 ) | ( n5584 & ~n5588 ) | ( n5587 & ~n5588 ) ;
  assign n5590 = x27 & x49 ;
  assign n5591 = x18 & x58 ;
  assign n5592 = ( ~n2731 & n5590 ) | ( ~n2731 & n5591 ) | ( n5590 & n5591 ) ;
  assign n5593 = ( n2731 & n5590 ) | ( n2731 & n5591 ) | ( n5590 & n5591 ) ;
  assign n5594 = ( n2731 & n5592 ) | ( n2731 & ~n5593 ) | ( n5592 & ~n5593 ) ;
  assign n5595 = ( ~n5539 & n5589 ) | ( ~n5539 & n5594 ) | ( n5589 & n5594 ) ;
  assign n5596 = ( n5539 & n5589 ) | ( n5539 & n5594 ) | ( n5589 & n5594 ) ;
  assign n5597 = ( n5539 & n5595 ) | ( n5539 & ~n5596 ) | ( n5595 & ~n5596 ) ;
  assign n5598 = x36 & x40 ;
  assign n5599 = x34 & x42 ;
  assign n5600 = x35 & x41 ;
  assign n5601 = ( ~n5598 & n5599 ) | ( ~n5598 & n5600 ) | ( n5599 & n5600 ) ;
  assign n5602 = ( n5598 & n5599 ) | ( n5598 & n5600 ) | ( n5599 & n5600 ) ;
  assign n5603 = ( n5598 & n5601 ) | ( n5598 & ~n5602 ) | ( n5601 & ~n5602 ) ;
  assign n5604 = x30 & x46 ;
  assign n5605 = x29 & x47 ;
  assign n5606 = x28 & x48 ;
  assign n5607 = ( ~n5604 & n5605 ) | ( ~n5604 & n5606 ) | ( n5605 & n5606 ) ;
  assign n5608 = ( n5604 & n5605 ) | ( n5604 & n5606 ) | ( n5605 & n5606 ) ;
  assign n5609 = ( n5604 & n5607 ) | ( n5604 & ~n5608 ) | ( n5607 & ~n5608 ) ;
  assign n5610 = x37 & x39 ;
  assign n5611 = x25 & x51 ;
  assign n5612 = x24 & x52 ;
  assign n5613 = ( ~n5610 & n5611 ) | ( ~n5610 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5614 = ( n5610 & n5611 ) | ( n5610 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5615 = ( n5610 & n5613 ) | ( n5610 & ~n5614 ) | ( n5613 & ~n5614 ) ;
  assign n5616 = ( ~n5603 & n5609 ) | ( ~n5603 & n5615 ) | ( n5609 & n5615 ) ;
  assign n5617 = ( n5603 & n5609 ) | ( n5603 & n5615 ) | ( n5609 & n5615 ) ;
  assign n5618 = ( n5603 & n5616 ) | ( n5603 & ~n5617 ) | ( n5616 & ~n5617 ) ;
  assign n5619 = ( n5518 & n5597 ) | ( n5518 & n5618 ) | ( n5597 & n5618 ) ;
  assign n5620 = ( ~n5518 & n5597 ) | ( ~n5518 & n5618 ) | ( n5597 & n5618 ) ;
  assign n5621 = ( n5518 & ~n5619 ) | ( n5518 & n5620 ) | ( ~n5619 & n5620 ) ;
  assign n5622 = ( n5469 & n5480 ) | ( n5469 & ~n5545 ) | ( n5480 & ~n5545 ) ;
  assign n5623 = ( n5469 & n5480 ) | ( n5469 & n5545 ) | ( n5480 & n5545 ) ;
  assign n5624 = ( n5545 & n5622 ) | ( n5545 & ~n5623 ) | ( n5622 & ~n5623 ) ;
  assign n5625 = ( n5483 & n5503 ) | ( n5483 & n5624 ) | ( n5503 & n5624 ) ;
  assign n5626 = ( n5483 & n5503 ) | ( n5483 & ~n5624 ) | ( n5503 & ~n5624 ) ;
  assign n5627 = ( n5624 & ~n5625 ) | ( n5624 & n5626 ) | ( ~n5625 & n5626 ) ;
  assign n5628 = ( n5556 & n5621 ) | ( n5556 & n5627 ) | ( n5621 & n5627 ) ;
  assign n5629 = ( ~n5556 & n5621 ) | ( ~n5556 & n5627 ) | ( n5621 & n5627 ) ;
  assign n5630 = ( n5556 & ~n5628 ) | ( n5556 & n5629 ) | ( ~n5628 & n5629 ) ;
  assign n5631 = ( n5559 & n5583 ) | ( n5559 & n5630 ) | ( n5583 & n5630 ) ;
  assign n5632 = ( ~n5559 & n5583 ) | ( ~n5559 & n5630 ) | ( n5583 & n5630 ) ;
  assign n5633 = ( n5559 & ~n5631 ) | ( n5559 & n5632 ) | ( ~n5631 & n5632 ) ;
  assign n5634 = x13 & x63 ;
  assign n5635 = x32 & x44 ;
  assign n5636 = x31 & x45 ;
  assign n5637 = ( ~n5634 & n5635 ) | ( ~n5634 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5638 = ( n5634 & n5635 ) | ( n5634 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5639 = ( n5634 & n5637 ) | ( n5634 & ~n5638 ) | ( n5637 & ~n5638 ) ;
  assign n5640 = x20 & x56 ;
  assign n5641 = x22 & x54 ;
  assign n5642 = x21 & x55 ;
  assign n5643 = ( ~n5640 & n5641 ) | ( ~n5640 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5644 = ( n5640 & n5641 ) | ( n5640 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5645 = ( n5640 & n5643 ) | ( n5640 & ~n5644 ) | ( n5643 & ~n5644 ) ;
  assign n5646 = x33 & x43 ;
  assign n5647 = x23 & x53 ;
  assign n5648 = x19 & x57 ;
  assign n5649 = ( ~n5646 & n5647 ) | ( ~n5646 & n5648 ) | ( n5647 & n5648 ) ;
  assign n5650 = ( n5646 & n5647 ) | ( n5646 & n5648 ) | ( n5647 & n5648 ) ;
  assign n5651 = ( n5646 & n5649 ) | ( n5646 & ~n5650 ) | ( n5649 & ~n5650 ) ;
  assign n5652 = ( ~n5639 & n5645 ) | ( ~n5639 & n5651 ) | ( n5645 & n5651 ) ;
  assign n5653 = ( n5639 & n5645 ) | ( n5639 & n5651 ) | ( n5645 & n5651 ) ;
  assign n5654 = ( n5639 & n5652 ) | ( n5639 & ~n5653 ) | ( n5652 & ~n5653 ) ;
  assign n5655 = ( n5511 & n5526 ) | ( n5511 & n5654 ) | ( n5526 & n5654 ) ;
  assign n5656 = ( n5511 & ~n5526 ) | ( n5511 & n5654 ) | ( ~n5526 & n5654 ) ;
  assign n5657 = ( n5526 & ~n5655 ) | ( n5526 & n5656 ) | ( ~n5655 & n5656 ) ;
  assign n5658 = ( n5514 & n5529 ) | ( n5514 & n5657 ) | ( n5529 & n5657 ) ;
  assign n5659 = ( ~n5514 & n5529 ) | ( ~n5514 & n5657 ) | ( n5529 & n5657 ) ;
  assign n5660 = ( n5514 & ~n5658 ) | ( n5514 & n5659 ) | ( ~n5658 & n5659 ) ;
  assign n5661 = ( n5533 & n5633 ) | ( n5533 & n5660 ) | ( n5633 & n5660 ) ;
  assign n5662 = ( n5533 & ~n5633 ) | ( n5533 & n5660 ) | ( ~n5633 & n5660 ) ;
  assign n5663 = ( n5633 & ~n5661 ) | ( n5633 & n5662 ) | ( ~n5661 & n5662 ) ;
  assign n5664 = ( n5563 & n5566 ) | ( n5563 & n5663 ) | ( n5566 & n5663 ) ;
  assign n5665 = ( n5563 & ~n5566 ) | ( n5563 & n5663 ) | ( ~n5566 & n5663 ) ;
  assign n5666 = ( n5566 & ~n5664 ) | ( n5566 & n5665 ) | ( ~n5664 & n5665 ) ;
  assign n5667 = x17 & x60 ;
  assign n5668 = x18 & x59 ;
  assign n5669 = ( n5614 & n5667 ) | ( n5614 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5670 = ( ~n5614 & n5667 ) | ( ~n5614 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5671 = ( n5614 & ~n5669 ) | ( n5614 & n5670 ) | ( ~n5669 & n5670 ) ;
  assign n5672 = ( n5569 & n5623 ) | ( n5569 & n5671 ) | ( n5623 & n5671 ) ;
  assign n5673 = ( n5569 & n5623 ) | ( n5569 & ~n5671 ) | ( n5623 & ~n5671 ) ;
  assign n5674 = ( n5671 & ~n5672 ) | ( n5671 & n5673 ) | ( ~n5672 & n5673 ) ;
  assign n5675 = ( n5608 & ~n5638 ) | ( n5608 & n5644 ) | ( ~n5638 & n5644 ) ;
  assign n5676 = ( n5608 & n5638 ) | ( n5608 & n5644 ) | ( n5638 & n5644 ) ;
  assign n5677 = ( n5638 & n5675 ) | ( n5638 & ~n5676 ) | ( n5675 & ~n5676 ) ;
  assign n5678 = ( ~n5588 & n5593 ) | ( ~n5588 & n5650 ) | ( n5593 & n5650 ) ;
  assign n5679 = ( n5588 & n5593 ) | ( n5588 & n5650 ) | ( n5593 & n5650 ) ;
  assign n5680 = ( n5588 & n5678 ) | ( n5588 & ~n5679 ) | ( n5678 & ~n5679 ) ;
  assign n5681 = ( n5653 & n5677 ) | ( n5653 & n5680 ) | ( n5677 & n5680 ) ;
  assign n5682 = ( n5653 & ~n5677 ) | ( n5653 & n5680 ) | ( ~n5677 & n5680 ) ;
  assign n5683 = ( n5677 & ~n5681 ) | ( n5677 & n5682 ) | ( ~n5681 & n5682 ) ;
  assign n5684 = ( ~n5619 & n5674 ) | ( ~n5619 & n5683 ) | ( n5674 & n5683 ) ;
  assign n5685 = ( n5619 & n5674 ) | ( n5619 & n5683 ) | ( n5674 & n5683 ) ;
  assign n5686 = ( n5619 & n5684 ) | ( n5619 & ~n5685 ) | ( n5684 & ~n5685 ) ;
  assign n5687 = x15 & x62 ;
  assign n5688 = x38 & x39 ;
  assign n5689 = ( x39 & n5687 ) | ( x39 & n5688 ) | ( n5687 & n5688 ) ;
  assign n5690 = ( x39 & ~n5687 ) | ( x39 & n5688 ) | ( ~n5687 & n5688 ) ;
  assign n5691 = ( n5687 & ~n5689 ) | ( n5687 & n5690 ) | ( ~n5689 & n5690 ) ;
  assign n5692 = x14 & x63 ;
  assign n5693 = x30 & x47 ;
  assign n5694 = x31 & x46 ;
  assign n5695 = ( ~n5692 & n5693 ) | ( ~n5692 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5696 = ( n5692 & n5693 ) | ( n5692 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5697 = ( n5692 & n5695 ) | ( n5692 & ~n5696 ) | ( n5695 & ~n5696 ) ;
  assign n5698 = x35 & x42 ;
  assign n5699 = x37 & x40 ;
  assign n5700 = x36 & x41 ;
  assign n5701 = ( ~n5698 & n5699 ) | ( ~n5698 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5702 = ( n5698 & n5699 ) | ( n5698 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5703 = ( n5698 & n5701 ) | ( n5698 & ~n5702 ) | ( n5701 & ~n5702 ) ;
  assign n5704 = ( ~n5691 & n5697 ) | ( ~n5691 & n5703 ) | ( n5697 & n5703 ) ;
  assign n5705 = ( n5691 & n5697 ) | ( n5691 & n5703 ) | ( n5697 & n5703 ) ;
  assign n5706 = ( n5691 & n5704 ) | ( n5691 & ~n5705 ) | ( n5704 & ~n5705 ) ;
  assign n5707 = x20 & x57 ;
  assign n5708 = x21 & x56 ;
  assign n5709 = x19 & x58 ;
  assign n5710 = ( ~n5707 & n5708 ) | ( ~n5707 & n5709 ) | ( n5708 & n5709 ) ;
  assign n5711 = ( n5707 & n5708 ) | ( n5707 & n5709 ) | ( n5708 & n5709 ) ;
  assign n5712 = ( n5707 & n5710 ) | ( n5707 & ~n5711 ) | ( n5710 & ~n5711 ) ;
  assign n5713 = x29 & x48 ;
  assign n5714 = x27 & x50 ;
  assign n5715 = x28 & x49 ;
  assign n5716 = ( ~n5713 & n5714 ) | ( ~n5713 & n5715 ) | ( n5714 & n5715 ) ;
  assign n5717 = ( n5713 & n5714 ) | ( n5713 & n5715 ) | ( n5714 & n5715 ) ;
  assign n5718 = ( n5713 & n5716 ) | ( n5713 & ~n5717 ) | ( n5716 & ~n5717 ) ;
  assign n5719 = ( ~n5602 & n5712 ) | ( ~n5602 & n5718 ) | ( n5712 & n5718 ) ;
  assign n5720 = ( n5602 & n5712 ) | ( n5602 & n5718 ) | ( n5712 & n5718 ) ;
  assign n5721 = ( n5602 & n5719 ) | ( n5602 & ~n5720 ) | ( n5719 & ~n5720 ) ;
  assign n5722 = ( n5579 & n5706 ) | ( n5579 & n5721 ) | ( n5706 & n5721 ) ;
  assign n5723 = ( ~n5579 & n5706 ) | ( ~n5579 & n5721 ) | ( n5706 & n5721 ) ;
  assign n5724 = ( n5579 & ~n5722 ) | ( n5579 & n5723 ) | ( ~n5722 & n5723 ) ;
  assign n5725 = ( ~n5572 & n5596 ) | ( ~n5572 & n5617 ) | ( n5596 & n5617 ) ;
  assign n5726 = ( n5572 & n5596 ) | ( n5572 & n5617 ) | ( n5596 & n5617 ) ;
  assign n5727 = ( n5572 & n5725 ) | ( n5572 & ~n5726 ) | ( n5725 & ~n5726 ) ;
  assign n5728 = ( n5655 & n5724 ) | ( n5655 & n5727 ) | ( n5724 & n5727 ) ;
  assign n5729 = ( ~n5655 & n5724 ) | ( ~n5655 & n5727 ) | ( n5724 & n5727 ) ;
  assign n5730 = ( n5655 & ~n5728 ) | ( n5655 & n5729 ) | ( ~n5728 & n5729 ) ;
  assign n5731 = ( n5658 & n5686 ) | ( n5658 & n5730 ) | ( n5686 & n5730 ) ;
  assign n5732 = ( ~n5658 & n5686 ) | ( ~n5658 & n5730 ) | ( n5686 & n5730 ) ;
  assign n5733 = ( n5658 & ~n5731 ) | ( n5658 & n5732 ) | ( ~n5731 & n5732 ) ;
  assign n5734 = x32 & x45 ;
  assign n5735 = x16 & x61 ;
  assign n5736 = x33 & x44 ;
  assign n5737 = ( ~n5734 & n5735 ) | ( ~n5734 & n5736 ) | ( n5735 & n5736 ) ;
  assign n5738 = ( n5734 & n5735 ) | ( n5734 & n5736 ) | ( n5735 & n5736 ) ;
  assign n5739 = ( n5734 & n5737 ) | ( n5734 & ~n5738 ) | ( n5737 & ~n5738 ) ;
  assign n5740 = x22 & x55 ;
  assign n5741 = x34 & x43 ;
  assign n5742 = x26 & x51 ;
  assign n5743 = ( ~n5740 & n5741 ) | ( ~n5740 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5744 = ( n5740 & n5741 ) | ( n5740 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5745 = ( n5740 & n5743 ) | ( n5740 & ~n5744 ) | ( n5743 & ~n5744 ) ;
  assign n5746 = x23 & x54 ;
  assign n5747 = x25 & x52 ;
  assign n5748 = x24 & x53 ;
  assign n5749 = ( ~n5746 & n5747 ) | ( ~n5746 & n5748 ) | ( n5747 & n5748 ) ;
  assign n5750 = ( n5746 & n5747 ) | ( n5746 & n5748 ) | ( n5747 & n5748 ) ;
  assign n5751 = ( n5746 & n5749 ) | ( n5746 & ~n5750 ) | ( n5749 & ~n5750 ) ;
  assign n5752 = ( ~n5739 & n5745 ) | ( ~n5739 & n5751 ) | ( n5745 & n5751 ) ;
  assign n5753 = ( n5739 & n5745 ) | ( n5739 & n5751 ) | ( n5745 & n5751 ) ;
  assign n5754 = ( n5739 & n5752 ) | ( n5739 & ~n5753 ) | ( n5752 & ~n5753 ) ;
  assign n5755 = ( n5575 & n5625 ) | ( n5575 & n5754 ) | ( n5625 & n5754 ) ;
  assign n5756 = ( n5575 & ~n5625 ) | ( n5575 & n5754 ) | ( ~n5625 & n5754 ) ;
  assign n5757 = ( n5625 & ~n5755 ) | ( n5625 & n5756 ) | ( ~n5755 & n5756 ) ;
  assign n5758 = ( n5582 & n5628 ) | ( n5582 & n5757 ) | ( n5628 & n5757 ) ;
  assign n5759 = ( n5582 & ~n5628 ) | ( n5582 & n5757 ) | ( ~n5628 & n5757 ) ;
  assign n5760 = ( n5628 & ~n5758 ) | ( n5628 & n5759 ) | ( ~n5758 & n5759 ) ;
  assign n5761 = ( n5631 & n5733 ) | ( n5631 & n5760 ) | ( n5733 & n5760 ) ;
  assign n5762 = ( ~n5631 & n5733 ) | ( ~n5631 & n5760 ) | ( n5733 & n5760 ) ;
  assign n5763 = ( n5631 & ~n5761 ) | ( n5631 & n5762 ) | ( ~n5761 & n5762 ) ;
  assign n5764 = ( n5661 & n5664 ) | ( n5661 & n5763 ) | ( n5664 & n5763 ) ;
  assign n5765 = ( n5661 & ~n5664 ) | ( n5661 & n5763 ) | ( ~n5664 & n5763 ) ;
  assign n5766 = ( n5664 & ~n5764 ) | ( n5664 & n5765 ) | ( ~n5764 & n5765 ) ;
  assign n5767 = ( ~n5669 & n5711 ) | ( ~n5669 & n5744 ) | ( n5711 & n5744 ) ;
  assign n5768 = ( n5669 & n5711 ) | ( n5669 & n5744 ) | ( n5711 & n5744 ) ;
  assign n5769 = ( n5669 & n5767 ) | ( n5669 & ~n5768 ) | ( n5767 & ~n5768 ) ;
  assign n5770 = x35 & x43 ;
  assign n5771 = x36 & x42 ;
  assign n5772 = x23 & x55 ;
  assign n5773 = ( ~n5770 & n5771 ) | ( ~n5770 & n5772 ) | ( n5771 & n5772 ) ;
  assign n5774 = ( n5770 & n5771 ) | ( n5770 & n5772 ) | ( n5771 & n5772 ) ;
  assign n5775 = ( n5770 & n5773 ) | ( n5770 & ~n5774 ) | ( n5773 & ~n5774 ) ;
  assign n5776 = x38 & x40 ;
  assign n5777 = x26 & x52 ;
  assign n5778 = x37 & x41 ;
  assign n5779 = ( ~n5776 & n5777 ) | ( ~n5776 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = ( n5776 & n5777 ) | ( n5776 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5781 = ( n5776 & n5779 ) | ( n5776 & ~n5780 ) | ( n5779 & ~n5780 ) ;
  assign n5782 = ( ~n5676 & n5775 ) | ( ~n5676 & n5781 ) | ( n5775 & n5781 ) ;
  assign n5783 = ( n5676 & n5775 ) | ( n5676 & n5781 ) | ( n5775 & n5781 ) ;
  assign n5784 = ( n5676 & n5782 ) | ( n5676 & ~n5783 ) | ( n5782 & ~n5783 ) ;
  assign n5785 = ( ~n5672 & n5769 ) | ( ~n5672 & n5784 ) | ( n5769 & n5784 ) ;
  assign n5786 = ( n5672 & n5769 ) | ( n5672 & n5784 ) | ( n5769 & n5784 ) ;
  assign n5787 = ( n5672 & n5785 ) | ( n5672 & ~n5786 ) | ( n5785 & ~n5786 ) ;
  assign n5788 = ( n5722 & n5755 ) | ( n5722 & n5787 ) | ( n5755 & n5787 ) ;
  assign n5789 = ( n5722 & n5755 ) | ( n5722 & ~n5787 ) | ( n5755 & ~n5787 ) ;
  assign n5790 = ( n5787 & ~n5788 ) | ( n5787 & n5789 ) | ( ~n5788 & n5789 ) ;
  assign n5791 = ( n5705 & n5720 ) | ( n5705 & ~n5753 ) | ( n5720 & ~n5753 ) ;
  assign n5792 = ( n5705 & n5720 ) | ( n5705 & n5753 ) | ( n5720 & n5753 ) ;
  assign n5793 = ( n5753 & n5791 ) | ( n5753 & ~n5792 ) | ( n5791 & ~n5792 ) ;
  assign n5794 = ( n5696 & n5717 ) | ( n5696 & ~n5738 ) | ( n5717 & ~n5738 ) ;
  assign n5795 = ( n5696 & n5717 ) | ( n5696 & n5738 ) | ( n5717 & n5738 ) ;
  assign n5796 = ( n5738 & n5794 ) | ( n5738 & ~n5795 ) | ( n5794 & ~n5795 ) ;
  assign n5797 = ( n5689 & n5702 ) | ( n5689 & n5750 ) | ( n5702 & n5750 ) ;
  assign n5798 = ( n5689 & n5702 ) | ( n5689 & ~n5750 ) | ( n5702 & ~n5750 ) ;
  assign n5799 = ( n5750 & ~n5797 ) | ( n5750 & n5798 ) | ( ~n5797 & n5798 ) ;
  assign n5800 = ( n5679 & n5796 ) | ( n5679 & n5799 ) | ( n5796 & n5799 ) ;
  assign n5801 = ( n5679 & ~n5796 ) | ( n5679 & n5799 ) | ( ~n5796 & n5799 ) ;
  assign n5802 = ( n5796 & ~n5800 ) | ( n5796 & n5801 ) | ( ~n5800 & n5801 ) ;
  assign n5803 = ( n5681 & n5793 ) | ( n5681 & n5802 ) | ( n5793 & n5802 ) ;
  assign n5804 = ( n5681 & ~n5793 ) | ( n5681 & n5802 ) | ( ~n5793 & n5802 ) ;
  assign n5805 = ( n5793 & ~n5803 ) | ( n5793 & n5804 ) | ( ~n5803 & n5804 ) ;
  assign n5806 = ( ~n5758 & n5790 ) | ( ~n5758 & n5805 ) | ( n5790 & n5805 ) ;
  assign n5807 = ( n5758 & n5790 ) | ( n5758 & n5805 ) | ( n5790 & n5805 ) ;
  assign n5808 = ( n5758 & n5806 ) | ( n5758 & ~n5807 ) | ( n5806 & ~n5807 ) ;
  assign n5809 = x31 & x47 ;
  assign n5810 = x20 & x58 ;
  assign n5811 = x30 & x48 ;
  assign n5812 = ( ~n5809 & n5810 ) | ( ~n5809 & n5811 ) | ( n5810 & n5811 ) ;
  assign n5813 = ( n5809 & n5810 ) | ( n5809 & n5811 ) | ( n5810 & n5811 ) ;
  assign n5814 = ( n5809 & n5812 ) | ( n5809 & ~n5813 ) | ( n5812 & ~n5813 ) ;
  assign n5815 = x25 & x53 ;
  assign n5816 = x24 & x54 ;
  assign n5817 = x22 & x56 ;
  assign n5818 = ( ~n5815 & n5816 ) | ( ~n5815 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5819 = ( n5815 & n5816 ) | ( n5815 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5820 = ( n5815 & n5818 ) | ( n5815 & ~n5819 ) | ( n5818 & ~n5819 ) ;
  assign n5821 = x32 & x46 ;
  assign n5822 = x33 & x45 ;
  assign n5823 = x34 & x44 ;
  assign n5824 = ( ~n5821 & n5822 ) | ( ~n5821 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5825 = ( n5821 & n5822 ) | ( n5821 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5826 = ( n5821 & n5824 ) | ( n5821 & ~n5825 ) | ( n5824 & ~n5825 ) ;
  assign n5827 = ( ~n5814 & n5820 ) | ( ~n5814 & n5826 ) | ( n5820 & n5826 ) ;
  assign n5828 = ( n5814 & n5820 ) | ( n5814 & n5826 ) | ( n5820 & n5826 ) ;
  assign n5829 = ( n5814 & n5827 ) | ( n5814 & ~n5828 ) | ( n5827 & ~n5828 ) ;
  assign n5830 = x28 & x50 ;
  assign n5831 = x29 & x49 ;
  assign n5832 = ( ~n2844 & n5830 ) | ( ~n2844 & n5831 ) | ( n5830 & n5831 ) ;
  assign n5833 = ( n2844 & n5830 ) | ( n2844 & n5831 ) | ( n5830 & n5831 ) ;
  assign n5834 = ( n2844 & n5832 ) | ( n2844 & ~n5833 ) | ( n5832 & ~n5833 ) ;
  assign n5835 = x16 & x62 ;
  assign n5836 = x17 & x61 ;
  assign n5837 = x15 & x63 ;
  assign n5838 = ( ~n5835 & n5836 ) | ( ~n5835 & n5837 ) | ( n5836 & n5837 ) ;
  assign n5839 = ( n5835 & n5836 ) | ( n5835 & n5837 ) | ( n5836 & n5837 ) ;
  assign n5840 = ( n5835 & n5838 ) | ( n5835 & ~n5839 ) | ( n5838 & ~n5839 ) ;
  assign n5841 = x18 & x60 ;
  assign n5842 = x19 & x59 ;
  assign n5843 = x21 & x57 ;
  assign n5844 = ( ~n5841 & n5842 ) | ( ~n5841 & n5843 ) | ( n5842 & n5843 ) ;
  assign n5845 = ( n5841 & n5842 ) | ( n5841 & n5843 ) | ( n5842 & n5843 ) ;
  assign n5846 = ( n5841 & n5844 ) | ( n5841 & ~n5845 ) | ( n5844 & ~n5845 ) ;
  assign n5847 = ( ~n5834 & n5840 ) | ( ~n5834 & n5846 ) | ( n5840 & n5846 ) ;
  assign n5848 = ( n5834 & n5840 ) | ( n5834 & n5846 ) | ( n5840 & n5846 ) ;
  assign n5849 = ( n5834 & n5847 ) | ( n5834 & ~n5848 ) | ( n5847 & ~n5848 ) ;
  assign n5850 = ( n5726 & n5829 ) | ( n5726 & n5849 ) | ( n5829 & n5849 ) ;
  assign n5851 = ( ~n5726 & n5829 ) | ( ~n5726 & n5849 ) | ( n5829 & n5849 ) ;
  assign n5852 = ( n5726 & ~n5850 ) | ( n5726 & n5851 ) | ( ~n5850 & n5851 ) ;
  assign n5853 = ( n5685 & ~n5728 ) | ( n5685 & n5852 ) | ( ~n5728 & n5852 ) ;
  assign n5854 = ( n5685 & n5728 ) | ( n5685 & n5852 ) | ( n5728 & n5852 ) ;
  assign n5855 = ( n5728 & n5853 ) | ( n5728 & ~n5854 ) | ( n5853 & ~n5854 ) ;
  assign n5856 = ( n5731 & n5808 ) | ( n5731 & n5855 ) | ( n5808 & n5855 ) ;
  assign n5857 = ( n5731 & ~n5808 ) | ( n5731 & n5855 ) | ( ~n5808 & n5855 ) ;
  assign n5858 = ( n5808 & ~n5856 ) | ( n5808 & n5857 ) | ( ~n5856 & n5857 ) ;
  assign n5859 = ( n5761 & ~n5764 ) | ( n5761 & n5858 ) | ( ~n5764 & n5858 ) ;
  assign n5860 = ( n5761 & n5764 ) | ( n5761 & n5858 ) | ( n5764 & n5858 ) ;
  assign n5861 = ( n5764 & n5859 ) | ( n5764 & ~n5860 ) | ( n5859 & ~n5860 ) ;
  assign n5862 = ( n5795 & n5797 ) | ( n5795 & ~n5848 ) | ( n5797 & ~n5848 ) ;
  assign n5863 = ( n5795 & n5797 ) | ( n5795 & n5848 ) | ( n5797 & n5848 ) ;
  assign n5864 = ( n5848 & n5862 ) | ( n5848 & ~n5863 ) | ( n5862 & ~n5863 ) ;
  assign n5865 = ( ~n5786 & n5792 ) | ( ~n5786 & n5864 ) | ( n5792 & n5864 ) ;
  assign n5866 = ( n5786 & n5792 ) | ( n5786 & n5864 ) | ( n5792 & n5864 ) ;
  assign n5867 = ( n5786 & n5865 ) | ( n5786 & ~n5866 ) | ( n5865 & ~n5866 ) ;
  assign n5868 = x28 & x51 ;
  assign n5869 = x17 & x62 ;
  assign n5870 = ( ~x40 & n5868 ) | ( ~x40 & n5869 ) | ( n5868 & n5869 ) ;
  assign n5871 = ( x40 & n5868 ) | ( x40 & n5869 ) | ( n5868 & n5869 ) ;
  assign n5872 = ( x40 & n5870 ) | ( x40 & ~n5871 ) | ( n5870 & ~n5871 ) ;
  assign n5873 = x38 & x41 ;
  assign n5874 = x39 & x40 ;
  assign n5875 = x37 & x42 ;
  assign n5876 = ( ~n5873 & n5874 ) | ( ~n5873 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5877 = ( n5873 & n5874 ) | ( n5873 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5878 = ( n5873 & n5876 ) | ( n5873 & ~n5877 ) | ( n5876 & ~n5877 ) ;
  assign n5879 = x26 & x53 ;
  assign n5880 = x24 & x55 ;
  assign n5881 = x25 & x54 ;
  assign n5882 = ( ~n5879 & n5880 ) | ( ~n5879 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5883 = ( n5879 & n5880 ) | ( n5879 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5884 = ( n5879 & n5882 ) | ( n5879 & ~n5883 ) | ( n5882 & ~n5883 ) ;
  assign n5885 = ( ~n5872 & n5878 ) | ( ~n5872 & n5884 ) | ( n5878 & n5884 ) ;
  assign n5886 = ( n5872 & n5878 ) | ( n5872 & n5884 ) | ( n5878 & n5884 ) ;
  assign n5887 = ( n5872 & n5885 ) | ( n5872 & ~n5886 ) | ( n5885 & ~n5886 ) ;
  assign n5888 = x20 & x59 ;
  assign n5889 = x21 & x58 ;
  assign n5890 = x19 & x60 ;
  assign n5891 = ( ~n5888 & n5889 ) | ( ~n5888 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5892 = ( n5888 & n5889 ) | ( n5888 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5893 = ( n5888 & n5891 ) | ( n5888 & ~n5892 ) | ( n5891 & ~n5892 ) ;
  assign n5894 = x33 & x46 ;
  assign n5895 = x31 & x48 ;
  assign n5896 = x32 & x47 ;
  assign n5897 = ( ~n5894 & n5895 ) | ( ~n5894 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5898 = ( n5894 & n5895 ) | ( n5894 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5899 = ( n5894 & n5897 ) | ( n5894 & ~n5898 ) | ( n5897 & ~n5898 ) ;
  assign n5900 = x30 & x49 ;
  assign n5901 = x22 & x57 ;
  assign n5902 = x29 & x50 ;
  assign n5903 = ( ~n5900 & n5901 ) | ( ~n5900 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5904 = ( n5900 & n5901 ) | ( n5900 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5905 = ( n5900 & n5903 ) | ( n5900 & ~n5904 ) | ( n5903 & ~n5904 ) ;
  assign n5906 = ( ~n5893 & n5899 ) | ( ~n5893 & n5905 ) | ( n5899 & n5905 ) ;
  assign n5907 = ( n5893 & n5899 ) | ( n5893 & n5905 ) | ( n5899 & n5905 ) ;
  assign n5908 = ( n5893 & n5906 ) | ( n5893 & ~n5907 ) | ( n5906 & ~n5907 ) ;
  assign n5909 = ( n5800 & n5887 ) | ( n5800 & n5908 ) | ( n5887 & n5908 ) ;
  assign n5910 = ( ~n5800 & n5887 ) | ( ~n5800 & n5908 ) | ( n5887 & n5908 ) ;
  assign n5911 = ( n5800 & ~n5909 ) | ( n5800 & n5910 ) | ( ~n5909 & n5910 ) ;
  assign n5912 = ( n5803 & ~n5867 ) | ( n5803 & n5911 ) | ( ~n5867 & n5911 ) ;
  assign n5913 = ( n5803 & n5867 ) | ( n5803 & n5911 ) | ( n5867 & n5911 ) ;
  assign n5914 = ( n5867 & n5912 ) | ( n5867 & ~n5913 ) | ( n5912 & ~n5913 ) ;
  assign n5915 = x35 & x44 ;
  assign n5916 = x16 & x63 ;
  assign n5917 = x34 & x45 ;
  assign n5918 = ( ~n5915 & n5916 ) | ( ~n5915 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5919 = ( n5915 & n5916 ) | ( n5915 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5920 = ( n5915 & n5918 ) | ( n5915 & ~n5919 ) | ( n5918 & ~n5919 ) ;
  assign n5921 = x23 & x56 ;
  assign n5922 = x36 & x43 ;
  assign n5923 = ( ~n2906 & n5921 ) | ( ~n2906 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5924 = ( n2906 & n5921 ) | ( n2906 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5925 = ( n2906 & n5923 ) | ( n2906 & ~n5924 ) | ( n5923 & ~n5924 ) ;
  assign n5926 = ( ~n5768 & n5920 ) | ( ~n5768 & n5925 ) | ( n5920 & n5925 ) ;
  assign n5927 = ( n5768 & n5920 ) | ( n5768 & n5925 ) | ( n5920 & n5925 ) ;
  assign n5928 = ( n5768 & n5926 ) | ( n5768 & ~n5927 ) | ( n5926 & ~n5927 ) ;
  assign n5929 = ( ~n5819 & n5833 ) | ( ~n5819 & n5845 ) | ( n5833 & n5845 ) ;
  assign n5930 = ( n5819 & n5833 ) | ( n5819 & n5845 ) | ( n5833 & n5845 ) ;
  assign n5931 = ( n5819 & n5929 ) | ( n5819 & ~n5930 ) | ( n5929 & ~n5930 ) ;
  assign n5932 = ( n5783 & n5928 ) | ( n5783 & n5931 ) | ( n5928 & n5931 ) ;
  assign n5933 = ( n5783 & ~n5928 ) | ( n5783 & n5931 ) | ( ~n5928 & n5931 ) ;
  assign n5934 = ( n5928 & ~n5932 ) | ( n5928 & n5933 ) | ( ~n5932 & n5933 ) ;
  assign n5935 = ( n5813 & ~n5825 ) | ( n5813 & n5839 ) | ( ~n5825 & n5839 ) ;
  assign n5936 = ( n5813 & n5825 ) | ( n5813 & n5839 ) | ( n5825 & n5839 ) ;
  assign n5937 = ( n5825 & n5935 ) | ( n5825 & ~n5936 ) | ( n5935 & ~n5936 ) ;
  assign n5938 = x18 & x61 ;
  assign n5939 = ( n5774 & n5780 ) | ( n5774 & n5938 ) | ( n5780 & n5938 ) ;
  assign n5940 = ( ~n5774 & n5780 ) | ( ~n5774 & n5938 ) | ( n5780 & n5938 ) ;
  assign n5941 = ( n5774 & ~n5939 ) | ( n5774 & n5940 ) | ( ~n5939 & n5940 ) ;
  assign n5942 = ( n5828 & n5937 ) | ( n5828 & n5941 ) | ( n5937 & n5941 ) ;
  assign n5943 = ( ~n5828 & n5937 ) | ( ~n5828 & n5941 ) | ( n5937 & n5941 ) ;
  assign n5944 = ( n5828 & ~n5942 ) | ( n5828 & n5943 ) | ( ~n5942 & n5943 ) ;
  assign n5945 = ( n5850 & ~n5934 ) | ( n5850 & n5944 ) | ( ~n5934 & n5944 ) ;
  assign n5946 = ( n5850 & n5934 ) | ( n5850 & n5944 ) | ( n5934 & n5944 ) ;
  assign n5947 = ( n5934 & n5945 ) | ( n5934 & ~n5946 ) | ( n5945 & ~n5946 ) ;
  assign n5948 = ( n5788 & n5854 ) | ( n5788 & n5947 ) | ( n5854 & n5947 ) ;
  assign n5949 = ( n5788 & ~n5854 ) | ( n5788 & n5947 ) | ( ~n5854 & n5947 ) ;
  assign n5950 = ( n5854 & ~n5948 ) | ( n5854 & n5949 ) | ( ~n5948 & n5949 ) ;
  assign n5951 = ( ~n5807 & n5914 ) | ( ~n5807 & n5950 ) | ( n5914 & n5950 ) ;
  assign n5952 = ( n5807 & n5914 ) | ( n5807 & n5950 ) | ( n5914 & n5950 ) ;
  assign n5953 = ( n5807 & n5951 ) | ( n5807 & ~n5952 ) | ( n5951 & ~n5952 ) ;
  assign n5954 = ( n5856 & n5860 ) | ( n5856 & n5953 ) | ( n5860 & n5953 ) ;
  assign n5955 = ( n5856 & ~n5860 ) | ( n5856 & n5953 ) | ( ~n5860 & n5953 ) ;
  assign n5956 = ( n5860 & ~n5954 ) | ( n5860 & n5955 ) | ( ~n5954 & n5955 ) ;
  assign n5957 = ( n5930 & n5936 ) | ( n5930 & ~n5939 ) | ( n5936 & ~n5939 ) ;
  assign n5958 = ( n5930 & n5936 ) | ( n5930 & n5939 ) | ( n5936 & n5939 ) ;
  assign n5959 = ( n5939 & n5957 ) | ( n5939 & ~n5958 ) | ( n5957 & ~n5958 ) ;
  assign n5960 = ( n5932 & n5942 ) | ( n5932 & n5959 ) | ( n5942 & n5959 ) ;
  assign n5961 = ( n5932 & n5942 ) | ( n5932 & ~n5959 ) | ( n5942 & ~n5959 ) ;
  assign n5962 = ( n5959 & ~n5960 ) | ( n5959 & n5961 ) | ( ~n5960 & n5961 ) ;
  assign n5963 = ( ~n5883 & n5919 ) | ( ~n5883 & n5924 ) | ( n5919 & n5924 ) ;
  assign n5964 = ( n5883 & n5919 ) | ( n5883 & n5924 ) | ( n5919 & n5924 ) ;
  assign n5965 = ( n5883 & n5963 ) | ( n5883 & ~n5964 ) | ( n5963 & ~n5964 ) ;
  assign n5966 = ( n5863 & n5927 ) | ( n5863 & n5965 ) | ( n5927 & n5965 ) ;
  assign n5967 = ( n5863 & ~n5927 ) | ( n5863 & n5965 ) | ( ~n5927 & n5965 ) ;
  assign n5968 = ( n5927 & ~n5966 ) | ( n5927 & n5967 ) | ( ~n5966 & n5967 ) ;
  assign n5969 = ( n5892 & ~n5898 ) | ( n5892 & n5904 ) | ( ~n5898 & n5904 ) ;
  assign n5970 = ( n5892 & n5898 ) | ( n5892 & n5904 ) | ( n5898 & n5904 ) ;
  assign n5971 = ( n5898 & n5969 ) | ( n5898 & ~n5970 ) | ( n5969 & ~n5970 ) ;
  assign n5972 = ( n5886 & n5907 ) | ( n5886 & n5971 ) | ( n5907 & n5971 ) ;
  assign n5973 = ( n5886 & n5907 ) | ( n5886 & ~n5971 ) | ( n5907 & ~n5971 ) ;
  assign n5974 = ( n5971 & ~n5972 ) | ( n5971 & n5973 ) | ( ~n5972 & n5973 ) ;
  assign n5975 = ( n5909 & n5968 ) | ( n5909 & n5974 ) | ( n5968 & n5974 ) ;
  assign n5976 = ( n5909 & ~n5968 ) | ( n5909 & n5974 ) | ( ~n5968 & n5974 ) ;
  assign n5977 = ( n5968 & ~n5975 ) | ( n5968 & n5976 ) | ( ~n5975 & n5976 ) ;
  assign n5978 = ( n5913 & n5962 ) | ( n5913 & n5977 ) | ( n5962 & n5977 ) ;
  assign n5979 = ( n5913 & ~n5962 ) | ( n5913 & n5977 ) | ( ~n5962 & n5977 ) ;
  assign n5980 = ( n5962 & ~n5978 ) | ( n5962 & n5979 ) | ( ~n5978 & n5979 ) ;
  assign n5981 = x19 & x61 ;
  assign n5982 = x18 & x62 ;
  assign n5983 = ( n5871 & n5981 ) | ( n5871 & n5982 ) | ( n5981 & n5982 ) ;
  assign n5984 = ( ~n5871 & n5981 ) | ( ~n5871 & n5982 ) | ( n5981 & n5982 ) ;
  assign n5985 = ( n5871 & ~n5983 ) | ( n5871 & n5984 ) | ( ~n5983 & n5984 ) ;
  assign n5986 = x33 & x47 ;
  assign n5987 = x17 & x63 ;
  assign n5988 = x29 & x51 ;
  assign n5989 = ( ~n5986 & n5987 ) | ( ~n5986 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5990 = ( n5986 & n5987 ) | ( n5986 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5991 = ( n5986 & n5989 ) | ( n5986 & ~n5990 ) | ( n5989 & ~n5990 ) ;
  assign n5992 = x35 & x45 ;
  assign n5993 = x36 & x44 ;
  assign n5994 = x34 & x46 ;
  assign n5995 = ( ~n5992 & n5993 ) | ( ~n5992 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5996 = ( n5992 & n5993 ) | ( n5992 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5997 = ( n5992 & n5995 ) | ( n5992 & ~n5996 ) | ( n5995 & ~n5996 ) ;
  assign n5998 = ( n5985 & n5991 ) | ( n5985 & n5997 ) | ( n5991 & n5997 ) ;
  assign n5999 = ( ~n5985 & n5991 ) | ( ~n5985 & n5997 ) | ( n5991 & n5997 ) ;
  assign n6000 = ( n5985 & ~n5998 ) | ( n5985 & n5999 ) | ( ~n5998 & n5999 ) ;
  assign n6001 = x22 & x58 ;
  assign n6002 = x20 & x60 ;
  assign n6003 = x21 & x59 ;
  assign n6004 = ( ~n6001 & n6002 ) | ( ~n6001 & n6003 ) | ( n6002 & n6003 ) ;
  assign n6005 = ( n6001 & n6002 ) | ( n6001 & n6003 ) | ( n6002 & n6003 ) ;
  assign n6006 = ( n6001 & n6004 ) | ( n6001 & ~n6005 ) | ( n6004 & ~n6005 ) ;
  assign n6007 = x32 & x48 ;
  assign n6008 = x31 & x49 ;
  assign n6009 = x30 & x50 ;
  assign n6010 = ( ~n6007 & n6008 ) | ( ~n6007 & n6009 ) | ( n6008 & n6009 ) ;
  assign n6011 = ( n6007 & n6008 ) | ( n6007 & n6009 ) | ( n6008 & n6009 ) ;
  assign n6012 = ( n6007 & n6010 ) | ( n6007 & ~n6011 ) | ( n6010 & ~n6011 ) ;
  assign n6013 = ( n5877 & ~n6006 ) | ( n5877 & n6012 ) | ( ~n6006 & n6012 ) ;
  assign n6014 = ( n5877 & n6006 ) | ( n5877 & n6012 ) | ( n6006 & n6012 ) ;
  assign n6015 = ( n6006 & n6013 ) | ( n6006 & ~n6014 ) | ( n6013 & ~n6014 ) ;
  assign n6016 = x39 & x41 ;
  assign n6017 = x27 & x53 ;
  assign n6018 = x28 & x52 ;
  assign n6019 = ( ~n6016 & n6017 ) | ( ~n6016 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6020 = ( n6016 & n6017 ) | ( n6016 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6021 = ( n6016 & n6019 ) | ( n6016 & ~n6020 ) | ( n6019 & ~n6020 ) ;
  assign n6022 = x25 & x55 ;
  assign n6023 = x37 & x43 ;
  assign n6024 = x38 & x42 ;
  assign n6025 = ( ~n6022 & n6023 ) | ( ~n6022 & n6024 ) | ( n6023 & n6024 ) ;
  assign n6026 = ( n6022 & n6023 ) | ( n6022 & n6024 ) | ( n6023 & n6024 ) ;
  assign n6027 = ( n6022 & n6025 ) | ( n6022 & ~n6026 ) | ( n6025 & ~n6026 ) ;
  assign n6028 = x26 & x54 ;
  assign n6029 = x23 & x57 ;
  assign n6030 = x24 & x56 ;
  assign n6031 = ( ~n6028 & n6029 ) | ( ~n6028 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6032 = ( n6028 & n6029 ) | ( n6028 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6033 = ( n6028 & n6031 ) | ( n6028 & ~n6032 ) | ( n6031 & ~n6032 ) ;
  assign n6034 = ( ~n6021 & n6027 ) | ( ~n6021 & n6033 ) | ( n6027 & n6033 ) ;
  assign n6035 = ( n6021 & n6027 ) | ( n6021 & n6033 ) | ( n6027 & n6033 ) ;
  assign n6036 = ( n6021 & n6034 ) | ( n6021 & ~n6035 ) | ( n6034 & ~n6035 ) ;
  assign n6037 = ( n6000 & n6015 ) | ( n6000 & n6036 ) | ( n6015 & n6036 ) ;
  assign n6038 = ( ~n6000 & n6015 ) | ( ~n6000 & n6036 ) | ( n6015 & n6036 ) ;
  assign n6039 = ( n6000 & ~n6037 ) | ( n6000 & n6038 ) | ( ~n6037 & n6038 ) ;
  assign n6040 = ( n5866 & n5946 ) | ( n5866 & n6039 ) | ( n5946 & n6039 ) ;
  assign n6041 = ( n5866 & ~n5946 ) | ( n5866 & n6039 ) | ( ~n5946 & n6039 ) ;
  assign n6042 = ( n5946 & ~n6040 ) | ( n5946 & n6041 ) | ( ~n6040 & n6041 ) ;
  assign n6043 = ( n5948 & n5980 ) | ( n5948 & n6042 ) | ( n5980 & n6042 ) ;
  assign n6044 = ( ~n5948 & n5980 ) | ( ~n5948 & n6042 ) | ( n5980 & n6042 ) ;
  assign n6045 = ( n5948 & ~n6043 ) | ( n5948 & n6044 ) | ( ~n6043 & n6044 ) ;
  assign n6046 = ( n5952 & n5954 ) | ( n5952 & n6045 ) | ( n5954 & n6045 ) ;
  assign n6047 = ( n5952 & ~n5954 ) | ( n5952 & n6045 ) | ( ~n5954 & n6045 ) ;
  assign n6048 = ( n5954 & ~n6046 ) | ( n5954 & n6047 ) | ( ~n6046 & n6047 ) ;
  assign n6049 = x31 & x50 ;
  assign n6050 = x32 & x49 ;
  assign n6051 = x30 & x51 ;
  assign n6052 = ( ~n6049 & n6050 ) | ( ~n6049 & n6051 ) | ( n6050 & n6051 ) ;
  assign n6053 = ( n6049 & n6050 ) | ( n6049 & n6051 ) | ( n6050 & n6051 ) ;
  assign n6054 = ( n6049 & n6052 ) | ( n6049 & ~n6053 ) | ( n6052 & ~n6053 ) ;
  assign n6055 = ( ~n5983 & n5996 ) | ( ~n5983 & n6054 ) | ( n5996 & n6054 ) ;
  assign n6056 = ( n5983 & n5996 ) | ( n5983 & n6054 ) | ( n5996 & n6054 ) ;
  assign n6057 = ( n5983 & n6055 ) | ( n5983 & ~n6056 ) | ( n6055 & ~n6056 ) ;
  assign n6058 = ( n5990 & ~n6005 ) | ( n5990 & n6011 ) | ( ~n6005 & n6011 ) ;
  assign n6059 = ( n5990 & n6005 ) | ( n5990 & n6011 ) | ( n6005 & n6011 ) ;
  assign n6060 = ( n6005 & n6058 ) | ( n6005 & ~n6059 ) | ( n6058 & ~n6059 ) ;
  assign n6061 = ( n5998 & ~n6057 ) | ( n5998 & n6060 ) | ( ~n6057 & n6060 ) ;
  assign n6062 = ( n5998 & n6057 ) | ( n5998 & n6060 ) | ( n6057 & n6060 ) ;
  assign n6063 = ( n6057 & n6061 ) | ( n6057 & ~n6062 ) | ( n6061 & ~n6062 ) ;
  assign n6064 = ( n6020 & ~n6026 ) | ( n6020 & n6032 ) | ( ~n6026 & n6032 ) ;
  assign n6065 = ( n6020 & n6026 ) | ( n6020 & n6032 ) | ( n6026 & n6032 ) ;
  assign n6066 = ( n6026 & n6064 ) | ( n6026 & ~n6065 ) | ( n6064 & ~n6065 ) ;
  assign n6067 = ( n6014 & n6035 ) | ( n6014 & n6066 ) | ( n6035 & n6066 ) ;
  assign n6068 = ( ~n6014 & n6035 ) | ( ~n6014 & n6066 ) | ( n6035 & n6066 ) ;
  assign n6069 = ( n6014 & ~n6067 ) | ( n6014 & n6068 ) | ( ~n6067 & n6068 ) ;
  assign n6070 = ( n6037 & n6063 ) | ( n6037 & n6069 ) | ( n6063 & n6069 ) ;
  assign n6071 = ( ~n6037 & n6063 ) | ( ~n6037 & n6069 ) | ( n6063 & n6069 ) ;
  assign n6072 = ( n6037 & ~n6070 ) | ( n6037 & n6071 ) | ( ~n6070 & n6071 ) ;
  assign n6073 = x38 & x43 ;
  assign n6074 = x39 & x42 ;
  assign n6075 = x27 & x54 ;
  assign n6076 = ( ~n6073 & n6074 ) | ( ~n6073 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6077 = ( n6073 & n6074 ) | ( n6073 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6078 = ( n6073 & n6076 ) | ( n6073 & ~n6077 ) | ( n6076 & ~n6077 ) ;
  assign n6079 = ( ~n5964 & n5970 ) | ( ~n5964 & n6078 ) | ( n5970 & n6078 ) ;
  assign n6080 = ( n5964 & n5970 ) | ( n5964 & n6078 ) | ( n5970 & n6078 ) ;
  assign n6081 = ( n5964 & n6079 ) | ( n5964 & ~n6080 ) | ( n6079 & ~n6080 ) ;
  assign n6082 = ( ~n5966 & n5972 ) | ( ~n5966 & n6081 ) | ( n5972 & n6081 ) ;
  assign n6083 = ( n5966 & n5972 ) | ( n5966 & n6081 ) | ( n5972 & n6081 ) ;
  assign n6084 = ( n5966 & n6082 ) | ( n5966 & ~n6083 ) | ( n6082 & ~n6083 ) ;
  assign n6085 = ( n6040 & ~n6072 ) | ( n6040 & n6084 ) | ( ~n6072 & n6084 ) ;
  assign n6086 = ( n6040 & n6072 ) | ( n6040 & n6084 ) | ( n6072 & n6084 ) ;
  assign n6087 = ( n6072 & n6085 ) | ( n6072 & ~n6086 ) | ( n6085 & ~n6086 ) ;
  assign n6088 = x37 & x44 ;
  assign n6089 = x35 & x46 ;
  assign n6090 = x36 & x45 ;
  assign n6091 = ( ~n6088 & n6089 ) | ( ~n6088 & n6090 ) | ( n6089 & n6090 ) ;
  assign n6092 = ( n6088 & n6089 ) | ( n6088 & n6090 ) | ( n6089 & n6090 ) ;
  assign n6093 = ( n6088 & n6091 ) | ( n6088 & ~n6092 ) | ( n6091 & ~n6092 ) ;
  assign n6094 = x21 & x60 ;
  assign n6095 = x20 & x61 ;
  assign n6096 = x18 & x63 ;
  assign n6097 = ( ~n6094 & n6095 ) | ( ~n6094 & n6096 ) | ( n6095 & n6096 ) ;
  assign n6098 = ( n6094 & n6095 ) | ( n6094 & n6096 ) | ( n6095 & n6096 ) ;
  assign n6099 = ( n6094 & n6097 ) | ( n6094 & ~n6098 ) | ( n6097 & ~n6098 ) ;
  assign n6100 = x29 & x52 ;
  assign n6101 = x26 & x55 ;
  assign n6102 = ( ~n3009 & n6100 ) | ( ~n3009 & n6101 ) | ( n6100 & n6101 ) ;
  assign n6103 = ( n3009 & n6100 ) | ( n3009 & n6101 ) | ( n6100 & n6101 ) ;
  assign n6104 = ( n3009 & n6102 ) | ( n3009 & ~n6103 ) | ( n6102 & ~n6103 ) ;
  assign n6105 = ( ~n6093 & n6099 ) | ( ~n6093 & n6104 ) | ( n6099 & n6104 ) ;
  assign n6106 = ( n6093 & n6099 ) | ( n6093 & n6104 ) | ( n6099 & n6104 ) ;
  assign n6107 = ( n6093 & n6105 ) | ( n6093 & ~n6106 ) | ( n6105 & ~n6106 ) ;
  assign n6108 = x19 & x62 ;
  assign n6109 = x40 & x41 ;
  assign n6110 = ( x41 & n6108 ) | ( x41 & n6109 ) | ( n6108 & n6109 ) ;
  assign n6111 = ( x41 & ~n6108 ) | ( x41 & n6109 ) | ( ~n6108 & n6109 ) ;
  assign n6112 = ( n6108 & ~n6110 ) | ( n6108 & n6111 ) | ( ~n6110 & n6111 ) ;
  assign n6113 = x34 & x47 ;
  assign n6114 = x24 & x57 ;
  assign n6115 = x33 & x48 ;
  assign n6116 = ( ~n6113 & n6114 ) | ( ~n6113 & n6115 ) | ( n6114 & n6115 ) ;
  assign n6117 = ( n6113 & n6114 ) | ( n6113 & n6115 ) | ( n6114 & n6115 ) ;
  assign n6118 = ( n6113 & n6116 ) | ( n6113 & ~n6117 ) | ( n6116 & ~n6117 ) ;
  assign n6119 = x25 & x56 ;
  assign n6120 = x22 & x59 ;
  assign n6121 = x23 & x58 ;
  assign n6122 = ( ~n6119 & n6120 ) | ( ~n6119 & n6121 ) | ( n6120 & n6121 ) ;
  assign n6123 = ( n6119 & n6120 ) | ( n6119 & n6121 ) | ( n6120 & n6121 ) ;
  assign n6124 = ( n6119 & n6122 ) | ( n6119 & ~n6123 ) | ( n6122 & ~n6123 ) ;
  assign n6125 = ( ~n6112 & n6118 ) | ( ~n6112 & n6124 ) | ( n6118 & n6124 ) ;
  assign n6126 = ( n6112 & n6118 ) | ( n6112 & n6124 ) | ( n6118 & n6124 ) ;
  assign n6127 = ( n6112 & n6125 ) | ( n6112 & ~n6126 ) | ( n6125 & ~n6126 ) ;
  assign n6128 = ( n5958 & n6107 ) | ( n5958 & n6127 ) | ( n6107 & n6127 ) ;
  assign n6129 = ( ~n5958 & n6107 ) | ( ~n5958 & n6127 ) | ( n6107 & n6127 ) ;
  assign n6130 = ( n5958 & ~n6128 ) | ( n5958 & n6129 ) | ( ~n6128 & n6129 ) ;
  assign n6131 = ( n5960 & n5975 ) | ( n5960 & n6130 ) | ( n5975 & n6130 ) ;
  assign n6132 = ( ~n5960 & n5975 ) | ( ~n5960 & n6130 ) | ( n5975 & n6130 ) ;
  assign n6133 = ( n5960 & ~n6131 ) | ( n5960 & n6132 ) | ( ~n6131 & n6132 ) ;
  assign n6134 = ( ~n5978 & n6087 ) | ( ~n5978 & n6133 ) | ( n6087 & n6133 ) ;
  assign n6135 = ( n5978 & n6087 ) | ( n5978 & n6133 ) | ( n6087 & n6133 ) ;
  assign n6136 = ( n5978 & n6134 ) | ( n5978 & ~n6135 ) | ( n6134 & ~n6135 ) ;
  assign n6137 = ( n6043 & ~n6046 ) | ( n6043 & n6136 ) | ( ~n6046 & n6136 ) ;
  assign n6138 = ( n6043 & n6046 ) | ( n6043 & n6136 ) | ( n6046 & n6136 ) ;
  assign n6139 = ( n6046 & n6137 ) | ( n6046 & ~n6138 ) | ( n6137 & ~n6138 ) ;
  assign n6140 = x25 & x57 ;
  assign n6141 = x28 & x54 ;
  assign n6142 = x27 & x55 ;
  assign n6143 = ( ~n6140 & n6141 ) | ( ~n6140 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6144 = ( n6140 & n6141 ) | ( n6140 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6145 = ( n6140 & n6143 ) | ( n6140 & ~n6144 ) | ( n6143 & ~n6144 ) ;
  assign n6146 = ( ~n6059 & n6065 ) | ( ~n6059 & n6145 ) | ( n6065 & n6145 ) ;
  assign n6147 = ( n6059 & n6065 ) | ( n6059 & n6145 ) | ( n6065 & n6145 ) ;
  assign n6148 = ( n6059 & n6146 ) | ( n6059 & ~n6147 ) | ( n6146 & ~n6147 ) ;
  assign n6149 = ( ~n6062 & n6067 ) | ( ~n6062 & n6148 ) | ( n6067 & n6148 ) ;
  assign n6150 = ( n6062 & n6067 ) | ( n6062 & n6148 ) | ( n6067 & n6148 ) ;
  assign n6151 = ( n6062 & n6149 ) | ( n6062 & ~n6150 ) | ( n6149 & ~n6150 ) ;
  assign n6152 = x19 & x63 ;
  assign n6153 = ( n6077 & n6110 ) | ( n6077 & n6152 ) | ( n6110 & n6152 ) ;
  assign n6154 = ( ~n6077 & n6110 ) | ( ~n6077 & n6152 ) | ( n6110 & n6152 ) ;
  assign n6155 = ( n6077 & ~n6153 ) | ( n6077 & n6154 ) | ( ~n6153 & n6154 ) ;
  assign n6156 = ( n6056 & n6126 ) | ( n6056 & n6155 ) | ( n6126 & n6155 ) ;
  assign n6157 = ( ~n6056 & n6126 ) | ( ~n6056 & n6155 ) | ( n6126 & n6155 ) ;
  assign n6158 = ( n6056 & ~n6156 ) | ( n6056 & n6157 ) | ( ~n6156 & n6157 ) ;
  assign n6159 = ( n6053 & ~n6103 ) | ( n6053 & n6117 ) | ( ~n6103 & n6117 ) ;
  assign n6160 = ( n6053 & n6103 ) | ( n6053 & n6117 ) | ( n6103 & n6117 ) ;
  assign n6161 = ( n6103 & n6159 ) | ( n6103 & ~n6160 ) | ( n6159 & ~n6160 ) ;
  assign n6162 = ( n6092 & ~n6098 ) | ( n6092 & n6123 ) | ( ~n6098 & n6123 ) ;
  assign n6163 = ( n6092 & n6098 ) | ( n6092 & n6123 ) | ( n6098 & n6123 ) ;
  assign n6164 = ( n6098 & n6162 ) | ( n6098 & ~n6163 ) | ( n6162 & ~n6163 ) ;
  assign n6165 = ( n6106 & n6161 ) | ( n6106 & n6164 ) | ( n6161 & n6164 ) ;
  assign n6166 = ( ~n6106 & n6161 ) | ( ~n6106 & n6164 ) | ( n6161 & n6164 ) ;
  assign n6167 = ( n6106 & ~n6165 ) | ( n6106 & n6166 ) | ( ~n6165 & n6166 ) ;
  assign n6168 = ( n6128 & ~n6158 ) | ( n6128 & n6167 ) | ( ~n6158 & n6167 ) ;
  assign n6169 = ( n6128 & n6158 ) | ( n6128 & n6167 ) | ( n6158 & n6167 ) ;
  assign n6170 = ( n6158 & n6168 ) | ( n6158 & ~n6169 ) | ( n6168 & ~n6169 ) ;
  assign n6171 = ( n6131 & n6151 ) | ( n6131 & n6170 ) | ( n6151 & n6170 ) ;
  assign n6172 = ( ~n6131 & n6151 ) | ( ~n6131 & n6170 ) | ( n6151 & n6170 ) ;
  assign n6173 = ( n6131 & ~n6171 ) | ( n6131 & n6172 ) | ( ~n6171 & n6172 ) ;
  assign n6174 = x39 & x43 ;
  assign n6175 = x38 & x44 ;
  assign n6176 = x26 & x56 ;
  assign n6177 = ( ~n6174 & n6175 ) | ( ~n6174 & n6176 ) | ( n6175 & n6176 ) ;
  assign n6178 = ( n6174 & n6175 ) | ( n6174 & n6176 ) | ( n6175 & n6176 ) ;
  assign n6179 = ( n6174 & n6177 ) | ( n6174 & ~n6178 ) | ( n6177 & ~n6178 ) ;
  assign n6180 = x36 & x46 ;
  assign n6181 = x37 & x45 ;
  assign n6182 = x35 & x47 ;
  assign n6183 = ( ~n6180 & n6181 ) | ( ~n6180 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6184 = ( n6180 & n6181 ) | ( n6180 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6185 = ( n6180 & n6183 ) | ( n6180 & ~n6184 ) | ( n6183 & ~n6184 ) ;
  assign n6186 = x40 & x42 ;
  assign n6187 = x30 & x52 ;
  assign n6188 = x29 & x53 ;
  assign n6189 = ( ~n6186 & n6187 ) | ( ~n6186 & n6188 ) | ( n6187 & n6188 ) ;
  assign n6190 = ( n6186 & n6187 ) | ( n6186 & n6188 ) | ( n6187 & n6188 ) ;
  assign n6191 = ( n6186 & n6189 ) | ( n6186 & ~n6190 ) | ( n6189 & ~n6190 ) ;
  assign n6192 = ( ~n6179 & n6185 ) | ( ~n6179 & n6191 ) | ( n6185 & n6191 ) ;
  assign n6193 = ( n6179 & n6185 ) | ( n6179 & n6191 ) | ( n6185 & n6191 ) ;
  assign n6194 = ( n6179 & n6192 ) | ( n6179 & ~n6193 ) | ( n6192 & ~n6193 ) ;
  assign n6195 = x23 & x59 ;
  assign n6196 = x24 & x58 ;
  assign n6197 = x22 & x60 ;
  assign n6198 = ( ~n6195 & n6196 ) | ( ~n6195 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = ( n6195 & n6196 ) | ( n6195 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6200 = ( n6195 & n6198 ) | ( n6195 & ~n6199 ) | ( n6198 & ~n6199 ) ;
  assign n6201 = x33 & x49 ;
  assign n6202 = x34 & x48 ;
  assign n6203 = x32 & x50 ;
  assign n6204 = ( ~n6201 & n6202 ) | ( ~n6201 & n6203 ) | ( n6202 & n6203 ) ;
  assign n6205 = ( n6201 & n6202 ) | ( n6201 & n6203 ) | ( n6202 & n6203 ) ;
  assign n6206 = ( n6201 & n6204 ) | ( n6201 & ~n6205 ) | ( n6204 & ~n6205 ) ;
  assign n6207 = x20 & x62 ;
  assign n6208 = x31 & x51 ;
  assign n6209 = x21 & x61 ;
  assign n6210 = ( ~n6207 & n6208 ) | ( ~n6207 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6211 = ( n6207 & n6208 ) | ( n6207 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6212 = ( n6207 & n6210 ) | ( n6207 & ~n6211 ) | ( n6210 & ~n6211 ) ;
  assign n6213 = ( ~n6200 & n6206 ) | ( ~n6200 & n6212 ) | ( n6206 & n6212 ) ;
  assign n6214 = ( n6200 & n6206 ) | ( n6200 & n6212 ) | ( n6206 & n6212 ) ;
  assign n6215 = ( n6200 & n6213 ) | ( n6200 & ~n6214 ) | ( n6213 & ~n6214 ) ;
  assign n6216 = ( n6080 & n6194 ) | ( n6080 & n6215 ) | ( n6194 & n6215 ) ;
  assign n6217 = ( ~n6080 & n6194 ) | ( ~n6080 & n6215 ) | ( n6194 & n6215 ) ;
  assign n6218 = ( n6080 & ~n6216 ) | ( n6080 & n6217 ) | ( ~n6216 & n6217 ) ;
  assign n6219 = ( n6070 & n6083 ) | ( n6070 & n6218 ) | ( n6083 & n6218 ) ;
  assign n6220 = ( n6070 & ~n6083 ) | ( n6070 & n6218 ) | ( ~n6083 & n6218 ) ;
  assign n6221 = ( n6083 & ~n6219 ) | ( n6083 & n6220 ) | ( ~n6219 & n6220 ) ;
  assign n6222 = ( n6086 & n6173 ) | ( n6086 & n6221 ) | ( n6173 & n6221 ) ;
  assign n6223 = ( ~n6086 & n6173 ) | ( ~n6086 & n6221 ) | ( n6173 & n6221 ) ;
  assign n6224 = ( n6086 & ~n6222 ) | ( n6086 & n6223 ) | ( ~n6222 & n6223 ) ;
  assign n6225 = ( n6135 & n6138 ) | ( n6135 & n6224 ) | ( n6138 & n6224 ) ;
  assign n6226 = ( n6135 & ~n6138 ) | ( n6135 & n6224 ) | ( ~n6138 & n6224 ) ;
  assign n6227 = ( n6138 & ~n6225 ) | ( n6138 & n6226 ) | ( ~n6225 & n6226 ) ;
  assign n6228 = ( n6160 & n6163 ) | ( n6160 & ~n6214 ) | ( n6163 & ~n6214 ) ;
  assign n6229 = ( n6160 & n6163 ) | ( n6160 & n6214 ) | ( n6163 & n6214 ) ;
  assign n6230 = ( n6214 & n6228 ) | ( n6214 & ~n6229 ) | ( n6228 & ~n6229 ) ;
  assign n6231 = x24 & x59 ;
  assign n6232 = x23 & x60 ;
  assign n6233 = ( n6190 & n6231 ) | ( n6190 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6234 = ( ~n6190 & n6231 ) | ( ~n6190 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6235 = ( n6190 & ~n6233 ) | ( n6190 & n6234 ) | ( ~n6233 & n6234 ) ;
  assign n6236 = x28 & x55 ;
  assign n6237 = x30 & x53 ;
  assign n6238 = x31 & x52 ;
  assign n6239 = ( ~n6236 & n6237 ) | ( ~n6236 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6240 = ( n6236 & n6237 ) | ( n6236 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6241 = ( n6236 & n6239 ) | ( n6236 & ~n6240 ) | ( n6239 & ~n6240 ) ;
  assign n6242 = ( n6153 & n6235 ) | ( n6153 & n6241 ) | ( n6235 & n6241 ) ;
  assign n6243 = ( n6153 & ~n6235 ) | ( n6153 & n6241 ) | ( ~n6235 & n6241 ) ;
  assign n6244 = ( n6235 & ~n6242 ) | ( n6235 & n6243 ) | ( ~n6242 & n6243 ) ;
  assign n6245 = ( n6156 & n6230 ) | ( n6156 & n6244 ) | ( n6230 & n6244 ) ;
  assign n6246 = ( ~n6156 & n6230 ) | ( ~n6156 & n6244 ) | ( n6230 & n6244 ) ;
  assign n6247 = ( n6156 & ~n6245 ) | ( n6156 & n6246 ) | ( ~n6245 & n6246 ) ;
  assign n6248 = ( n6178 & ~n6184 ) | ( n6178 & n6199 ) | ( ~n6184 & n6199 ) ;
  assign n6249 = ( n6178 & n6184 ) | ( n6178 & n6199 ) | ( n6184 & n6199 ) ;
  assign n6250 = ( n6184 & n6248 ) | ( n6184 & ~n6249 ) | ( n6248 & ~n6249 ) ;
  assign n6251 = ( n6144 & n6205 ) | ( n6144 & ~n6211 ) | ( n6205 & ~n6211 ) ;
  assign n6252 = ( n6144 & n6205 ) | ( n6144 & n6211 ) | ( n6205 & n6211 ) ;
  assign n6253 = ( n6211 & n6251 ) | ( n6211 & ~n6252 ) | ( n6251 & ~n6252 ) ;
  assign n6254 = ( n6193 & n6250 ) | ( n6193 & n6253 ) | ( n6250 & n6253 ) ;
  assign n6255 = ( ~n6193 & n6250 ) | ( ~n6193 & n6253 ) | ( n6250 & n6253 ) ;
  assign n6256 = ( n6193 & ~n6254 ) | ( n6193 & n6255 ) | ( ~n6254 & n6255 ) ;
  assign n6257 = ( n6165 & n6216 ) | ( n6165 & ~n6256 ) | ( n6216 & ~n6256 ) ;
  assign n6258 = ( n6165 & n6216 ) | ( n6165 & n6256 ) | ( n6216 & n6256 ) ;
  assign n6259 = ( n6256 & n6257 ) | ( n6256 & ~n6258 ) | ( n6257 & ~n6258 ) ;
  assign n6260 = ( n6219 & n6247 ) | ( n6219 & n6259 ) | ( n6247 & n6259 ) ;
  assign n6261 = ( ~n6219 & n6247 ) | ( ~n6219 & n6259 ) | ( n6247 & n6259 ) ;
  assign n6262 = ( n6219 & ~n6260 ) | ( n6219 & n6261 ) | ( ~n6260 & n6261 ) ;
  assign n6263 = x20 & x63 ;
  assign n6264 = x27 & x56 ;
  assign n6265 = x22 & x61 ;
  assign n6266 = ( ~n6263 & n6264 ) | ( ~n6263 & n6265 ) | ( n6264 & n6265 ) ;
  assign n6267 = ( n6263 & n6264 ) | ( n6263 & n6265 ) | ( n6264 & n6265 ) ;
  assign n6268 = ( n6263 & n6266 ) | ( n6263 & ~n6267 ) | ( n6266 & ~n6267 ) ;
  assign n6269 = x36 & x47 ;
  assign n6270 = x37 & x46 ;
  assign n6271 = x38 & x45 ;
  assign n6272 = ( ~n6269 & n6270 ) | ( ~n6269 & n6271 ) | ( n6270 & n6271 ) ;
  assign n6273 = ( n6269 & n6270 ) | ( n6269 & n6271 ) | ( n6270 & n6271 ) ;
  assign n6274 = ( n6269 & n6272 ) | ( n6269 & ~n6273 ) | ( n6272 & ~n6273 ) ;
  assign n6275 = x32 & x51 ;
  assign n6276 = x26 & x57 ;
  assign n6277 = x25 & x58 ;
  assign n6278 = ( ~n6275 & n6276 ) | ( ~n6275 & n6277 ) | ( n6276 & n6277 ) ;
  assign n6279 = ( n6275 & n6276 ) | ( n6275 & n6277 ) | ( n6276 & n6277 ) ;
  assign n6280 = ( n6275 & n6278 ) | ( n6275 & ~n6279 ) | ( n6278 & ~n6279 ) ;
  assign n6281 = ( ~n6268 & n6274 ) | ( ~n6268 & n6280 ) | ( n6274 & n6280 ) ;
  assign n6282 = ( n6268 & n6274 ) | ( n6268 & n6280 ) | ( n6274 & n6280 ) ;
  assign n6283 = ( n6268 & n6281 ) | ( n6268 & ~n6282 ) | ( n6281 & ~n6282 ) ;
  assign n6284 = x40 & x43 ;
  assign n6285 = x29 & x54 ;
  assign n6286 = x39 & x44 ;
  assign n6287 = ( ~n6284 & n6285 ) | ( ~n6284 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = ( n6284 & n6285 ) | ( n6284 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6289 = ( n6284 & n6287 ) | ( n6284 & ~n6288 ) | ( n6287 & ~n6288 ) ;
  assign n6290 = x34 & x49 ;
  assign n6291 = x33 & x50 ;
  assign n6292 = x35 & x48 ;
  assign n6293 = ( ~n6290 & n6291 ) | ( ~n6290 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6294 = ( n6290 & n6291 ) | ( n6290 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6295 = ( n6290 & n6293 ) | ( n6290 & ~n6294 ) | ( n6293 & ~n6294 ) ;
  assign n6296 = x21 & x62 ;
  assign n6297 = x41 & x42 ;
  assign n6298 = ( x42 & n6296 ) | ( x42 & n6297 ) | ( n6296 & n6297 ) ;
  assign n6299 = ( x42 & ~n6296 ) | ( x42 & n6297 ) | ( ~n6296 & n6297 ) ;
  assign n6300 = ( n6296 & ~n6298 ) | ( n6296 & n6299 ) | ( ~n6298 & n6299 ) ;
  assign n6301 = ( ~n6289 & n6295 ) | ( ~n6289 & n6300 ) | ( n6295 & n6300 ) ;
  assign n6302 = ( n6289 & n6295 ) | ( n6289 & n6300 ) | ( n6295 & n6300 ) ;
  assign n6303 = ( n6289 & n6301 ) | ( n6289 & ~n6302 ) | ( n6301 & ~n6302 ) ;
  assign n6304 = ( n6147 & n6283 ) | ( n6147 & n6303 ) | ( n6283 & n6303 ) ;
  assign n6305 = ( ~n6147 & n6283 ) | ( ~n6147 & n6303 ) | ( n6283 & n6303 ) ;
  assign n6306 = ( n6147 & ~n6304 ) | ( n6147 & n6305 ) | ( ~n6304 & n6305 ) ;
  assign n6307 = ( n6150 & n6169 ) | ( n6150 & n6306 ) | ( n6169 & n6306 ) ;
  assign n6308 = ( ~n6150 & n6169 ) | ( ~n6150 & n6306 ) | ( n6169 & n6306 ) ;
  assign n6309 = ( n6150 & ~n6307 ) | ( n6150 & n6308 ) | ( ~n6307 & n6308 ) ;
  assign n6310 = ( n6171 & n6262 ) | ( n6171 & n6309 ) | ( n6262 & n6309 ) ;
  assign n6311 = ( ~n6171 & n6262 ) | ( ~n6171 & n6309 ) | ( n6262 & n6309 ) ;
  assign n6312 = ( n6171 & ~n6310 ) | ( n6171 & n6311 ) | ( ~n6310 & n6311 ) ;
  assign n6313 = ( n6222 & n6225 ) | ( n6222 & n6312 ) | ( n6225 & n6312 ) ;
  assign n6314 = ( n6222 & ~n6225 ) | ( n6222 & n6312 ) | ( ~n6225 & n6312 ) ;
  assign n6315 = ( n6225 & ~n6313 ) | ( n6225 & n6314 ) | ( ~n6313 & n6314 ) ;
  assign n6316 = ( n6240 & n6288 ) | ( n6240 & n6298 ) | ( n6288 & n6298 ) ;
  assign n6317 = ( n6240 & ~n6288 ) | ( n6240 & n6298 ) | ( ~n6288 & n6298 ) ;
  assign n6318 = ( n6288 & ~n6316 ) | ( n6288 & n6317 ) | ( ~n6316 & n6317 ) ;
  assign n6319 = ( n6282 & n6302 ) | ( n6282 & n6318 ) | ( n6302 & n6318 ) ;
  assign n6320 = ( n6282 & n6302 ) | ( n6282 & ~n6318 ) | ( n6302 & ~n6318 ) ;
  assign n6321 = ( n6318 & ~n6319 ) | ( n6318 & n6320 ) | ( ~n6319 & n6320 ) ;
  assign n6322 = ( n6254 & ~n6304 ) | ( n6254 & n6321 ) | ( ~n6304 & n6321 ) ;
  assign n6323 = ( n6254 & n6304 ) | ( n6254 & n6321 ) | ( n6304 & n6321 ) ;
  assign n6324 = ( n6304 & n6322 ) | ( n6304 & ~n6323 ) | ( n6322 & ~n6323 ) ;
  assign n6325 = ( n6258 & n6307 ) | ( n6258 & ~n6324 ) | ( n6307 & ~n6324 ) ;
  assign n6326 = ( n6258 & n6307 ) | ( n6258 & n6324 ) | ( n6307 & n6324 ) ;
  assign n6327 = ( n6324 & n6325 ) | ( n6324 & ~n6326 ) | ( n6325 & ~n6326 ) ;
  assign n6328 = x26 & x58 ;
  assign n6329 = x31 & x53 ;
  assign n6330 = x32 & x52 ;
  assign n6331 = ( ~n6328 & n6329 ) | ( ~n6328 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6332 = ( n6328 & n6329 ) | ( n6328 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6333 = ( n6328 & n6331 ) | ( n6328 & ~n6332 ) | ( n6331 & ~n6332 ) ;
  assign n6334 = ( ~n6233 & n6267 ) | ( ~n6233 & n6333 ) | ( n6267 & n6333 ) ;
  assign n6335 = ( n6233 & n6267 ) | ( n6233 & n6333 ) | ( n6267 & n6333 ) ;
  assign n6336 = ( n6233 & n6334 ) | ( n6233 & ~n6335 ) | ( n6334 & ~n6335 ) ;
  assign n6337 = ( ~n6229 & n6242 ) | ( ~n6229 & n6336 ) | ( n6242 & n6336 ) ;
  assign n6338 = ( n6229 & n6242 ) | ( n6229 & n6336 ) | ( n6242 & n6336 ) ;
  assign n6339 = ( n6229 & n6337 ) | ( n6229 & ~n6338 ) | ( n6337 & ~n6338 ) ;
  assign n6340 = ( n6273 & n6279 ) | ( n6273 & ~n6294 ) | ( n6279 & ~n6294 ) ;
  assign n6341 = ( n6273 & n6279 ) | ( n6273 & n6294 ) | ( n6279 & n6294 ) ;
  assign n6342 = ( n6294 & n6340 ) | ( n6294 & ~n6341 ) | ( n6340 & ~n6341 ) ;
  assign n6343 = ( n6249 & n6252 ) | ( n6249 & n6342 ) | ( n6252 & n6342 ) ;
  assign n6344 = ( n6249 & n6252 ) | ( n6249 & ~n6342 ) | ( n6252 & ~n6342 ) ;
  assign n6345 = ( n6342 & ~n6343 ) | ( n6342 & n6344 ) | ( ~n6343 & n6344 ) ;
  assign n6346 = x21 & x63 ;
  assign n6347 = x22 & x62 ;
  assign n6348 = x23 & x61 ;
  assign n6349 = ( ~n6346 & n6347 ) | ( ~n6346 & n6348 ) | ( n6347 & n6348 ) ;
  assign n6350 = ( n6346 & n6347 ) | ( n6346 & n6348 ) | ( n6347 & n6348 ) ;
  assign n6351 = ( n6346 & n6349 ) | ( n6346 & ~n6350 ) | ( n6349 & ~n6350 ) ;
  assign n6352 = x24 & x60 ;
  assign n6353 = x25 & x59 ;
  assign n6354 = x33 & x51 ;
  assign n6355 = ( ~n6352 & n6353 ) | ( ~n6352 & n6354 ) | ( n6353 & n6354 ) ;
  assign n6356 = ( n6352 & n6353 ) | ( n6352 & n6354 ) | ( n6353 & n6354 ) ;
  assign n6357 = ( n6352 & n6355 ) | ( n6352 & ~n6356 ) | ( n6355 & ~n6356 ) ;
  assign n6358 = x35 & x49 ;
  assign n6359 = x36 & x48 ;
  assign n6360 = x34 & x50 ;
  assign n6361 = ( ~n6358 & n6359 ) | ( ~n6358 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6362 = ( n6358 & n6359 ) | ( n6358 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6363 = ( n6358 & n6361 ) | ( n6358 & ~n6362 ) | ( n6361 & ~n6362 ) ;
  assign n6364 = ( ~n6351 & n6357 ) | ( ~n6351 & n6363 ) | ( n6357 & n6363 ) ;
  assign n6365 = ( n6351 & n6357 ) | ( n6351 & n6363 ) | ( n6357 & n6363 ) ;
  assign n6366 = ( n6351 & n6364 ) | ( n6351 & ~n6365 ) | ( n6364 & ~n6365 ) ;
  assign n6367 = x38 & x46 ;
  assign n6368 = x28 & x56 ;
  assign n6369 = ( ~n3291 & n6367 ) | ( ~n3291 & n6368 ) | ( n6367 & n6368 ) ;
  assign n6370 = ( n3291 & n6367 ) | ( n3291 & n6368 ) | ( n6367 & n6368 ) ;
  assign n6371 = ( n3291 & n6369 ) | ( n3291 & ~n6370 ) | ( n6369 & ~n6370 ) ;
  assign n6372 = x27 & x57 ;
  assign n6373 = x37 & x47 ;
  assign n6374 = x30 & x54 ;
  assign n6375 = ( ~n6372 & n6373 ) | ( ~n6372 & n6374 ) | ( n6373 & n6374 ) ;
  assign n6376 = ( n6372 & n6373 ) | ( n6372 & n6374 ) | ( n6373 & n6374 ) ;
  assign n6377 = ( n6372 & n6375 ) | ( n6372 & ~n6376 ) | ( n6375 & ~n6376 ) ;
  assign n6378 = x39 & x45 ;
  assign n6379 = x41 & x43 ;
  assign n6380 = x40 & x44 ;
  assign n6381 = ( ~n6378 & n6379 ) | ( ~n6378 & n6380 ) | ( n6379 & n6380 ) ;
  assign n6382 = ( n6378 & n6379 ) | ( n6378 & n6380 ) | ( n6379 & n6380 ) ;
  assign n6383 = ( n6378 & n6381 ) | ( n6378 & ~n6382 ) | ( n6381 & ~n6382 ) ;
  assign n6384 = ( ~n6371 & n6377 ) | ( ~n6371 & n6383 ) | ( n6377 & n6383 ) ;
  assign n6385 = ( n6371 & n6377 ) | ( n6371 & n6383 ) | ( n6377 & n6383 ) ;
  assign n6386 = ( n6371 & n6384 ) | ( n6371 & ~n6385 ) | ( n6384 & ~n6385 ) ;
  assign n6387 = ( n6345 & n6366 ) | ( n6345 & n6386 ) | ( n6366 & n6386 ) ;
  assign n6388 = ( ~n6345 & n6366 ) | ( ~n6345 & n6386 ) | ( n6366 & n6386 ) ;
  assign n6389 = ( n6345 & ~n6387 ) | ( n6345 & n6388 ) | ( ~n6387 & n6388 ) ;
  assign n6390 = ( n6245 & n6339 ) | ( n6245 & n6389 ) | ( n6339 & n6389 ) ;
  assign n6391 = ( ~n6245 & n6339 ) | ( ~n6245 & n6389 ) | ( n6339 & n6389 ) ;
  assign n6392 = ( n6245 & ~n6390 ) | ( n6245 & n6391 ) | ( ~n6390 & n6391 ) ;
  assign n6393 = ( n6260 & n6327 ) | ( n6260 & n6392 ) | ( n6327 & n6392 ) ;
  assign n6394 = ( ~n6260 & n6327 ) | ( ~n6260 & n6392 ) | ( n6327 & n6392 ) ;
  assign n6395 = ( n6260 & ~n6393 ) | ( n6260 & n6394 ) | ( ~n6393 & n6394 ) ;
  assign n6396 = ( n6310 & n6313 ) | ( n6310 & n6395 ) | ( n6313 & n6395 ) ;
  assign n6397 = ( n6310 & ~n6313 ) | ( n6310 & n6395 ) | ( ~n6313 & n6395 ) ;
  assign n6398 = ( n6313 & ~n6396 ) | ( n6313 & n6397 ) | ( ~n6396 & n6397 ) ;
  assign n6399 = x40 & x45 ;
  assign n6400 = x41 & x44 ;
  assign n6401 = x39 & x46 ;
  assign n6402 = ( ~n6399 & n6400 ) | ( ~n6399 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6403 = ( n6399 & n6400 ) | ( n6399 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6404 = ( n6399 & n6402 ) | ( n6399 & ~n6403 ) | ( n6402 & ~n6403 ) ;
  assign n6405 = x35 & x50 ;
  assign n6406 = x22 & x63 ;
  assign n6407 = x28 & x57 ;
  assign n6408 = ( ~n6405 & n6406 ) | ( ~n6405 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6409 = ( n6405 & n6406 ) | ( n6405 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6410 = ( n6405 & n6408 ) | ( n6405 & ~n6409 ) | ( n6408 & ~n6409 ) ;
  assign n6411 = x32 & x53 ;
  assign n6412 = x33 & x52 ;
  assign n6413 = x34 & x51 ;
  assign n6414 = ( ~n6411 & n6412 ) | ( ~n6411 & n6413 ) | ( n6412 & n6413 ) ;
  assign n6415 = ( n6411 & n6412 ) | ( n6411 & n6413 ) | ( n6412 & n6413 ) ;
  assign n6416 = ( n6411 & n6414 ) | ( n6411 & ~n6415 ) | ( n6414 & ~n6415 ) ;
  assign n6417 = ( ~n6404 & n6410 ) | ( ~n6404 & n6416 ) | ( n6410 & n6416 ) ;
  assign n6418 = ( n6404 & n6410 ) | ( n6404 & n6416 ) | ( n6410 & n6416 ) ;
  assign n6419 = ( n6404 & n6417 ) | ( n6404 & ~n6418 ) | ( n6417 & ~n6418 ) ;
  assign n6420 = x38 & x47 ;
  assign n6421 = x37 & x48 ;
  assign n6422 = x36 & x49 ;
  assign n6423 = ( ~n6420 & n6421 ) | ( ~n6420 & n6422 ) | ( n6421 & n6422 ) ;
  assign n6424 = ( n6420 & n6421 ) | ( n6420 & n6422 ) | ( n6421 & n6422 ) ;
  assign n6425 = ( n6420 & n6423 ) | ( n6420 & ~n6424 ) | ( n6423 & ~n6424 ) ;
  assign n6426 = x30 & x55 ;
  assign n6427 = x31 & x54 ;
  assign n6428 = ( ~n3341 & n6426 ) | ( ~n3341 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6429 = ( n3341 & n6426 ) | ( n3341 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6430 = ( n3341 & n6428 ) | ( n3341 & ~n6429 ) | ( n6428 & ~n6429 ) ;
  assign n6431 = x23 & x62 ;
  assign n6432 = x42 & x43 ;
  assign n6433 = ( x43 & n6431 ) | ( x43 & n6432 ) | ( n6431 & n6432 ) ;
  assign n6434 = ( x43 & ~n6431 ) | ( x43 & n6432 ) | ( ~n6431 & n6432 ) ;
  assign n6435 = ( n6431 & ~n6433 ) | ( n6431 & n6434 ) | ( ~n6433 & n6434 ) ;
  assign n6436 = ( ~n6425 & n6430 ) | ( ~n6425 & n6435 ) | ( n6430 & n6435 ) ;
  assign n6437 = ( n6425 & n6430 ) | ( n6425 & n6435 ) | ( n6430 & n6435 ) ;
  assign n6438 = ( n6425 & n6436 ) | ( n6425 & ~n6437 ) | ( n6436 & ~n6437 ) ;
  assign n6439 = ( n6319 & n6419 ) | ( n6319 & n6438 ) | ( n6419 & n6438 ) ;
  assign n6440 = ( ~n6319 & n6419 ) | ( ~n6319 & n6438 ) | ( n6419 & n6438 ) ;
  assign n6441 = ( n6319 & ~n6439 ) | ( n6319 & n6440 ) | ( ~n6439 & n6440 ) ;
  assign n6442 = x26 & x59 ;
  assign n6443 = x27 & x58 ;
  assign n6444 = x25 & x60 ;
  assign n6445 = ( ~n6442 & n6443 ) | ( ~n6442 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6446 = ( n6442 & n6443 ) | ( n6442 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6447 = ( n6442 & n6445 ) | ( n6442 & ~n6446 ) | ( n6445 & ~n6446 ) ;
  assign n6448 = ( n6332 & n6376 ) | ( n6332 & ~n6447 ) | ( n6376 & ~n6447 ) ;
  assign n6449 = ( n6332 & n6376 ) | ( n6332 & n6447 ) | ( n6376 & n6447 ) ;
  assign n6450 = ( n6447 & n6448 ) | ( n6447 & ~n6449 ) | ( n6448 & ~n6449 ) ;
  assign n6451 = x24 & x61 ;
  assign n6452 = ( n6370 & n6382 ) | ( n6370 & n6451 ) | ( n6382 & n6451 ) ;
  assign n6453 = ( ~n6370 & n6382 ) | ( ~n6370 & n6451 ) | ( n6382 & n6451 ) ;
  assign n6454 = ( n6370 & ~n6452 ) | ( n6370 & n6453 ) | ( ~n6452 & n6453 ) ;
  assign n6455 = ( n6343 & n6450 ) | ( n6343 & n6454 ) | ( n6450 & n6454 ) ;
  assign n6456 = ( ~n6343 & n6450 ) | ( ~n6343 & n6454 ) | ( n6450 & n6454 ) ;
  assign n6457 = ( n6343 & ~n6455 ) | ( n6343 & n6456 ) | ( ~n6455 & n6456 ) ;
  assign n6458 = ( ~n6350 & n6356 ) | ( ~n6350 & n6362 ) | ( n6356 & n6362 ) ;
  assign n6459 = ( n6350 & n6356 ) | ( n6350 & n6362 ) | ( n6356 & n6362 ) ;
  assign n6460 = ( n6350 & n6458 ) | ( n6350 & ~n6459 ) | ( n6458 & ~n6459 ) ;
  assign n6461 = ( n6365 & n6385 ) | ( n6365 & n6460 ) | ( n6385 & n6460 ) ;
  assign n6462 = ( ~n6365 & n6385 ) | ( ~n6365 & n6460 ) | ( n6385 & n6460 ) ;
  assign n6463 = ( n6365 & ~n6461 ) | ( n6365 & n6462 ) | ( ~n6461 & n6462 ) ;
  assign n6464 = ( ~n6441 & n6457 ) | ( ~n6441 & n6463 ) | ( n6457 & n6463 ) ;
  assign n6465 = ( n6441 & n6457 ) | ( n6441 & n6463 ) | ( n6457 & n6463 ) ;
  assign n6466 = ( n6441 & n6464 ) | ( n6441 & ~n6465 ) | ( n6464 & ~n6465 ) ;
  assign n6467 = ( n6316 & ~n6335 ) | ( n6316 & n6341 ) | ( ~n6335 & n6341 ) ;
  assign n6468 = ( n6316 & n6335 ) | ( n6316 & n6341 ) | ( n6335 & n6341 ) ;
  assign n6469 = ( n6335 & n6467 ) | ( n6335 & ~n6468 ) | ( n6467 & ~n6468 ) ;
  assign n6470 = ( n6338 & n6387 ) | ( n6338 & n6469 ) | ( n6387 & n6469 ) ;
  assign n6471 = ( ~n6338 & n6387 ) | ( ~n6338 & n6469 ) | ( n6387 & n6469 ) ;
  assign n6472 = ( n6338 & ~n6470 ) | ( n6338 & n6471 ) | ( ~n6470 & n6471 ) ;
  assign n6473 = ( n6323 & n6390 ) | ( n6323 & n6472 ) | ( n6390 & n6472 ) ;
  assign n6474 = ( n6323 & ~n6390 ) | ( n6323 & n6472 ) | ( ~n6390 & n6472 ) ;
  assign n6475 = ( n6390 & ~n6473 ) | ( n6390 & n6474 ) | ( ~n6473 & n6474 ) ;
  assign n6476 = ( n6326 & n6466 ) | ( n6326 & n6475 ) | ( n6466 & n6475 ) ;
  assign n6477 = ( ~n6326 & n6466 ) | ( ~n6326 & n6475 ) | ( n6466 & n6475 ) ;
  assign n6478 = ( n6326 & ~n6476 ) | ( n6326 & n6477 ) | ( ~n6476 & n6477 ) ;
  assign n6479 = ( n6393 & n6396 ) | ( n6393 & n6478 ) | ( n6396 & n6478 ) ;
  assign n6480 = ( n6393 & ~n6396 ) | ( n6393 & n6478 ) | ( ~n6396 & n6478 ) ;
  assign n6481 = ( n6396 & ~n6479 ) | ( n6396 & n6480 ) | ( ~n6479 & n6480 ) ;
  assign n6482 = x25 & x61 ;
  assign n6483 = x24 & x62 ;
  assign n6484 = ( ~n6433 & n6482 ) | ( ~n6433 & n6483 ) | ( n6482 & n6483 ) ;
  assign n6485 = ( n6433 & n6482 ) | ( n6433 & n6483 ) | ( n6482 & n6483 ) ;
  assign n6486 = ( n6433 & n6484 ) | ( n6433 & ~n6485 ) | ( n6484 & ~n6485 ) ;
  assign n6487 = ( n6452 & n6459 ) | ( n6452 & ~n6486 ) | ( n6459 & ~n6486 ) ;
  assign n6488 = ( n6452 & n6459 ) | ( n6452 & n6486 ) | ( n6459 & n6486 ) ;
  assign n6489 = ( n6486 & n6487 ) | ( n6486 & ~n6488 ) | ( n6487 & ~n6488 ) ;
  assign n6490 = ( n6439 & n6455 ) | ( n6439 & n6489 ) | ( n6455 & n6489 ) ;
  assign n6491 = ( ~n6439 & n6455 ) | ( ~n6439 & n6489 ) | ( n6455 & n6489 ) ;
  assign n6492 = ( n6439 & ~n6490 ) | ( n6439 & n6491 ) | ( ~n6490 & n6491 ) ;
  assign n6493 = ( n6465 & n6470 ) | ( n6465 & n6492 ) | ( n6470 & n6492 ) ;
  assign n6494 = ( n6465 & ~n6470 ) | ( n6465 & n6492 ) | ( ~n6470 & n6492 ) ;
  assign n6495 = ( n6470 & ~n6493 ) | ( n6470 & n6494 ) | ( ~n6493 & n6494 ) ;
  assign n6496 = ( n6403 & ~n6424 ) | ( n6403 & n6429 ) | ( ~n6424 & n6429 ) ;
  assign n6497 = ( n6403 & n6424 ) | ( n6403 & n6429 ) | ( n6424 & n6429 ) ;
  assign n6498 = ( n6424 & n6496 ) | ( n6424 & ~n6497 ) | ( n6496 & ~n6497 ) ;
  assign n6499 = ( n6409 & n6415 ) | ( n6409 & ~n6446 ) | ( n6415 & ~n6446 ) ;
  assign n6500 = ( n6409 & n6415 ) | ( n6409 & n6446 ) | ( n6415 & n6446 ) ;
  assign n6501 = ( n6446 & n6499 ) | ( n6446 & ~n6500 ) | ( n6499 & ~n6500 ) ;
  assign n6502 = ( n6468 & n6498 ) | ( n6468 & n6501 ) | ( n6498 & n6501 ) ;
  assign n6503 = ( ~n6468 & n6498 ) | ( ~n6468 & n6501 ) | ( n6498 & n6501 ) ;
  assign n6504 = ( n6468 & ~n6502 ) | ( n6468 & n6503 ) | ( ~n6502 & n6503 ) ;
  assign n6505 = ( n6418 & n6437 ) | ( n6418 & ~n6449 ) | ( n6437 & ~n6449 ) ;
  assign n6506 = ( n6418 & n6437 ) | ( n6418 & n6449 ) | ( n6437 & n6449 ) ;
  assign n6507 = ( n6449 & n6505 ) | ( n6449 & ~n6506 ) | ( n6505 & ~n6506 ) ;
  assign n6508 = x29 & x57 ;
  assign n6509 = x31 & x55 ;
  assign n6510 = x38 & x48 ;
  assign n6511 = ( ~n6508 & n6509 ) | ( ~n6508 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6512 = ( n6508 & n6509 ) | ( n6508 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6513 = ( n6508 & n6511 ) | ( n6508 & ~n6512 ) | ( n6511 & ~n6512 ) ;
  assign n6514 = x35 & x51 ;
  assign n6515 = x33 & x53 ;
  assign n6516 = x34 & x52 ;
  assign n6517 = ( ~n6514 & n6515 ) | ( ~n6514 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6518 = ( n6514 & n6515 ) | ( n6514 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6519 = ( n6514 & n6517 ) | ( n6514 & ~n6518 ) | ( n6517 & ~n6518 ) ;
  assign n6520 = x37 & x49 ;
  assign n6521 = x23 & x63 ;
  assign n6522 = x36 & x50 ;
  assign n6523 = ( ~n6520 & n6521 ) | ( ~n6520 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6524 = ( n6520 & n6521 ) | ( n6520 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6525 = ( n6520 & n6523 ) | ( n6520 & ~n6524 ) | ( n6523 & ~n6524 ) ;
  assign n6526 = ( ~n6513 & n6519 ) | ( ~n6513 & n6525 ) | ( n6519 & n6525 ) ;
  assign n6527 = ( n6513 & n6519 ) | ( n6513 & n6525 ) | ( n6519 & n6525 ) ;
  assign n6528 = ( n6513 & n6526 ) | ( n6513 & ~n6527 ) | ( n6526 & ~n6527 ) ;
  assign n6529 = x30 & x56 ;
  assign n6530 = x39 & x47 ;
  assign n6531 = x40 & x46 ;
  assign n6532 = ( ~n6529 & n6530 ) | ( ~n6529 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6533 = ( n6529 & n6530 ) | ( n6529 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6534 = ( n6529 & n6532 ) | ( n6529 & ~n6533 ) | ( n6532 & ~n6533 ) ;
  assign n6535 = x28 & x58 ;
  assign n6536 = x26 & x60 ;
  assign n6537 = x27 & x59 ;
  assign n6538 = ( ~n6535 & n6536 ) | ( ~n6535 & n6537 ) | ( n6536 & n6537 ) ;
  assign n6539 = ( n6535 & n6536 ) | ( n6535 & n6537 ) | ( n6536 & n6537 ) ;
  assign n6540 = ( n6535 & n6538 ) | ( n6535 & ~n6539 ) | ( n6538 & ~n6539 ) ;
  assign n6541 = x42 & x44 ;
  assign n6542 = x41 & x45 ;
  assign n6543 = x32 & x54 ;
  assign n6544 = ( ~n6541 & n6542 ) | ( ~n6541 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6545 = ( n6541 & n6542 ) | ( n6541 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6546 = ( n6541 & n6544 ) | ( n6541 & ~n6545 ) | ( n6544 & ~n6545 ) ;
  assign n6547 = ( ~n6534 & n6540 ) | ( ~n6534 & n6546 ) | ( n6540 & n6546 ) ;
  assign n6548 = ( n6534 & n6540 ) | ( n6534 & n6546 ) | ( n6540 & n6546 ) ;
  assign n6549 = ( n6534 & n6547 ) | ( n6534 & ~n6548 ) | ( n6547 & ~n6548 ) ;
  assign n6550 = ( n6461 & n6528 ) | ( n6461 & n6549 ) | ( n6528 & n6549 ) ;
  assign n6551 = ( ~n6461 & n6528 ) | ( ~n6461 & n6549 ) | ( n6528 & n6549 ) ;
  assign n6552 = ( n6461 & ~n6550 ) | ( n6461 & n6551 ) | ( ~n6550 & n6551 ) ;
  assign n6553 = ( ~n6504 & n6507 ) | ( ~n6504 & n6552 ) | ( n6507 & n6552 ) ;
  assign n6554 = ( n6504 & n6507 ) | ( n6504 & n6552 ) | ( n6507 & n6552 ) ;
  assign n6555 = ( n6504 & n6553 ) | ( n6504 & ~n6554 ) | ( n6553 & ~n6554 ) ;
  assign n6556 = ( n6473 & ~n6495 ) | ( n6473 & n6555 ) | ( ~n6495 & n6555 ) ;
  assign n6557 = ( n6473 & n6495 ) | ( n6473 & n6555 ) | ( n6495 & n6555 ) ;
  assign n6558 = ( n6495 & n6556 ) | ( n6495 & ~n6557 ) | ( n6556 & ~n6557 ) ;
  assign n6559 = ( n6476 & n6479 ) | ( n6476 & n6558 ) | ( n6479 & n6558 ) ;
  assign n6560 = ( n6476 & ~n6479 ) | ( n6476 & n6558 ) | ( ~n6479 & n6558 ) ;
  assign n6561 = ( n6479 & ~n6559 ) | ( n6479 & n6560 ) | ( ~n6559 & n6560 ) ;
  assign n6562 = x40 & x47 ;
  assign n6563 = x33 & x54 ;
  assign n6564 = x31 & x56 ;
  assign n6565 = ( ~n6562 & n6563 ) | ( ~n6562 & n6564 ) | ( n6563 & n6564 ) ;
  assign n6566 = ( n6562 & n6563 ) | ( n6562 & n6564 ) | ( n6563 & n6564 ) ;
  assign n6567 = ( n6562 & n6565 ) | ( n6562 & ~n6566 ) | ( n6565 & ~n6566 ) ;
  assign n6568 = x25 & x62 ;
  assign n6569 = x43 & x44 ;
  assign n6570 = ( x44 & n6568 ) | ( x44 & n6569 ) | ( n6568 & n6569 ) ;
  assign n6571 = ( x44 & ~n6568 ) | ( x44 & n6569 ) | ( ~n6568 & n6569 ) ;
  assign n6572 = ( n6568 & ~n6570 ) | ( n6568 & n6571 ) | ( ~n6570 & n6571 ) ;
  assign n6573 = ( ~n6500 & n6567 ) | ( ~n6500 & n6572 ) | ( n6567 & n6572 ) ;
  assign n6574 = ( n6500 & n6567 ) | ( n6500 & n6572 ) | ( n6567 & n6572 ) ;
  assign n6575 = ( n6500 & n6573 ) | ( n6500 & ~n6574 ) | ( n6573 & ~n6574 ) ;
  assign n6576 = x34 & x53 ;
  assign n6577 = x28 & x59 ;
  assign n6578 = ( ~n3535 & n6576 ) | ( ~n3535 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6579 = ( n3535 & n6576 ) | ( n3535 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6580 = ( n3535 & n6578 ) | ( n3535 & ~n6579 ) | ( n6578 & ~n6579 ) ;
  assign n6581 = x35 & x52 ;
  assign n6582 = x29 & x58 ;
  assign n6583 = x36 & x51 ;
  assign n6584 = ( ~n6581 & n6582 ) | ( ~n6581 & n6583 ) | ( n6582 & n6583 ) ;
  assign n6585 = ( n6581 & n6582 ) | ( n6581 & n6583 ) | ( n6582 & n6583 ) ;
  assign n6586 = ( n6581 & n6584 ) | ( n6581 & ~n6585 ) | ( n6584 & ~n6585 ) ;
  assign n6587 = ( ~n6485 & n6580 ) | ( ~n6485 & n6586 ) | ( n6580 & n6586 ) ;
  assign n6588 = ( n6485 & n6580 ) | ( n6485 & n6586 ) | ( n6580 & n6586 ) ;
  assign n6589 = ( n6485 & n6587 ) | ( n6485 & ~n6588 ) | ( n6587 & ~n6588 ) ;
  assign n6590 = x37 & x50 ;
  assign n6591 = x39 & x48 ;
  assign n6592 = x38 & x49 ;
  assign n6593 = ( ~n6590 & n6591 ) | ( ~n6590 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6594 = ( n6590 & n6591 ) | ( n6590 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6595 = ( n6590 & n6593 ) | ( n6590 & ~n6594 ) | ( n6593 & ~n6594 ) ;
  assign n6596 = x27 & x60 ;
  assign n6597 = x24 & x63 ;
  assign n6598 = x26 & x61 ;
  assign n6599 = ( ~n6596 & n6597 ) | ( ~n6596 & n6598 ) | ( n6597 & n6598 ) ;
  assign n6600 = ( n6596 & n6597 ) | ( n6596 & n6598 ) | ( n6597 & n6598 ) ;
  assign n6601 = ( n6596 & n6599 ) | ( n6596 & ~n6600 ) | ( n6599 & ~n6600 ) ;
  assign n6602 = x32 & x55 ;
  assign n6603 = x41 & x46 ;
  assign n6604 = x42 & x45 ;
  assign n6605 = ( ~n6602 & n6603 ) | ( ~n6602 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6606 = ( n6602 & n6603 ) | ( n6602 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6607 = ( n6602 & n6605 ) | ( n6602 & ~n6606 ) | ( n6605 & ~n6606 ) ;
  assign n6608 = ( ~n6595 & n6601 ) | ( ~n6595 & n6607 ) | ( n6601 & n6607 ) ;
  assign n6609 = ( n6595 & n6601 ) | ( n6595 & n6607 ) | ( n6601 & n6607 ) ;
  assign n6610 = ( n6595 & n6608 ) | ( n6595 & ~n6609 ) | ( n6608 & ~n6609 ) ;
  assign n6611 = ( ~n6575 & n6589 ) | ( ~n6575 & n6610 ) | ( n6589 & n6610 ) ;
  assign n6612 = ( n6575 & n6589 ) | ( n6575 & n6610 ) | ( n6589 & n6610 ) ;
  assign n6613 = ( n6575 & n6611 ) | ( n6575 & ~n6612 ) | ( n6611 & ~n6612 ) ;
  assign n6614 = ( n6518 & ~n6524 ) | ( n6518 & n6539 ) | ( ~n6524 & n6539 ) ;
  assign n6615 = ( n6518 & n6524 ) | ( n6518 & n6539 ) | ( n6524 & n6539 ) ;
  assign n6616 = ( n6524 & n6614 ) | ( n6524 & ~n6615 ) | ( n6614 & ~n6615 ) ;
  assign n6617 = ( ~n6512 & n6533 ) | ( ~n6512 & n6545 ) | ( n6533 & n6545 ) ;
  assign n6618 = ( n6512 & n6533 ) | ( n6512 & n6545 ) | ( n6533 & n6545 ) ;
  assign n6619 = ( n6512 & n6617 ) | ( n6512 & ~n6618 ) | ( n6617 & ~n6618 ) ;
  assign n6620 = ( n6488 & n6616 ) | ( n6488 & n6619 ) | ( n6616 & n6619 ) ;
  assign n6621 = ( ~n6488 & n6616 ) | ( ~n6488 & n6619 ) | ( n6616 & n6619 ) ;
  assign n6622 = ( n6488 & ~n6620 ) | ( n6488 & n6621 ) | ( ~n6620 & n6621 ) ;
  assign n6623 = ( n6502 & n6506 ) | ( n6502 & n6622 ) | ( n6506 & n6622 ) ;
  assign n6624 = ( ~n6502 & n6506 ) | ( ~n6502 & n6622 ) | ( n6506 & n6622 ) ;
  assign n6625 = ( n6502 & ~n6623 ) | ( n6502 & n6624 ) | ( ~n6623 & n6624 ) ;
  assign n6626 = ( n6554 & n6613 ) | ( n6554 & n6625 ) | ( n6613 & n6625 ) ;
  assign n6627 = ( ~n6554 & n6613 ) | ( ~n6554 & n6625 ) | ( n6613 & n6625 ) ;
  assign n6628 = ( n6554 & ~n6626 ) | ( n6554 & n6627 ) | ( ~n6626 & n6627 ) ;
  assign n6629 = ( n6497 & ~n6527 ) | ( n6497 & n6548 ) | ( ~n6527 & n6548 ) ;
  assign n6630 = ( n6497 & n6527 ) | ( n6497 & n6548 ) | ( n6527 & n6548 ) ;
  assign n6631 = ( n6527 & n6629 ) | ( n6527 & ~n6630 ) | ( n6629 & ~n6630 ) ;
  assign n6632 = ( n6490 & n6550 ) | ( n6490 & n6631 ) | ( n6550 & n6631 ) ;
  assign n6633 = ( ~n6490 & n6550 ) | ( ~n6490 & n6631 ) | ( n6550 & n6631 ) ;
  assign n6634 = ( n6490 & ~n6632 ) | ( n6490 & n6633 ) | ( ~n6632 & n6633 ) ;
  assign n6635 = ( ~n6493 & n6628 ) | ( ~n6493 & n6634 ) | ( n6628 & n6634 ) ;
  assign n6636 = ( n6493 & n6628 ) | ( n6493 & n6634 ) | ( n6628 & n6634 ) ;
  assign n6637 = ( n6493 & n6635 ) | ( n6493 & ~n6636 ) | ( n6635 & ~n6636 ) ;
  assign n6638 = ( n6557 & ~n6559 ) | ( n6557 & n6637 ) | ( ~n6559 & n6637 ) ;
  assign n6639 = ( n6557 & n6559 ) | ( n6557 & n6637 ) | ( n6559 & n6637 ) ;
  assign n6640 = ( n6559 & n6638 ) | ( n6559 & ~n6639 ) | ( n6638 & ~n6639 ) ;
  assign n6641 = x43 & x45 ;
  assign n6642 = x34 & x54 ;
  assign n6643 = x33 & x55 ;
  assign n6644 = ( ~n6641 & n6642 ) | ( ~n6641 & n6643 ) | ( n6642 & n6643 ) ;
  assign n6645 = ( n6641 & n6642 ) | ( n6641 & n6643 ) | ( n6642 & n6643 ) ;
  assign n6646 = ( n6641 & n6644 ) | ( n6641 & ~n6645 ) | ( n6644 & ~n6645 ) ;
  assign n6647 = ( n6566 & n6585 ) | ( n6566 & ~n6646 ) | ( n6585 & ~n6646 ) ;
  assign n6648 = ( n6566 & n6585 ) | ( n6566 & n6646 ) | ( n6585 & n6646 ) ;
  assign n6649 = ( n6646 & n6647 ) | ( n6646 & ~n6648 ) | ( n6647 & ~n6648 ) ;
  assign n6650 = ( n6579 & ~n6594 ) | ( n6579 & n6600 ) | ( ~n6594 & n6600 ) ;
  assign n6651 = ( n6579 & n6594 ) | ( n6579 & n6600 ) | ( n6594 & n6600 ) ;
  assign n6652 = ( n6594 & n6650 ) | ( n6594 & ~n6651 ) | ( n6650 & ~n6651 ) ;
  assign n6653 = ( n6574 & n6649 ) | ( n6574 & n6652 ) | ( n6649 & n6652 ) ;
  assign n6654 = ( ~n6574 & n6649 ) | ( ~n6574 & n6652 ) | ( n6649 & n6652 ) ;
  assign n6655 = ( n6574 & ~n6653 ) | ( n6574 & n6654 ) | ( ~n6653 & n6654 ) ;
  assign n6656 = ( n6620 & n6630 ) | ( n6620 & n6655 ) | ( n6630 & n6655 ) ;
  assign n6657 = ( n6620 & n6630 ) | ( n6620 & ~n6655 ) | ( n6630 & ~n6655 ) ;
  assign n6658 = ( n6655 & ~n6656 ) | ( n6655 & n6657 ) | ( ~n6656 & n6657 ) ;
  assign n6659 = x39 & x49 ;
  assign n6660 = x29 & x59 ;
  assign n6661 = x38 & x50 ;
  assign n6662 = ( ~n6659 & n6660 ) | ( ~n6659 & n6661 ) | ( n6660 & n6661 ) ;
  assign n6663 = ( n6659 & n6660 ) | ( n6659 & n6661 ) | ( n6660 & n6661 ) ;
  assign n6664 = ( n6659 & n6662 ) | ( n6659 & ~n6663 ) | ( n6662 & ~n6663 ) ;
  assign n6665 = x40 & x48 ;
  assign n6666 = x32 & x56 ;
  assign n6667 = ( n3666 & ~n6665 ) | ( n3666 & n6666 ) | ( ~n6665 & n6666 ) ;
  assign n6668 = ( n3666 & n6665 ) | ( n3666 & n6666 ) | ( n6665 & n6666 ) ;
  assign n6669 = ( n6665 & n6667 ) | ( n6665 & ~n6668 ) | ( n6667 & ~n6668 ) ;
  assign n6670 = ( ~n6618 & n6664 ) | ( ~n6618 & n6669 ) | ( n6664 & n6669 ) ;
  assign n6671 = ( n6618 & n6664 ) | ( n6618 & n6669 ) | ( n6664 & n6669 ) ;
  assign n6672 = ( n6618 & n6670 ) | ( n6618 & ~n6671 ) | ( n6670 & ~n6671 ) ;
  assign n6673 = x25 & x63 ;
  assign n6674 = n6570 | n6673 ;
  assign n6675 = x44 & x63 ;
  assign n6676 = n4696 | n6568 ;
  assign n6677 = n6675 & n6676 ;
  assign n6678 = ( n6606 & n6674 ) | ( n6606 & n6677 ) | ( n6674 & n6677 ) ;
  assign n6679 = n6606 | n6674 ;
  assign n6680 = ( n6606 & ~n6674 ) | ( n6606 & n6677 ) | ( ~n6674 & n6677 ) ;
  assign n6681 = ( ~n6678 & n6679 ) | ( ~n6678 & n6680 ) | ( n6679 & n6680 ) ;
  assign n6682 = x37 & x51 ;
  assign n6683 = x35 & x53 ;
  assign n6684 = x36 & x52 ;
  assign n6685 = ( ~n6682 & n6683 ) | ( ~n6682 & n6684 ) | ( n6683 & n6684 ) ;
  assign n6686 = ( n6682 & n6683 ) | ( n6682 & n6684 ) | ( n6683 & n6684 ) ;
  assign n6687 = ( n6682 & n6685 ) | ( n6682 & ~n6686 ) | ( n6685 & ~n6686 ) ;
  assign n6688 = x42 & x46 ;
  assign n6689 = x31 & x57 ;
  assign n6690 = x41 & x47 ;
  assign n6691 = ( ~n6688 & n6689 ) | ( ~n6688 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6692 = ( n6688 & n6689 ) | ( n6688 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6693 = ( n6688 & n6691 ) | ( n6688 & ~n6692 ) | ( n6691 & ~n6692 ) ;
  assign n6694 = x26 & x62 ;
  assign n6695 = x27 & x61 ;
  assign n6696 = x28 & x60 ;
  assign n6697 = ( ~n6694 & n6695 ) | ( ~n6694 & n6696 ) | ( n6695 & n6696 ) ;
  assign n6698 = ( n6694 & n6695 ) | ( n6694 & n6696 ) | ( n6695 & n6696 ) ;
  assign n6699 = ( n6694 & n6697 ) | ( n6694 & ~n6698 ) | ( n6697 & ~n6698 ) ;
  assign n6700 = ( ~n6687 & n6693 ) | ( ~n6687 & n6699 ) | ( n6693 & n6699 ) ;
  assign n6701 = ( n6687 & n6693 ) | ( n6687 & n6699 ) | ( n6693 & n6699 ) ;
  assign n6702 = ( n6687 & n6700 ) | ( n6687 & ~n6701 ) | ( n6700 & ~n6701 ) ;
  assign n6703 = ( ~n6672 & n6681 ) | ( ~n6672 & n6702 ) | ( n6681 & n6702 ) ;
  assign n6704 = ( n6672 & n6681 ) | ( n6672 & n6702 ) | ( n6681 & n6702 ) ;
  assign n6705 = ( n6672 & n6703 ) | ( n6672 & ~n6704 ) | ( n6703 & ~n6704 ) ;
  assign n6706 = ( ~n6632 & n6658 ) | ( ~n6632 & n6705 ) | ( n6658 & n6705 ) ;
  assign n6707 = ( n6632 & n6658 ) | ( n6632 & n6705 ) | ( n6658 & n6705 ) ;
  assign n6708 = ( n6632 & n6706 ) | ( n6632 & ~n6707 ) | ( n6706 & ~n6707 ) ;
  assign n6709 = ( ~n6588 & n6609 ) | ( ~n6588 & n6615 ) | ( n6609 & n6615 ) ;
  assign n6710 = ( n6588 & n6609 ) | ( n6588 & n6615 ) | ( n6609 & n6615 ) ;
  assign n6711 = ( n6588 & n6709 ) | ( n6588 & ~n6710 ) | ( n6709 & ~n6710 ) ;
  assign n6712 = ( n6612 & n6623 ) | ( n6612 & n6711 ) | ( n6623 & n6711 ) ;
  assign n6713 = ( n6612 & n6623 ) | ( n6612 & ~n6711 ) | ( n6623 & ~n6711 ) ;
  assign n6714 = ( n6711 & ~n6712 ) | ( n6711 & n6713 ) | ( ~n6712 & n6713 ) ;
  assign n6715 = ( n6626 & ~n6708 ) | ( n6626 & n6714 ) | ( ~n6708 & n6714 ) ;
  assign n6716 = ( n6626 & n6708 ) | ( n6626 & n6714 ) | ( n6708 & n6714 ) ;
  assign n6717 = ( n6708 & n6715 ) | ( n6708 & ~n6716 ) | ( n6715 & ~n6716 ) ;
  assign n6718 = ( n6636 & n6639 ) | ( n6636 & n6717 ) | ( n6639 & n6717 ) ;
  assign n6719 = ( n6636 & ~n6639 ) | ( n6636 & n6717 ) | ( ~n6639 & n6717 ) ;
  assign n6720 = ( n6639 & ~n6718 ) | ( n6639 & n6719 ) | ( ~n6718 & n6719 ) ;
  assign n6721 = x26 & x63 ;
  assign n6722 = x39 & x50 ;
  assign n6723 = x40 & x49 ;
  assign n6724 = ( ~n6721 & n6722 ) | ( ~n6721 & n6723 ) | ( n6722 & n6723 ) ;
  assign n6725 = ( n6721 & n6722 ) | ( n6721 & n6723 ) | ( n6722 & n6723 ) ;
  assign n6726 = ( n6721 & n6724 ) | ( n6721 & ~n6725 ) | ( n6724 & ~n6725 ) ;
  assign n6727 = ( n6663 & n6692 ) | ( n6663 & ~n6726 ) | ( n6692 & ~n6726 ) ;
  assign n6728 = ( n6663 & n6692 ) | ( n6663 & n6726 ) | ( n6692 & n6726 ) ;
  assign n6729 = ( n6726 & n6727 ) | ( n6726 & ~n6728 ) | ( n6727 & ~n6728 ) ;
  assign n6730 = ( n6671 & n6701 ) | ( n6671 & n6729 ) | ( n6701 & n6729 ) ;
  assign n6731 = ( n6671 & n6701 ) | ( n6671 & ~n6729 ) | ( n6701 & ~n6729 ) ;
  assign n6732 = ( n6729 & ~n6730 ) | ( n6729 & n6731 ) | ( ~n6730 & n6731 ) ;
  assign n6733 = ( n6656 & n6704 ) | ( n6656 & n6732 ) | ( n6704 & n6732 ) ;
  assign n6734 = ( ~n6656 & n6704 ) | ( ~n6656 & n6732 ) | ( n6704 & n6732 ) ;
  assign n6735 = ( n6656 & ~n6733 ) | ( n6656 & n6734 ) | ( ~n6733 & n6734 ) ;
  assign n6736 = x28 & x61 ;
  assign n6737 = x29 & x60 ;
  assign n6738 = ( n6645 & n6736 ) | ( n6645 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6739 = ( ~n6645 & n6736 ) | ( ~n6645 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6740 = ( n6645 & ~n6738 ) | ( n6645 & n6739 ) | ( ~n6738 & n6739 ) ;
  assign n6741 = x43 & x46 ;
  assign n6742 = x42 & x47 ;
  assign n6743 = x34 & x55 ;
  assign n6744 = ( ~n6741 & n6742 ) | ( ~n6741 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6745 = ( n6741 & n6742 ) | ( n6741 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6746 = ( n6741 & n6744 ) | ( n6741 & ~n6745 ) | ( n6744 & ~n6745 ) ;
  assign n6747 = x27 & x62 ;
  assign n6748 = x44 & x45 ;
  assign n6749 = ( x45 & n6747 ) | ( x45 & n6748 ) | ( n6747 & n6748 ) ;
  assign n6750 = ( x45 & ~n6747 ) | ( x45 & n6748 ) | ( ~n6747 & n6748 ) ;
  assign n6751 = ( n6747 & ~n6749 ) | ( n6747 & n6750 ) | ( ~n6749 & n6750 ) ;
  assign n6752 = ( n6740 & n6746 ) | ( n6740 & n6751 ) | ( n6746 & n6751 ) ;
  assign n6753 = ( ~n6740 & n6746 ) | ( ~n6740 & n6751 ) | ( n6746 & n6751 ) ;
  assign n6754 = ( n6740 & ~n6752 ) | ( n6740 & n6753 ) | ( ~n6752 & n6753 ) ;
  assign n6755 = x37 & x52 ;
  assign n6756 = x38 & x51 ;
  assign n6757 = x36 & x53 ;
  assign n6758 = ( ~n6755 & n6756 ) | ( ~n6755 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6759 = ( n6755 & n6756 ) | ( n6755 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6760 = ( n6755 & n6758 ) | ( n6755 & ~n6759 ) | ( n6758 & ~n6759 ) ;
  assign n6761 = x35 & x54 ;
  assign n6762 = x33 & x56 ;
  assign n6763 = x41 & x48 ;
  assign n6764 = ( ~n6761 & n6762 ) | ( ~n6761 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6765 = ( n6761 & n6762 ) | ( n6761 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6766 = ( n6761 & n6764 ) | ( n6761 & ~n6765 ) | ( n6764 & ~n6765 ) ;
  assign n6767 = x31 & x58 ;
  assign n6768 = x30 & x59 ;
  assign n6769 = x32 & x57 ;
  assign n6770 = ( ~n6767 & n6768 ) | ( ~n6767 & n6769 ) | ( n6768 & n6769 ) ;
  assign n6771 = ( n6767 & n6768 ) | ( n6767 & n6769 ) | ( n6768 & n6769 ) ;
  assign n6772 = ( n6767 & n6770 ) | ( n6767 & ~n6771 ) | ( n6770 & ~n6771 ) ;
  assign n6773 = ( ~n6760 & n6766 ) | ( ~n6760 & n6772 ) | ( n6766 & n6772 ) ;
  assign n6774 = ( n6760 & n6766 ) | ( n6760 & n6772 ) | ( n6766 & n6772 ) ;
  assign n6775 = ( n6760 & n6773 ) | ( n6760 & ~n6774 ) | ( n6773 & ~n6774 ) ;
  assign n6776 = ( n6668 & ~n6686 ) | ( n6668 & n6698 ) | ( ~n6686 & n6698 ) ;
  assign n6777 = ( n6668 & n6686 ) | ( n6668 & n6698 ) | ( n6686 & n6698 ) ;
  assign n6778 = ( n6686 & n6776 ) | ( n6686 & ~n6777 ) | ( n6776 & ~n6777 ) ;
  assign n6779 = ( n6754 & n6775 ) | ( n6754 & n6778 ) | ( n6775 & n6778 ) ;
  assign n6780 = ( ~n6754 & n6775 ) | ( ~n6754 & n6778 ) | ( n6775 & n6778 ) ;
  assign n6781 = ( n6754 & ~n6779 ) | ( n6754 & n6780 ) | ( ~n6779 & n6780 ) ;
  assign n6782 = ( n6674 & n6678 ) | ( n6674 & ~n6681 ) | ( n6678 & ~n6681 ) ;
  assign n6783 = ( n6648 & n6651 ) | ( n6648 & n6782 ) | ( n6651 & n6782 ) ;
  assign n6784 = ( n6648 & n6651 ) | ( n6648 & ~n6782 ) | ( n6651 & ~n6782 ) ;
  assign n6785 = ( n6782 & ~n6783 ) | ( n6782 & n6784 ) | ( ~n6783 & n6784 ) ;
  assign n6786 = ( ~n6653 & n6710 ) | ( ~n6653 & n6785 ) | ( n6710 & n6785 ) ;
  assign n6787 = ( n6653 & n6710 ) | ( n6653 & n6785 ) | ( n6710 & n6785 ) ;
  assign n6788 = ( n6653 & n6786 ) | ( n6653 & ~n6787 ) | ( n6786 & ~n6787 ) ;
  assign n6789 = ( n6712 & n6781 ) | ( n6712 & n6788 ) | ( n6781 & n6788 ) ;
  assign n6790 = ( ~n6712 & n6781 ) | ( ~n6712 & n6788 ) | ( n6781 & n6788 ) ;
  assign n6791 = ( n6712 & ~n6789 ) | ( n6712 & n6790 ) | ( ~n6789 & n6790 ) ;
  assign n6792 = ( ~n6707 & n6735 ) | ( ~n6707 & n6791 ) | ( n6735 & n6791 ) ;
  assign n6793 = ( n6707 & n6735 ) | ( n6707 & n6791 ) | ( n6735 & n6791 ) ;
  assign n6794 = ( n6707 & n6792 ) | ( n6707 & ~n6793 ) | ( n6792 & ~n6793 ) ;
  assign n6795 = ( n6716 & n6718 ) | ( n6716 & n6794 ) | ( n6718 & n6794 ) ;
  assign n6796 = ( n6716 & ~n6718 ) | ( n6716 & n6794 ) | ( ~n6718 & n6794 ) ;
  assign n6797 = ( n6718 & ~n6795 ) | ( n6718 & n6796 ) | ( ~n6795 & n6796 ) ;
  assign n6798 = ( n6745 & n6749 ) | ( n6745 & n6765 ) | ( n6749 & n6765 ) ;
  assign n6799 = ( n6745 & n6749 ) | ( n6745 & ~n6765 ) | ( n6749 & ~n6765 ) ;
  assign n6800 = ( n6765 & ~n6798 ) | ( n6765 & n6799 ) | ( ~n6798 & n6799 ) ;
  assign n6801 = ( n6752 & n6774 ) | ( n6752 & n6800 ) | ( n6774 & n6800 ) ;
  assign n6802 = ( ~n6752 & n6774 ) | ( ~n6752 & n6800 ) | ( n6774 & n6800 ) ;
  assign n6803 = ( n6752 & ~n6801 ) | ( n6752 & n6802 ) | ( ~n6801 & n6802 ) ;
  assign n6804 = ( n6779 & ~n6787 ) | ( n6779 & n6803 ) | ( ~n6787 & n6803 ) ;
  assign n6805 = ( n6779 & n6787 ) | ( n6779 & n6803 ) | ( n6787 & n6803 ) ;
  assign n6806 = ( n6787 & n6804 ) | ( n6787 & ~n6805 ) | ( n6804 & ~n6805 ) ;
  assign n6807 = ( ~n6725 & n6759 ) | ( ~n6725 & n6771 ) | ( n6759 & n6771 ) ;
  assign n6808 = ( n6725 & n6759 ) | ( n6725 & n6771 ) | ( n6759 & n6771 ) ;
  assign n6809 = ( n6725 & n6807 ) | ( n6725 & ~n6808 ) | ( n6807 & ~n6808 ) ;
  assign n6810 = x37 & x53 ;
  assign n6811 = x38 & x52 ;
  assign n6812 = x36 & x54 ;
  assign n6813 = ( ~n6810 & n6811 ) | ( ~n6810 & n6812 ) | ( n6811 & n6812 ) ;
  assign n6814 = ( n6810 & n6811 ) | ( n6810 & n6812 ) | ( n6811 & n6812 ) ;
  assign n6815 = ( n6810 & n6813 ) | ( n6810 & ~n6814 ) | ( n6813 & ~n6814 ) ;
  assign n6816 = x34 & x56 ;
  assign n6817 = x33 & x57 ;
  assign n6818 = x35 & x55 ;
  assign n6819 = ( ~n6816 & n6817 ) | ( ~n6816 & n6818 ) | ( n6817 & n6818 ) ;
  assign n6820 = ( n6816 & n6817 ) | ( n6816 & n6818 ) | ( n6817 & n6818 ) ;
  assign n6821 = ( n6816 & n6819 ) | ( n6816 & ~n6820 ) | ( n6819 & ~n6820 ) ;
  assign n6822 = x42 & x48 ;
  assign n6823 = x44 & x46 ;
  assign n6824 = x43 & x47 ;
  assign n6825 = ( ~n6822 & n6823 ) | ( ~n6822 & n6824 ) | ( n6823 & n6824 ) ;
  assign n6826 = ( n6822 & n6823 ) | ( n6822 & n6824 ) | ( n6823 & n6824 ) ;
  assign n6827 = ( n6822 & n6825 ) | ( n6822 & ~n6826 ) | ( n6825 & ~n6826 ) ;
  assign n6828 = ( ~n6815 & n6821 ) | ( ~n6815 & n6827 ) | ( n6821 & n6827 ) ;
  assign n6829 = ( n6815 & n6821 ) | ( n6815 & n6827 ) | ( n6821 & n6827 ) ;
  assign n6830 = ( n6815 & n6828 ) | ( n6815 & ~n6829 ) | ( n6828 & ~n6829 ) ;
  assign n6831 = ( n6783 & n6809 ) | ( n6783 & n6830 ) | ( n6809 & n6830 ) ;
  assign n6832 = ( ~n6783 & n6809 ) | ( ~n6783 & n6830 ) | ( n6809 & n6830 ) ;
  assign n6833 = ( n6783 & ~n6831 ) | ( n6783 & n6832 ) | ( ~n6831 & n6832 ) ;
  assign n6834 = x27 & x63 ;
  assign n6835 = x28 & x62 ;
  assign n6836 = x29 & x61 ;
  assign n6837 = ( ~n6834 & n6835 ) | ( ~n6834 & n6836 ) | ( n6835 & n6836 ) ;
  assign n6838 = ( n6834 & n6835 ) | ( n6834 & n6836 ) | ( n6835 & n6836 ) ;
  assign n6839 = ( n6834 & n6837 ) | ( n6834 & ~n6838 ) | ( n6837 & ~n6838 ) ;
  assign n6840 = x30 & x60 ;
  assign n6841 = x32 & x58 ;
  assign n6842 = ( ~n3736 & n6840 ) | ( ~n3736 & n6841 ) | ( n6840 & n6841 ) ;
  assign n6843 = ( n3736 & n6840 ) | ( n3736 & n6841 ) | ( n6840 & n6841 ) ;
  assign n6844 = ( n3736 & n6842 ) | ( n3736 & ~n6843 ) | ( n6842 & ~n6843 ) ;
  assign n6845 = ( ~n6738 & n6839 ) | ( ~n6738 & n6844 ) | ( n6839 & n6844 ) ;
  assign n6846 = ( n6738 & n6839 ) | ( n6738 & n6844 ) | ( n6839 & n6844 ) ;
  assign n6847 = ( n6738 & n6845 ) | ( n6738 & ~n6846 ) | ( n6845 & ~n6846 ) ;
  assign n6848 = x41 & x49 ;
  assign n6849 = x40 & x50 ;
  assign n6850 = x39 & x51 ;
  assign n6851 = ( ~n6848 & n6849 ) | ( ~n6848 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6852 = ( n6848 & n6849 ) | ( n6848 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6853 = ( n6848 & n6851 ) | ( n6848 & ~n6852 ) | ( n6851 & ~n6852 ) ;
  assign n6854 = ( n6728 & n6777 ) | ( n6728 & n6853 ) | ( n6777 & n6853 ) ;
  assign n6855 = ( ~n6728 & n6777 ) | ( ~n6728 & n6853 ) | ( n6777 & n6853 ) ;
  assign n6856 = ( n6728 & ~n6854 ) | ( n6728 & n6855 ) | ( ~n6854 & n6855 ) ;
  assign n6857 = ( n6730 & n6847 ) | ( n6730 & n6856 ) | ( n6847 & n6856 ) ;
  assign n6858 = ( ~n6730 & n6847 ) | ( ~n6730 & n6856 ) | ( n6847 & n6856 ) ;
  assign n6859 = ( n6730 & ~n6857 ) | ( n6730 & n6858 ) | ( ~n6857 & n6858 ) ;
  assign n6860 = ( n6733 & n6833 ) | ( n6733 & n6859 ) | ( n6833 & n6859 ) ;
  assign n6861 = ( ~n6733 & n6833 ) | ( ~n6733 & n6859 ) | ( n6833 & n6859 ) ;
  assign n6862 = ( n6733 & ~n6860 ) | ( n6733 & n6861 ) | ( ~n6860 & n6861 ) ;
  assign n6863 = ( n6789 & ~n6806 ) | ( n6789 & n6862 ) | ( ~n6806 & n6862 ) ;
  assign n6864 = ( n6789 & n6806 ) | ( n6789 & n6862 ) | ( n6806 & n6862 ) ;
  assign n6865 = ( n6806 & n6863 ) | ( n6806 & ~n6864 ) | ( n6863 & ~n6864 ) ;
  assign n6866 = ( n6793 & n6795 ) | ( n6793 & n6865 ) | ( n6795 & n6865 ) ;
  assign n6867 = ( n6793 & ~n6795 ) | ( n6793 & n6865 ) | ( ~n6795 & n6865 ) ;
  assign n6868 = ( n6795 & ~n6866 ) | ( n6795 & n6867 ) | ( ~n6866 & n6867 ) ;
  assign n6869 = x34 & x57 ;
  assign n6870 = x42 & x49 ;
  assign n6871 = x36 & x55 ;
  assign n6872 = ( ~n6869 & n6870 ) | ( ~n6869 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = ( n6869 & n6870 ) | ( n6869 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6874 = ( n6869 & n6872 ) | ( n6869 & ~n6873 ) | ( n6872 & ~n6873 ) ;
  assign n6875 = ( n6798 & ~n6808 ) | ( n6798 & n6874 ) | ( ~n6808 & n6874 ) ;
  assign n6876 = ( n6798 & n6808 ) | ( n6798 & n6874 ) | ( n6808 & n6874 ) ;
  assign n6877 = ( n6808 & n6875 ) | ( n6808 & ~n6876 ) | ( n6875 & ~n6876 ) ;
  assign n6878 = x32 & x59 ;
  assign n6879 = x33 & x58 ;
  assign n6880 = x31 & x60 ;
  assign n6881 = ( ~n6878 & n6879 ) | ( ~n6878 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6882 = ( n6878 & n6879 ) | ( n6878 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6883 = ( n6878 & n6881 ) | ( n6878 & ~n6882 ) | ( n6881 & ~n6882 ) ;
  assign n6884 = x39 & x52 ;
  assign n6885 = x38 & x53 ;
  assign n6886 = x37 & x54 ;
  assign n6887 = ( ~n6884 & n6885 ) | ( ~n6884 & n6886 ) | ( n6885 & n6886 ) ;
  assign n6888 = ( n6884 & n6885 ) | ( n6884 & n6886 ) | ( n6885 & n6886 ) ;
  assign n6889 = ( n6884 & n6887 ) | ( n6884 & ~n6888 ) | ( n6887 & ~n6888 ) ;
  assign n6890 = ( ~n6852 & n6883 ) | ( ~n6852 & n6889 ) | ( n6883 & n6889 ) ;
  assign n6891 = ( n6852 & n6883 ) | ( n6852 & n6889 ) | ( n6883 & n6889 ) ;
  assign n6892 = ( n6852 & n6890 ) | ( n6852 & ~n6891 ) | ( n6890 & ~n6891 ) ;
  assign n6893 = ( n6801 & n6877 ) | ( n6801 & n6892 ) | ( n6877 & n6892 ) ;
  assign n6894 = ( ~n6801 & n6877 ) | ( ~n6801 & n6892 ) | ( n6877 & n6892 ) ;
  assign n6895 = ( n6801 & ~n6893 ) | ( n6801 & n6894 ) | ( ~n6893 & n6894 ) ;
  assign n6896 = ( ~n6814 & n6838 ) | ( ~n6814 & n6843 ) | ( n6838 & n6843 ) ;
  assign n6897 = ( n6814 & n6838 ) | ( n6814 & n6843 ) | ( n6838 & n6843 ) ;
  assign n6898 = ( n6814 & n6896 ) | ( n6814 & ~n6897 ) | ( n6896 & ~n6897 ) ;
  assign n6899 = x43 & x48 ;
  assign n6900 = x44 & x47 ;
  assign n6901 = x35 & x56 ;
  assign n6902 = ( ~n6899 & n6900 ) | ( ~n6899 & n6901 ) | ( n6900 & n6901 ) ;
  assign n6903 = ( n6899 & n6900 ) | ( n6899 & n6901 ) | ( n6900 & n6901 ) ;
  assign n6904 = ( n6899 & n6902 ) | ( n6899 & ~n6903 ) | ( n6902 & ~n6903 ) ;
  assign n6905 = x40 & x51 ;
  assign n6906 = x41 & x50 ;
  assign n6907 = x28 & x63 ;
  assign n6908 = ( ~n6905 & n6906 ) | ( ~n6905 & n6907 ) | ( n6906 & n6907 ) ;
  assign n6909 = ( n6905 & n6906 ) | ( n6905 & n6907 ) | ( n6906 & n6907 ) ;
  assign n6910 = ( n6905 & n6908 ) | ( n6905 & ~n6909 ) | ( n6908 & ~n6909 ) ;
  assign n6911 = x29 & x62 ;
  assign n6912 = x45 & x46 ;
  assign n6913 = ( x46 & n6911 ) | ( x46 & n6912 ) | ( n6911 & n6912 ) ;
  assign n6914 = ( x46 & ~n6911 ) | ( x46 & n6912 ) | ( ~n6911 & n6912 ) ;
  assign n6915 = ( n6911 & ~n6913 ) | ( n6911 & n6914 ) | ( ~n6913 & n6914 ) ;
  assign n6916 = ( ~n6904 & n6910 ) | ( ~n6904 & n6915 ) | ( n6910 & n6915 ) ;
  assign n6917 = ( n6904 & n6910 ) | ( n6904 & n6915 ) | ( n6910 & n6915 ) ;
  assign n6918 = ( n6904 & n6916 ) | ( n6904 & ~n6917 ) | ( n6916 & ~n6917 ) ;
  assign n6919 = ( n6854 & n6898 ) | ( n6854 & n6918 ) | ( n6898 & n6918 ) ;
  assign n6920 = ( ~n6854 & n6898 ) | ( ~n6854 & n6918 ) | ( n6898 & n6918 ) ;
  assign n6921 = ( n6854 & ~n6919 ) | ( n6854 & n6920 ) | ( ~n6919 & n6920 ) ;
  assign n6922 = ( n6805 & ~n6895 ) | ( n6805 & n6921 ) | ( ~n6895 & n6921 ) ;
  assign n6923 = ( n6805 & n6895 ) | ( n6805 & n6921 ) | ( n6895 & n6921 ) ;
  assign n6924 = ( n6895 & n6922 ) | ( n6895 & ~n6923 ) | ( n6922 & ~n6923 ) ;
  assign n6925 = ( n4131 & n6820 ) | ( n4131 & n6826 ) | ( n6820 & n6826 ) ;
  assign n6926 = ( ~n4131 & n6820 ) | ( ~n4131 & n6826 ) | ( n6820 & n6826 ) ;
  assign n6927 = ( n4131 & ~n6925 ) | ( n4131 & n6926 ) | ( ~n6925 & n6926 ) ;
  assign n6928 = ( n6829 & n6846 ) | ( n6829 & ~n6927 ) | ( n6846 & ~n6927 ) ;
  assign n6929 = ( n6829 & n6846 ) | ( n6829 & n6927 ) | ( n6846 & n6927 ) ;
  assign n6930 = ( n6927 & n6928 ) | ( n6927 & ~n6929 ) | ( n6928 & ~n6929 ) ;
  assign n6931 = ( n6831 & n6857 ) | ( n6831 & n6930 ) | ( n6857 & n6930 ) ;
  assign n6932 = ( n6831 & ~n6857 ) | ( n6831 & n6930 ) | ( ~n6857 & n6930 ) ;
  assign n6933 = ( n6857 & ~n6931 ) | ( n6857 & n6932 ) | ( ~n6931 & n6932 ) ;
  assign n6934 = ( ~n6860 & n6924 ) | ( ~n6860 & n6933 ) | ( n6924 & n6933 ) ;
  assign n6935 = ( n6860 & n6924 ) | ( n6860 & n6933 ) | ( n6924 & n6933 ) ;
  assign n6936 = ( n6860 & n6934 ) | ( n6860 & ~n6935 ) | ( n6934 & ~n6935 ) ;
  assign n6937 = ( n6864 & ~n6866 ) | ( n6864 & n6936 ) | ( ~n6866 & n6936 ) ;
  assign n6938 = ( n6864 & n6866 ) | ( n6864 & n6936 ) | ( n6866 & n6936 ) ;
  assign n6939 = ( n6866 & n6937 ) | ( n6866 & ~n6938 ) | ( n6937 & ~n6938 ) ;
  assign n6940 = x31 & x61 ;
  assign n6941 = x30 & x62 ;
  assign n6942 = ( ~n6913 & n6940 ) | ( ~n6913 & n6941 ) | ( n6940 & n6941 ) ;
  assign n6943 = ( n6913 & n6940 ) | ( n6913 & n6941 ) | ( n6940 & n6941 ) ;
  assign n6944 = ( n6913 & n6942 ) | ( n6913 & ~n6943 ) | ( n6942 & ~n6943 ) ;
  assign n6945 = x41 & x51 ;
  assign n6946 = x40 & x52 ;
  assign n6947 = x39 & x53 ;
  assign n6948 = ( ~n6945 & n6946 ) | ( ~n6945 & n6947 ) | ( n6946 & n6947 ) ;
  assign n6949 = ( n6945 & n6946 ) | ( n6945 & n6947 ) | ( n6946 & n6947 ) ;
  assign n6950 = ( n6945 & n6948 ) | ( n6945 & ~n6949 ) | ( n6948 & ~n6949 ) ;
  assign n6951 = ( ~n6925 & n6944 ) | ( ~n6925 & n6950 ) | ( n6944 & n6950 ) ;
  assign n6952 = ( n6925 & n6944 ) | ( n6925 & n6950 ) | ( n6944 & n6950 ) ;
  assign n6953 = ( n6925 & n6951 ) | ( n6925 & ~n6952 ) | ( n6951 & ~n6952 ) ;
  assign n6954 = x42 & x50 ;
  assign n6955 = x35 & x57 ;
  assign n6956 = x34 & x58 ;
  assign n6957 = ( ~n6954 & n6955 ) | ( ~n6954 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6958 = ( n6954 & n6955 ) | ( n6954 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6959 = ( n6954 & n6957 ) | ( n6954 & ~n6958 ) | ( n6957 & ~n6958 ) ;
  assign n6960 = x36 & x56 ;
  assign n6961 = x33 & x59 ;
  assign n6962 = x29 & x63 ;
  assign n6963 = ( ~n6960 & n6961 ) | ( ~n6960 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = ( n6960 & n6961 ) | ( n6960 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6965 = ( n6960 & n6963 ) | ( n6960 & ~n6964 ) | ( n6963 & ~n6964 ) ;
  assign n6966 = x45 & x47 ;
  assign n6967 = x44 & x48 ;
  assign n6968 = x43 & x49 ;
  assign n6969 = ( ~n6966 & n6967 ) | ( ~n6966 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = ( n6966 & n6967 ) | ( n6966 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6971 = ( n6966 & n6969 ) | ( n6966 & ~n6970 ) | ( n6969 & ~n6970 ) ;
  assign n6972 = ( ~n6959 & n6965 ) | ( ~n6959 & n6971 ) | ( n6965 & n6971 ) ;
  assign n6973 = ( n6959 & n6965 ) | ( n6959 & n6971 ) | ( n6965 & n6971 ) ;
  assign n6974 = ( n6959 & n6972 ) | ( n6959 & ~n6973 ) | ( n6972 & ~n6973 ) ;
  assign n6975 = ( n6929 & n6953 ) | ( n6929 & n6974 ) | ( n6953 & n6974 ) ;
  assign n6976 = ( ~n6929 & n6953 ) | ( ~n6929 & n6974 ) | ( n6953 & n6974 ) ;
  assign n6977 = ( n6929 & ~n6975 ) | ( n6929 & n6976 ) | ( ~n6975 & n6976 ) ;
  assign n6978 = ( n6893 & n6931 ) | ( n6893 & n6977 ) | ( n6931 & n6977 ) ;
  assign n6979 = ( n6893 & ~n6931 ) | ( n6893 & n6977 ) | ( ~n6931 & n6977 ) ;
  assign n6980 = ( n6931 & ~n6978 ) | ( n6931 & n6979 ) | ( ~n6978 & n6979 ) ;
  assign n6981 = ( n6891 & ~n6897 ) | ( n6891 & n6917 ) | ( ~n6897 & n6917 ) ;
  assign n6982 = ( n6891 & n6897 ) | ( n6891 & n6917 ) | ( n6897 & n6917 ) ;
  assign n6983 = ( n6897 & n6981 ) | ( n6897 & ~n6982 ) | ( n6981 & ~n6982 ) ;
  assign n6984 = ( n6882 & ~n6888 ) | ( n6882 & n6909 ) | ( ~n6888 & n6909 ) ;
  assign n6985 = ( n6882 & n6888 ) | ( n6882 & n6909 ) | ( n6888 & n6909 ) ;
  assign n6986 = ( n6888 & n6984 ) | ( n6888 & ~n6985 ) | ( n6984 & ~n6985 ) ;
  assign n6987 = x32 & x60 ;
  assign n6988 = x38 & x54 ;
  assign n6989 = x37 & x55 ;
  assign n6990 = ( ~n6987 & n6988 ) | ( ~n6987 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6991 = ( n6987 & n6988 ) | ( n6987 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6992 = ( n6987 & n6990 ) | ( n6987 & ~n6991 ) | ( n6990 & ~n6991 ) ;
  assign n6993 = ( n6873 & n6903 ) | ( n6873 & ~n6992 ) | ( n6903 & ~n6992 ) ;
  assign n6994 = ( n6873 & n6903 ) | ( n6873 & n6992 ) | ( n6903 & n6992 ) ;
  assign n6995 = ( n6992 & n6993 ) | ( n6992 & ~n6994 ) | ( n6993 & ~n6994 ) ;
  assign n6996 = ( n6876 & n6986 ) | ( n6876 & n6995 ) | ( n6986 & n6995 ) ;
  assign n6997 = ( ~n6876 & n6986 ) | ( ~n6876 & n6995 ) | ( n6986 & n6995 ) ;
  assign n6998 = ( n6876 & ~n6996 ) | ( n6876 & n6997 ) | ( ~n6996 & n6997 ) ;
  assign n6999 = ( n6919 & n6983 ) | ( n6919 & n6998 ) | ( n6983 & n6998 ) ;
  assign n7000 = ( n6919 & ~n6983 ) | ( n6919 & n6998 ) | ( ~n6983 & n6998 ) ;
  assign n7001 = ( n6983 & ~n6999 ) | ( n6983 & n7000 ) | ( ~n6999 & n7000 ) ;
  assign n7002 = ( n6923 & n6980 ) | ( n6923 & n7001 ) | ( n6980 & n7001 ) ;
  assign n7003 = ( n6923 & ~n6980 ) | ( n6923 & n7001 ) | ( ~n6980 & n7001 ) ;
  assign n7004 = ( n6980 & ~n7002 ) | ( n6980 & n7003 ) | ( ~n7002 & n7003 ) ;
  assign n7005 = ( n6935 & n6938 ) | ( n6935 & n7004 ) | ( n6938 & n7004 ) ;
  assign n7006 = ( n6935 & ~n6938 ) | ( n6935 & n7004 ) | ( ~n6938 & n7004 ) ;
  assign n7007 = ( n6938 & ~n7005 ) | ( n6938 & n7006 ) | ( ~n7005 & n7006 ) ;
  assign n7008 = x44 & x49 ;
  assign n7009 = x42 & x51 ;
  assign n7010 = x43 & x50 ;
  assign n7011 = ( ~n7008 & n7009 ) | ( ~n7008 & n7010 ) | ( n7009 & n7010 ) ;
  assign n7012 = ( n7008 & n7009 ) | ( n7008 & n7010 ) | ( n7009 & n7010 ) ;
  assign n7013 = ( n7008 & n7011 ) | ( n7008 & ~n7012 ) | ( n7011 & ~n7012 ) ;
  assign n7014 = x45 & x48 ;
  assign n7015 = x38 & x55 ;
  assign n7016 = x37 & x56 ;
  assign n7017 = ( ~n7014 & n7015 ) | ( ~n7014 & n7016 ) | ( n7015 & n7016 ) ;
  assign n7018 = ( n7014 & n7015 ) | ( n7014 & n7016 ) | ( n7015 & n7016 ) ;
  assign n7019 = ( n7014 & n7017 ) | ( n7014 & ~n7018 ) | ( n7017 & ~n7018 ) ;
  assign n7020 = x31 & x62 ;
  assign n7021 = x46 & x47 ;
  assign n7022 = ( x47 & n7020 ) | ( x47 & n7021 ) | ( n7020 & n7021 ) ;
  assign n7023 = ( x47 & ~n7020 ) | ( x47 & n7021 ) | ( ~n7020 & n7021 ) ;
  assign n7024 = ( n7020 & ~n7022 ) | ( n7020 & n7023 ) | ( ~n7022 & n7023 ) ;
  assign n7025 = ( ~n7013 & n7019 ) | ( ~n7013 & n7024 ) | ( n7019 & n7024 ) ;
  assign n7026 = ( n7013 & n7019 ) | ( n7013 & n7024 ) | ( n7019 & n7024 ) ;
  assign n7027 = ( n7013 & n7025 ) | ( n7013 & ~n7026 ) | ( n7025 & ~n7026 ) ;
  assign n7028 = x32 & x61 ;
  assign n7029 = x30 & x63 ;
  assign n7030 = x33 & x60 ;
  assign n7031 = ( ~n7028 & n7029 ) | ( ~n7028 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7032 = ( n7028 & n7029 ) | ( n7028 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7033 = ( n7028 & n7031 ) | ( n7028 & ~n7032 ) | ( n7031 & ~n7032 ) ;
  assign n7034 = x41 & x52 ;
  assign n7035 = x40 & x53 ;
  assign n7036 = x34 & x59 ;
  assign n7037 = ( ~n7034 & n7035 ) | ( ~n7034 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7038 = ( n7034 & n7035 ) | ( n7034 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7039 = ( n7034 & n7037 ) | ( n7034 & ~n7038 ) | ( n7037 & ~n7038 ) ;
  assign n7040 = x35 & x58 ;
  assign n7041 = x36 & x57 ;
  assign n7042 = x39 & x54 ;
  assign n7043 = ( ~n7040 & n7041 ) | ( ~n7040 & n7042 ) | ( n7041 & n7042 ) ;
  assign n7044 = ( n7040 & n7041 ) | ( n7040 & n7042 ) | ( n7041 & n7042 ) ;
  assign n7045 = ( n7040 & n7043 ) | ( n7040 & ~n7044 ) | ( n7043 & ~n7044 ) ;
  assign n7046 = ( ~n7033 & n7039 ) | ( ~n7033 & n7045 ) | ( n7039 & n7045 ) ;
  assign n7047 = ( n7033 & n7039 ) | ( n7033 & n7045 ) | ( n7039 & n7045 ) ;
  assign n7048 = ( n7033 & n7046 ) | ( n7033 & ~n7047 ) | ( n7046 & ~n7047 ) ;
  assign n7049 = ( n6982 & n7027 ) | ( n6982 & n7048 ) | ( n7027 & n7048 ) ;
  assign n7050 = ( ~n6982 & n7027 ) | ( ~n6982 & n7048 ) | ( n7027 & n7048 ) ;
  assign n7051 = ( n6982 & ~n7049 ) | ( n6982 & n7050 ) | ( ~n7049 & n7050 ) ;
  assign n7052 = ( n6975 & n6999 ) | ( n6975 & n7051 ) | ( n6999 & n7051 ) ;
  assign n7053 = ( n6975 & ~n6999 ) | ( n6975 & n7051 ) | ( ~n6999 & n7051 ) ;
  assign n7054 = ( n6999 & ~n7052 ) | ( n6999 & n7053 ) | ( ~n7052 & n7053 ) ;
  assign n7055 = ( ~n6943 & n6964 ) | ( ~n6943 & n6991 ) | ( n6964 & n6991 ) ;
  assign n7056 = ( n6943 & n6964 ) | ( n6943 & n6991 ) | ( n6964 & n6991 ) ;
  assign n7057 = ( n6943 & n7055 ) | ( n6943 & ~n7056 ) | ( n7055 & ~n7056 ) ;
  assign n7058 = ( n6949 & ~n6958 ) | ( n6949 & n6970 ) | ( ~n6958 & n6970 ) ;
  assign n7059 = ( n6949 & n6958 ) | ( n6949 & n6970 ) | ( n6958 & n6970 ) ;
  assign n7060 = ( n6958 & n7058 ) | ( n6958 & ~n7059 ) | ( n7058 & ~n7059 ) ;
  assign n7061 = ( n6952 & n7057 ) | ( n6952 & n7060 ) | ( n7057 & n7060 ) ;
  assign n7062 = ( ~n6952 & n7057 ) | ( ~n6952 & n7060 ) | ( n7057 & n7060 ) ;
  assign n7063 = ( n6952 & ~n7061 ) | ( n6952 & n7062 ) | ( ~n7061 & n7062 ) ;
  assign n7064 = ( ~n6973 & n6985 ) | ( ~n6973 & n6994 ) | ( n6985 & n6994 ) ;
  assign n7065 = ( n6973 & n6985 ) | ( n6973 & n6994 ) | ( n6985 & n6994 ) ;
  assign n7066 = ( n6973 & n7064 ) | ( n6973 & ~n7065 ) | ( n7064 & ~n7065 ) ;
  assign n7067 = ( n6996 & n7063 ) | ( n6996 & n7066 ) | ( n7063 & n7066 ) ;
  assign n7068 = ( n6996 & ~n7063 ) | ( n6996 & n7066 ) | ( ~n7063 & n7066 ) ;
  assign n7069 = ( n7063 & ~n7067 ) | ( n7063 & n7068 ) | ( ~n7067 & n7068 ) ;
  assign n7070 = ( n6978 & n7054 ) | ( n6978 & n7069 ) | ( n7054 & n7069 ) ;
  assign n7071 = ( ~n6978 & n7054 ) | ( ~n6978 & n7069 ) | ( n7054 & n7069 ) ;
  assign n7072 = ( n6978 & ~n7070 ) | ( n6978 & n7071 ) | ( ~n7070 & n7071 ) ;
  assign n7073 = ( n7002 & n7005 ) | ( n7002 & n7072 ) | ( n7005 & n7072 ) ;
  assign n7074 = ( n7002 & ~n7005 ) | ( n7002 & n7072 ) | ( ~n7005 & n7072 ) ;
  assign n7075 = ( n7005 & ~n7073 ) | ( n7005 & n7074 ) | ( ~n7073 & n7074 ) ;
  assign n7076 = x33 & x61 ;
  assign n7077 = x35 & x59 ;
  assign n7078 = ( ~n4197 & n7076 ) | ( ~n4197 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7079 = ( n4197 & n7076 ) | ( n4197 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7080 = ( n4197 & n7078 ) | ( n4197 & ~n7079 ) | ( n7078 & ~n7079 ) ;
  assign n7081 = x37 & x57 ;
  assign n7082 = x39 & x55 ;
  assign n7083 = x34 & x60 ;
  assign n7084 = ( ~n7081 & n7082 ) | ( ~n7081 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7085 = ( n7081 & n7082 ) | ( n7081 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7086 = ( n7081 & n7084 ) | ( n7081 & ~n7085 ) | ( n7084 & ~n7085 ) ;
  assign n7087 = ( ~n7012 & n7080 ) | ( ~n7012 & n7086 ) | ( n7080 & n7086 ) ;
  assign n7088 = ( n7012 & n7080 ) | ( n7012 & n7086 ) | ( n7080 & n7086 ) ;
  assign n7089 = ( n7012 & n7087 ) | ( n7012 & ~n7088 ) | ( n7087 & ~n7088 ) ;
  assign n7090 = x43 & x51 ;
  assign n7091 = x36 & x58 ;
  assign n7092 = x44 & x50 ;
  assign n7093 = ( ~n7090 & n7091 ) | ( ~n7090 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7094 = ( n7090 & n7091 ) | ( n7090 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7095 = ( n7090 & n7093 ) | ( n7090 & ~n7094 ) | ( n7093 & ~n7094 ) ;
  assign n7096 = x41 & x53 ;
  assign n7097 = x42 & x52 ;
  assign n7098 = x40 & x54 ;
  assign n7099 = ( ~n7096 & n7097 ) | ( ~n7096 & n7098 ) | ( n7097 & n7098 ) ;
  assign n7100 = ( n7096 & n7097 ) | ( n7096 & n7098 ) | ( n7097 & n7098 ) ;
  assign n7101 = ( n7096 & n7099 ) | ( n7096 & ~n7100 ) | ( n7099 & ~n7100 ) ;
  assign n7102 = x38 & x56 ;
  assign n7103 = x46 & x48 ;
  assign n7104 = x45 & x49 ;
  assign n7105 = ( ~n7102 & n7103 ) | ( ~n7102 & n7104 ) | ( n7103 & n7104 ) ;
  assign n7106 = ( n7102 & n7103 ) | ( n7102 & n7104 ) | ( n7103 & n7104 ) ;
  assign n7107 = ( n7102 & n7105 ) | ( n7102 & ~n7106 ) | ( n7105 & ~n7106 ) ;
  assign n7108 = ( ~n7095 & n7101 ) | ( ~n7095 & n7107 ) | ( n7101 & n7107 ) ;
  assign n7109 = ( n7095 & n7101 ) | ( n7095 & n7107 ) | ( n7101 & n7107 ) ;
  assign n7110 = ( n7095 & n7108 ) | ( n7095 & ~n7109 ) | ( n7108 & ~n7109 ) ;
  assign n7111 = ( ~n7065 & n7089 ) | ( ~n7065 & n7110 ) | ( n7089 & n7110 ) ;
  assign n7112 = ( n7065 & n7089 ) | ( n7065 & n7110 ) | ( n7089 & n7110 ) ;
  assign n7113 = ( n7065 & n7111 ) | ( n7065 & ~n7112 ) | ( n7111 & ~n7112 ) ;
  assign n7114 = x31 & x63 ;
  assign n7115 = ( n7018 & n7022 ) | ( n7018 & n7114 ) | ( n7022 & n7114 ) ;
  assign n7116 = ( ~n7018 & n7022 ) | ( ~n7018 & n7114 ) | ( n7022 & n7114 ) ;
  assign n7117 = ( n7018 & ~n7115 ) | ( n7018 & n7116 ) | ( ~n7115 & n7116 ) ;
  assign n7118 = ( ~n7032 & n7038 ) | ( ~n7032 & n7044 ) | ( n7038 & n7044 ) ;
  assign n7119 = ( n7032 & n7038 ) | ( n7032 & n7044 ) | ( n7038 & n7044 ) ;
  assign n7120 = ( n7032 & n7118 ) | ( n7032 & ~n7119 ) | ( n7118 & ~n7119 ) ;
  assign n7121 = ( n7026 & n7117 ) | ( n7026 & n7120 ) | ( n7117 & n7120 ) ;
  assign n7122 = ( ~n7026 & n7117 ) | ( ~n7026 & n7120 ) | ( n7117 & n7120 ) ;
  assign n7123 = ( n7026 & ~n7121 ) | ( n7026 & n7122 ) | ( ~n7121 & n7122 ) ;
  assign n7124 = ( ~n7067 & n7113 ) | ( ~n7067 & n7123 ) | ( n7113 & n7123 ) ;
  assign n7125 = ( n7067 & n7113 ) | ( n7067 & n7123 ) | ( n7113 & n7123 ) ;
  assign n7126 = ( n7067 & n7124 ) | ( n7067 & ~n7125 ) | ( n7124 & ~n7125 ) ;
  assign n7127 = ( n7047 & ~n7056 ) | ( n7047 & n7059 ) | ( ~n7056 & n7059 ) ;
  assign n7128 = ( n7047 & n7056 ) | ( n7047 & n7059 ) | ( n7056 & n7059 ) ;
  assign n7129 = ( n7056 & n7127 ) | ( n7056 & ~n7128 ) | ( n7127 & ~n7128 ) ;
  assign n7130 = ( n7049 & n7061 ) | ( n7049 & n7129 ) | ( n7061 & n7129 ) ;
  assign n7131 = ( ~n7049 & n7061 ) | ( ~n7049 & n7129 ) | ( n7061 & n7129 ) ;
  assign n7132 = ( n7049 & ~n7130 ) | ( n7049 & n7131 ) | ( ~n7130 & n7131 ) ;
  assign n7133 = ( n7052 & n7126 ) | ( n7052 & n7132 ) | ( n7126 & n7132 ) ;
  assign n7134 = ( n7052 & ~n7126 ) | ( n7052 & n7132 ) | ( ~n7126 & n7132 ) ;
  assign n7135 = ( n7126 & ~n7133 ) | ( n7126 & n7134 ) | ( ~n7133 & n7134 ) ;
  assign n7136 = ( n7070 & n7073 ) | ( n7070 & n7135 ) | ( n7073 & n7135 ) ;
  assign n7137 = ( n7070 & ~n7073 ) | ( n7070 & n7135 ) | ( ~n7073 & n7135 ) ;
  assign n7138 = ( n7073 & ~n7136 ) | ( n7073 & n7137 ) | ( ~n7136 & n7137 ) ;
  assign n7139 = x40 & x55 ;
  assign n7140 = x38 & x57 ;
  assign n7141 = x37 & x58 ;
  assign n7142 = ( ~n7139 & n7140 ) | ( ~n7139 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7143 = ( n7139 & n7140 ) | ( n7139 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7144 = ( n7139 & n7142 ) | ( n7139 & ~n7143 ) | ( n7142 & ~n7143 ) ;
  assign n7145 = x41 & x54 ;
  assign n7146 = x34 & x61 ;
  assign n7147 = ( ~n4325 & n7145 ) | ( ~n4325 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7148 = ( n4325 & n7145 ) | ( n4325 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7149 = ( n4325 & n7147 ) | ( n4325 & ~n7148 ) | ( n7147 & ~n7148 ) ;
  assign n7150 = ( ~n7094 & n7144 ) | ( ~n7094 & n7149 ) | ( n7144 & n7149 ) ;
  assign n7151 = ( n7094 & n7144 ) | ( n7094 & n7149 ) | ( n7144 & n7149 ) ;
  assign n7152 = ( n7094 & n7150 ) | ( n7094 & ~n7151 ) | ( n7150 & ~n7151 ) ;
  assign n7153 = x46 & x49 ;
  assign n7154 = x39 & x56 ;
  assign n7155 = x45 & x50 ;
  assign n7156 = ( ~n7153 & n7154 ) | ( ~n7153 & n7155 ) | ( n7154 & n7155 ) ;
  assign n7157 = ( n7153 & n7154 ) | ( n7153 & n7155 ) | ( n7154 & n7155 ) ;
  assign n7158 = ( n7153 & n7156 ) | ( n7153 & ~n7157 ) | ( n7156 & ~n7157 ) ;
  assign n7159 = x42 & x53 ;
  assign n7160 = x43 & x52 ;
  assign n7161 = x44 & x51 ;
  assign n7162 = ( ~n7159 & n7160 ) | ( ~n7159 & n7161 ) | ( n7160 & n7161 ) ;
  assign n7163 = ( n7159 & n7160 ) | ( n7159 & n7161 ) | ( n7160 & n7161 ) ;
  assign n7164 = ( n7159 & n7162 ) | ( n7159 & ~n7163 ) | ( n7162 & ~n7163 ) ;
  assign n7165 = x33 & x62 ;
  assign n7166 = x47 & x48 ;
  assign n7167 = ( x48 & n7165 ) | ( x48 & n7166 ) | ( n7165 & n7166 ) ;
  assign n7168 = ( x48 & ~n7165 ) | ( x48 & n7166 ) | ( ~n7165 & n7166 ) ;
  assign n7169 = ( n7165 & ~n7167 ) | ( n7165 & n7168 ) | ( ~n7167 & n7168 ) ;
  assign n7170 = ( ~n7158 & n7164 ) | ( ~n7158 & n7169 ) | ( n7164 & n7169 ) ;
  assign n7171 = ( n7158 & n7164 ) | ( n7158 & n7169 ) | ( n7164 & n7169 ) ;
  assign n7172 = ( n7158 & n7170 ) | ( n7158 & ~n7171 ) | ( n7170 & ~n7171 ) ;
  assign n7173 = ( n7128 & n7152 ) | ( n7128 & n7172 ) | ( n7152 & n7172 ) ;
  assign n7174 = ( ~n7128 & n7152 ) | ( ~n7128 & n7172 ) | ( n7152 & n7172 ) ;
  assign n7175 = ( n7128 & ~n7173 ) | ( n7128 & n7174 ) | ( ~n7173 & n7174 ) ;
  assign n7176 = ( ~n7079 & n7085 ) | ( ~n7079 & n7100 ) | ( n7085 & n7100 ) ;
  assign n7177 = ( n7079 & n7085 ) | ( n7079 & n7100 ) | ( n7085 & n7100 ) ;
  assign n7178 = ( n7079 & n7176 ) | ( n7079 & ~n7177 ) | ( n7176 & ~n7177 ) ;
  assign n7179 = ( n7088 & n7109 ) | ( n7088 & n7178 ) | ( n7109 & n7178 ) ;
  assign n7180 = ( ~n7088 & n7109 ) | ( ~n7088 & n7178 ) | ( n7109 & n7178 ) ;
  assign n7181 = ( n7088 & ~n7179 ) | ( n7088 & n7180 ) | ( ~n7179 & n7180 ) ;
  assign n7182 = ( n7130 & n7175 ) | ( n7130 & n7181 ) | ( n7175 & n7181 ) ;
  assign n7183 = ( ~n7130 & n7175 ) | ( ~n7130 & n7181 ) | ( n7175 & n7181 ) ;
  assign n7184 = ( n7130 & ~n7182 ) | ( n7130 & n7183 ) | ( ~n7182 & n7183 ) ;
  assign n7185 = x36 & x59 ;
  assign n7186 = x35 & x60 ;
  assign n7187 = ( n7106 & n7185 ) | ( n7106 & n7186 ) | ( n7185 & n7186 ) ;
  assign n7188 = ( ~n7106 & n7185 ) | ( ~n7106 & n7186 ) | ( n7185 & n7186 ) ;
  assign n7189 = ( n7106 & ~n7187 ) | ( n7106 & n7188 ) | ( ~n7187 & n7188 ) ;
  assign n7190 = ( n7115 & n7119 ) | ( n7115 & n7189 ) | ( n7119 & n7189 ) ;
  assign n7191 = ( n7115 & n7119 ) | ( n7115 & ~n7189 ) | ( n7119 & ~n7189 ) ;
  assign n7192 = ( n7189 & ~n7190 ) | ( n7189 & n7191 ) | ( ~n7190 & n7191 ) ;
  assign n7193 = ( ~n7112 & n7121 ) | ( ~n7112 & n7192 ) | ( n7121 & n7192 ) ;
  assign n7194 = ( n7112 & n7121 ) | ( n7112 & n7192 ) | ( n7121 & n7192 ) ;
  assign n7195 = ( n7112 & n7193 ) | ( n7112 & ~n7194 ) | ( n7193 & ~n7194 ) ;
  assign n7196 = ( n7125 & n7184 ) | ( n7125 & n7195 ) | ( n7184 & n7195 ) ;
  assign n7197 = ( n7125 & ~n7184 ) | ( n7125 & n7195 ) | ( ~n7184 & n7195 ) ;
  assign n7198 = ( n7184 & ~n7196 ) | ( n7184 & n7197 ) | ( ~n7196 & n7197 ) ;
  assign n7199 = ( n7133 & ~n7136 ) | ( n7133 & n7198 ) | ( ~n7136 & n7198 ) ;
  assign n7200 = ( n7133 & n7136 ) | ( n7133 & n7198 ) | ( n7136 & n7198 ) ;
  assign n7201 = ( n7136 & n7199 ) | ( n7136 & ~n7200 ) | ( n7199 & ~n7200 ) ;
  assign n7202 = ( n7143 & n7148 ) | ( n7143 & ~n7187 ) | ( n7148 & ~n7187 ) ;
  assign n7203 = ( n7143 & n7148 ) | ( n7143 & n7187 ) | ( n7148 & n7187 ) ;
  assign n7204 = ( n7187 & n7202 ) | ( n7187 & ~n7203 ) | ( n7202 & ~n7203 ) ;
  assign n7205 = x41 & x55 ;
  assign n7206 = x43 & x53 ;
  assign n7207 = x42 & x54 ;
  assign n7208 = ( ~n7205 & n7206 ) | ( ~n7205 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( n7205 & n7206 ) | ( n7205 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7210 = ( n7205 & n7208 ) | ( n7205 & ~n7209 ) | ( n7208 & ~n7209 ) ;
  assign n7211 = x33 & x63 ;
  assign n7212 = x34 & x62 ;
  assign n7213 = x35 & x61 ;
  assign n7214 = ( ~n7211 & n7212 ) | ( ~n7211 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7215 = ( n7211 & n7212 ) | ( n7211 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7216 = ( n7211 & n7214 ) | ( n7211 & ~n7215 ) | ( n7214 & ~n7215 ) ;
  assign n7217 = ( ~n7177 & n7210 ) | ( ~n7177 & n7216 ) | ( n7210 & n7216 ) ;
  assign n7218 = ( n7177 & n7210 ) | ( n7177 & n7216 ) | ( n7210 & n7216 ) ;
  assign n7219 = ( n7177 & n7217 ) | ( n7177 & ~n7218 ) | ( n7217 & ~n7218 ) ;
  assign n7220 = ( n7190 & n7204 ) | ( n7190 & n7219 ) | ( n7204 & n7219 ) ;
  assign n7221 = ( ~n7190 & n7204 ) | ( ~n7190 & n7219 ) | ( n7204 & n7219 ) ;
  assign n7222 = ( n7190 & ~n7220 ) | ( n7190 & n7221 ) | ( ~n7220 & n7221 ) ;
  assign n7223 = ( n7157 & n7163 ) | ( n7157 & n7167 ) | ( n7163 & n7167 ) ;
  assign n7224 = ( ~n7157 & n7163 ) | ( ~n7157 & n7167 ) | ( n7163 & n7167 ) ;
  assign n7225 = ( n7157 & ~n7223 ) | ( n7157 & n7224 ) | ( ~n7223 & n7224 ) ;
  assign n7226 = ( n7151 & n7171 ) | ( n7151 & n7225 ) | ( n7171 & n7225 ) ;
  assign n7227 = ( ~n7151 & n7171 ) | ( ~n7151 & n7225 ) | ( n7171 & n7225 ) ;
  assign n7228 = ( n7151 & ~n7226 ) | ( n7151 & n7227 ) | ( ~n7226 & n7227 ) ;
  assign n7229 = ( n7194 & ~n7222 ) | ( n7194 & n7228 ) | ( ~n7222 & n7228 ) ;
  assign n7230 = ( n7194 & n7222 ) | ( n7194 & n7228 ) | ( n7222 & n7228 ) ;
  assign n7231 = ( n7222 & n7229 ) | ( n7222 & ~n7230 ) | ( n7229 & ~n7230 ) ;
  assign n7232 = x47 & x49 ;
  assign n7233 = x46 & x50 ;
  assign n7234 = x45 & x51 ;
  assign n7235 = ( ~n7232 & n7233 ) | ( ~n7232 & n7234 ) | ( n7233 & n7234 ) ;
  assign n7236 = ( n7232 & n7233 ) | ( n7232 & n7234 ) | ( n7233 & n7234 ) ;
  assign n7237 = ( n7232 & n7235 ) | ( n7232 & ~n7236 ) | ( n7235 & ~n7236 ) ;
  assign n7238 = x39 & x57 ;
  assign n7239 = x44 & x52 ;
  assign n7240 = x38 & x58 ;
  assign n7241 = ( ~n7238 & n7239 ) | ( ~n7238 & n7240 ) | ( n7239 & n7240 ) ;
  assign n7242 = ( n7238 & n7239 ) | ( n7238 & n7240 ) | ( n7239 & n7240 ) ;
  assign n7243 = ( n7238 & n7241 ) | ( n7238 & ~n7242 ) | ( n7241 & ~n7242 ) ;
  assign n7244 = x40 & x56 ;
  assign n7245 = x36 & x60 ;
  assign n7246 = x37 & x59 ;
  assign n7247 = ( ~n7244 & n7245 ) | ( ~n7244 & n7246 ) | ( n7245 & n7246 ) ;
  assign n7248 = ( n7244 & n7245 ) | ( n7244 & n7246 ) | ( n7245 & n7246 ) ;
  assign n7249 = ( n7244 & n7247 ) | ( n7244 & ~n7248 ) | ( n7247 & ~n7248 ) ;
  assign n7250 = ( ~n7237 & n7243 ) | ( ~n7237 & n7249 ) | ( n7243 & n7249 ) ;
  assign n7251 = ( n7237 & n7243 ) | ( n7237 & n7249 ) | ( n7243 & n7249 ) ;
  assign n7252 = ( n7237 & n7250 ) | ( n7237 & ~n7251 ) | ( n7250 & ~n7251 ) ;
  assign n7253 = ( n7173 & n7179 ) | ( n7173 & ~n7252 ) | ( n7179 & ~n7252 ) ;
  assign n7254 = ( n7173 & n7179 ) | ( n7173 & n7252 ) | ( n7179 & n7252 ) ;
  assign n7255 = ( n7252 & n7253 ) | ( n7252 & ~n7254 ) | ( n7253 & ~n7254 ) ;
  assign n7256 = ( ~n7182 & n7231 ) | ( ~n7182 & n7255 ) | ( n7231 & n7255 ) ;
  assign n7257 = ( n7182 & n7231 ) | ( n7182 & n7255 ) | ( n7231 & n7255 ) ;
  assign n7258 = ( n7182 & n7256 ) | ( n7182 & ~n7257 ) | ( n7256 & ~n7257 ) ;
  assign n7259 = ( n7196 & ~n7200 ) | ( n7196 & n7258 ) | ( ~n7200 & n7258 ) ;
  assign n7260 = ( n7196 & n7200 ) | ( n7196 & n7258 ) | ( n7200 & n7258 ) ;
  assign n7261 = ( n7200 & n7259 ) | ( n7200 & ~n7260 ) | ( n7259 & ~n7260 ) ;
  assign n7262 = x36 & x61 ;
  assign n7263 = ( n7236 & n7242 ) | ( n7236 & n7262 ) | ( n7242 & n7262 ) ;
  assign n7264 = ( ~n7236 & n7242 ) | ( ~n7236 & n7262 ) | ( n7242 & n7262 ) ;
  assign n7265 = ( n7236 & ~n7263 ) | ( n7236 & n7264 ) | ( ~n7263 & n7264 ) ;
  assign n7266 = ( n7203 & n7251 ) | ( n7203 & n7265 ) | ( n7251 & n7265 ) ;
  assign n7267 = ( ~n7203 & n7251 ) | ( ~n7203 & n7265 ) | ( n7251 & n7265 ) ;
  assign n7268 = ( n7203 & ~n7266 ) | ( n7203 & n7267 ) | ( ~n7266 & n7267 ) ;
  assign n7269 = x46 & x51 ;
  assign n7270 = x40 & x57 ;
  assign n7271 = x47 & x50 ;
  assign n7272 = ( ~n7269 & n7270 ) | ( ~n7269 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7273 = ( n7269 & n7270 ) | ( n7269 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7274 = ( n7269 & n7272 ) | ( n7269 & ~n7273 ) | ( n7272 & ~n7273 ) ;
  assign n7275 = x35 & x62 ;
  assign n7276 = x48 & x49 ;
  assign n7277 = ( x49 & n7275 ) | ( x49 & n7276 ) | ( n7275 & n7276 ) ;
  assign n7278 = ( x49 & ~n7275 ) | ( x49 & n7276 ) | ( ~n7275 & n7276 ) ;
  assign n7279 = ( n7275 & ~n7277 ) | ( n7275 & n7278 ) | ( ~n7277 & n7278 ) ;
  assign n7280 = ( ~n7223 & n7274 ) | ( ~n7223 & n7279 ) | ( n7274 & n7279 ) ;
  assign n7281 = ( n7223 & n7274 ) | ( n7223 & n7279 ) | ( n7274 & n7279 ) ;
  assign n7282 = ( n7223 & n7280 ) | ( n7223 & ~n7281 ) | ( n7280 & ~n7281 ) ;
  assign n7283 = ( n7209 & n7215 ) | ( n7209 & ~n7248 ) | ( n7215 & ~n7248 ) ;
  assign n7284 = ( n7209 & n7215 ) | ( n7209 & n7248 ) | ( n7215 & n7248 ) ;
  assign n7285 = ( n7248 & n7283 ) | ( n7248 & ~n7284 ) | ( n7283 & ~n7284 ) ;
  assign n7286 = ( n7218 & n7282 ) | ( n7218 & n7285 ) | ( n7282 & n7285 ) ;
  assign n7287 = ( n7218 & ~n7282 ) | ( n7218 & n7285 ) | ( ~n7282 & n7285 ) ;
  assign n7288 = ( n7282 & ~n7286 ) | ( n7282 & n7287 ) | ( ~n7286 & n7287 ) ;
  assign n7289 = ( n7254 & n7268 ) | ( n7254 & n7288 ) | ( n7268 & n7288 ) ;
  assign n7290 = ( ~n7254 & n7268 ) | ( ~n7254 & n7288 ) | ( n7268 & n7288 ) ;
  assign n7291 = ( n7254 & ~n7289 ) | ( n7254 & n7290 ) | ( ~n7289 & n7290 ) ;
  assign n7292 = x45 & x52 ;
  assign n7293 = x43 & x54 ;
  assign n7294 = x44 & x53 ;
  assign n7295 = ( ~n7292 & n7293 ) | ( ~n7292 & n7294 ) | ( n7293 & n7294 ) ;
  assign n7296 = ( n7292 & n7293 ) | ( n7292 & n7294 ) | ( n7293 & n7294 ) ;
  assign n7297 = ( n7292 & n7295 ) | ( n7292 & ~n7296 ) | ( n7295 & ~n7296 ) ;
  assign n7298 = x38 & x59 ;
  assign n7299 = x39 & x58 ;
  assign n7300 = x37 & x60 ;
  assign n7301 = ( ~n7298 & n7299 ) | ( ~n7298 & n7300 ) | ( n7299 & n7300 ) ;
  assign n7302 = ( n7298 & n7299 ) | ( n7298 & n7300 ) | ( n7299 & n7300 ) ;
  assign n7303 = ( n7298 & n7301 ) | ( n7298 & ~n7302 ) | ( n7301 & ~n7302 ) ;
  assign n7304 = x34 & x63 ;
  assign n7305 = x42 & x55 ;
  assign n7306 = x41 & x56 ;
  assign n7307 = ( ~n7304 & n7305 ) | ( ~n7304 & n7306 ) | ( n7305 & n7306 ) ;
  assign n7308 = ( n7304 & n7305 ) | ( n7304 & n7306 ) | ( n7305 & n7306 ) ;
  assign n7309 = ( n7304 & n7307 ) | ( n7304 & ~n7308 ) | ( n7307 & ~n7308 ) ;
  assign n7310 = ( ~n7297 & n7303 ) | ( ~n7297 & n7309 ) | ( n7303 & n7309 ) ;
  assign n7311 = ( n7297 & n7303 ) | ( n7297 & n7309 ) | ( n7303 & n7309 ) ;
  assign n7312 = ( n7297 & n7310 ) | ( n7297 & ~n7311 ) | ( n7310 & ~n7311 ) ;
  assign n7313 = ( n7220 & n7226 ) | ( n7220 & n7312 ) | ( n7226 & n7312 ) ;
  assign n7314 = ( ~n7220 & n7226 ) | ( ~n7220 & n7312 ) | ( n7226 & n7312 ) ;
  assign n7315 = ( n7220 & ~n7313 ) | ( n7220 & n7314 ) | ( ~n7313 & n7314 ) ;
  assign n7316 = ( ~n7230 & n7291 ) | ( ~n7230 & n7315 ) | ( n7291 & n7315 ) ;
  assign n7317 = ( n7230 & n7291 ) | ( n7230 & n7315 ) | ( n7291 & n7315 ) ;
  assign n7318 = ( n7230 & n7316 ) | ( n7230 & ~n7317 ) | ( n7316 & ~n7317 ) ;
  assign n7319 = ( n7257 & ~n7260 ) | ( n7257 & n7318 ) | ( ~n7260 & n7318 ) ;
  assign n7320 = ( n7257 & n7260 ) | ( n7257 & n7318 ) | ( n7260 & n7318 ) ;
  assign n7321 = ( n7260 & n7319 ) | ( n7260 & ~n7320 ) | ( n7319 & ~n7320 ) ;
  assign n7322 = ( n7263 & n7284 ) | ( n7263 & ~n7311 ) | ( n7284 & ~n7311 ) ;
  assign n7323 = ( n7263 & n7284 ) | ( n7263 & n7311 ) | ( n7284 & n7311 ) ;
  assign n7324 = ( n7311 & n7322 ) | ( n7311 & ~n7323 ) | ( n7322 & ~n7323 ) ;
  assign n7325 = x36 & x62 ;
  assign n7326 = x37 & x61 ;
  assign n7327 = ( ~n7277 & n7325 ) | ( ~n7277 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7328 = ( n7277 & n7325 ) | ( n7277 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7329 = ( n7277 & n7327 ) | ( n7277 & ~n7328 ) | ( n7327 & ~n7328 ) ;
  assign n7330 = x40 & x58 ;
  assign n7331 = x39 & x59 ;
  assign n7332 = x45 & x53 ;
  assign n7333 = ( ~n7330 & n7331 ) | ( ~n7330 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7334 = ( n7330 & n7331 ) | ( n7330 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7335 = ( n7330 & n7333 ) | ( n7330 & ~n7334 ) | ( n7333 & ~n7334 ) ;
  assign n7336 = x48 & x50 ;
  assign n7337 = x46 & x52 ;
  assign n7338 = x47 & x51 ;
  assign n7339 = ( ~n7336 & n7337 ) | ( ~n7336 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7340 = ( n7336 & n7337 ) | ( n7336 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7341 = ( n7336 & n7339 ) | ( n7336 & ~n7340 ) | ( n7339 & ~n7340 ) ;
  assign n7342 = ( ~n7329 & n7335 ) | ( ~n7329 & n7341 ) | ( n7335 & n7341 ) ;
  assign n7343 = ( n7329 & n7335 ) | ( n7329 & n7341 ) | ( n7335 & n7341 ) ;
  assign n7344 = ( n7329 & n7342 ) | ( n7329 & ~n7343 ) | ( n7342 & ~n7343 ) ;
  assign n7345 = ( ~n7296 & n7302 ) | ( ~n7296 & n7308 ) | ( n7302 & n7308 ) ;
  assign n7346 = ( n7296 & n7302 ) | ( n7296 & n7308 ) | ( n7302 & n7308 ) ;
  assign n7347 = ( n7296 & n7345 ) | ( n7296 & ~n7346 ) | ( n7345 & ~n7346 ) ;
  assign n7348 = ( n7281 & n7344 ) | ( n7281 & n7347 ) | ( n7344 & n7347 ) ;
  assign n7349 = ( n7281 & ~n7344 ) | ( n7281 & n7347 ) | ( ~n7344 & n7347 ) ;
  assign n7350 = ( n7344 & ~n7348 ) | ( n7344 & n7349 ) | ( ~n7348 & n7349 ) ;
  assign n7351 = ( n7313 & n7324 ) | ( n7313 & n7350 ) | ( n7324 & n7350 ) ;
  assign n7352 = ( ~n7313 & n7324 ) | ( ~n7313 & n7350 ) | ( n7324 & n7350 ) ;
  assign n7353 = ( n7313 & ~n7351 ) | ( n7313 & n7352 ) | ( ~n7351 & n7352 ) ;
  assign n7354 = x42 & x56 ;
  assign n7355 = x38 & x60 ;
  assign n7356 = x41 & x57 ;
  assign n7357 = ( ~n7354 & n7355 ) | ( ~n7354 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7358 = ( n7354 & n7355 ) | ( n7354 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7359 = ( n7354 & n7357 ) | ( n7354 & ~n7358 ) | ( n7357 & ~n7358 ) ;
  assign n7360 = x44 & x54 ;
  assign n7361 = x43 & x55 ;
  assign n7362 = x35 & x63 ;
  assign n7363 = ( ~n7360 & n7361 ) | ( ~n7360 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7364 = ( n7360 & n7361 ) | ( n7360 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7365 = ( n7360 & n7363 ) | ( n7360 & ~n7364 ) | ( n7363 & ~n7364 ) ;
  assign n7366 = ( ~n7273 & n7359 ) | ( ~n7273 & n7365 ) | ( n7359 & n7365 ) ;
  assign n7367 = ( n7273 & n7359 ) | ( n7273 & n7365 ) | ( n7359 & n7365 ) ;
  assign n7368 = ( n7273 & n7366 ) | ( n7273 & ~n7367 ) | ( n7366 & ~n7367 ) ;
  assign n7369 = ( n7266 & n7286 ) | ( n7266 & n7368 ) | ( n7286 & n7368 ) ;
  assign n7370 = ( n7266 & ~n7286 ) | ( n7266 & n7368 ) | ( ~n7286 & n7368 ) ;
  assign n7371 = ( n7286 & ~n7369 ) | ( n7286 & n7370 ) | ( ~n7369 & n7370 ) ;
  assign n7372 = ( n7289 & n7353 ) | ( n7289 & n7371 ) | ( n7353 & n7371 ) ;
  assign n7373 = ( n7289 & ~n7353 ) | ( n7289 & n7371 ) | ( ~n7353 & n7371 ) ;
  assign n7374 = ( n7353 & ~n7372 ) | ( n7353 & n7373 ) | ( ~n7372 & n7373 ) ;
  assign n7375 = ( n7317 & ~n7320 ) | ( n7317 & n7374 ) | ( ~n7320 & n7374 ) ;
  assign n7376 = ( n7317 & n7320 ) | ( n7317 & n7374 ) | ( n7320 & n7374 ) ;
  assign n7377 = ( n7320 & n7375 ) | ( n7320 & ~n7376 ) | ( n7375 & ~n7376 ) ;
  assign n7378 = x40 & x59 ;
  assign n7379 = x44 & x55 ;
  assign n7380 = x41 & x58 ;
  assign n7381 = ( ~n7378 & n7379 ) | ( ~n7378 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7382 = ( n7378 & n7379 ) | ( n7378 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7383 = ( n7378 & n7381 ) | ( n7378 & ~n7382 ) | ( n7381 & ~n7382 ) ;
  assign n7384 = x47 & x52 ;
  assign n7385 = x45 & x54 ;
  assign n7386 = x46 & x53 ;
  assign n7387 = ( ~n7384 & n7385 ) | ( ~n7384 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7388 = ( n7384 & n7385 ) | ( n7384 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7389 = ( n7384 & n7387 ) | ( n7384 & ~n7388 ) | ( n7387 & ~n7388 ) ;
  assign n7390 = x43 & x56 ;
  assign n7391 = x48 & x51 ;
  assign n7392 = x42 & x57 ;
  assign n7393 = ( ~n7390 & n7391 ) | ( ~n7390 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7394 = ( n7390 & n7391 ) | ( n7390 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7395 = ( n7390 & n7393 ) | ( n7390 & ~n7394 ) | ( n7393 & ~n7394 ) ;
  assign n7396 = ( ~n7383 & n7389 ) | ( ~n7383 & n7395 ) | ( n7389 & n7395 ) ;
  assign n7397 = ( n7383 & n7389 ) | ( n7383 & n7395 ) | ( n7389 & n7395 ) ;
  assign n7398 = ( n7383 & n7396 ) | ( n7383 & ~n7397 ) | ( n7396 & ~n7397 ) ;
  assign n7399 = ( n7323 & n7348 ) | ( n7323 & n7398 ) | ( n7348 & n7398 ) ;
  assign n7400 = ( n7323 & ~n7348 ) | ( n7323 & n7398 ) | ( ~n7348 & n7398 ) ;
  assign n7401 = ( n7348 & ~n7399 ) | ( n7348 & n7400 ) | ( ~n7399 & n7400 ) ;
  assign n7402 = x37 & x62 ;
  assign n7403 = x49 & x50 ;
  assign n7404 = ( x50 & n7402 ) | ( x50 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7405 = ( x50 & ~n7402 ) | ( x50 & n7403 ) | ( ~n7402 & n7403 ) ;
  assign n7406 = ( n7402 & ~n7404 ) | ( n7402 & n7405 ) | ( ~n7404 & n7405 ) ;
  assign n7407 = ( n7346 & ~n7367 ) | ( n7346 & n7406 ) | ( ~n7367 & n7406 ) ;
  assign n7408 = ( n7346 & n7367 ) | ( n7346 & n7406 ) | ( n7367 & n7406 ) ;
  assign n7409 = ( n7367 & n7407 ) | ( n7367 & ~n7408 ) | ( n7407 & ~n7408 ) ;
  assign n7410 = x39 & x60 ;
  assign n7411 = x36 & x63 ;
  assign n7412 = x38 & x61 ;
  assign n7413 = ( ~n7410 & n7411 ) | ( ~n7410 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = ( n7410 & n7411 ) | ( n7410 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7415 = ( n7410 & n7413 ) | ( n7410 & ~n7414 ) | ( n7413 & ~n7414 ) ;
  assign n7416 = ( ~n7328 & n7358 ) | ( ~n7328 & n7415 ) | ( n7358 & n7415 ) ;
  assign n7417 = ( n7328 & n7358 ) | ( n7328 & n7415 ) | ( n7358 & n7415 ) ;
  assign n7418 = ( n7328 & n7416 ) | ( n7328 & ~n7417 ) | ( n7416 & ~n7417 ) ;
  assign n7419 = ( ~n7334 & n7340 ) | ( ~n7334 & n7364 ) | ( n7340 & n7364 ) ;
  assign n7420 = ( n7334 & n7340 ) | ( n7334 & n7364 ) | ( n7340 & n7364 ) ;
  assign n7421 = ( n7334 & n7419 ) | ( n7334 & ~n7420 ) | ( n7419 & ~n7420 ) ;
  assign n7422 = ( n7343 & ~n7418 ) | ( n7343 & n7421 ) | ( ~n7418 & n7421 ) ;
  assign n7423 = ( n7343 & n7418 ) | ( n7343 & n7421 ) | ( n7418 & n7421 ) ;
  assign n7424 = ( n7418 & n7422 ) | ( n7418 & ~n7423 ) | ( n7422 & ~n7423 ) ;
  assign n7425 = ( n7369 & n7409 ) | ( n7369 & n7424 ) | ( n7409 & n7424 ) ;
  assign n7426 = ( ~n7369 & n7409 ) | ( ~n7369 & n7424 ) | ( n7409 & n7424 ) ;
  assign n7427 = ( n7369 & ~n7425 ) | ( n7369 & n7426 ) | ( ~n7425 & n7426 ) ;
  assign n7428 = ( ~n7351 & n7401 ) | ( ~n7351 & n7427 ) | ( n7401 & n7427 ) ;
  assign n7429 = ( n7351 & n7401 ) | ( n7351 & n7427 ) | ( n7401 & n7427 ) ;
  assign n7430 = ( n7351 & n7428 ) | ( n7351 & ~n7429 ) | ( n7428 & ~n7429 ) ;
  assign n7431 = ( n7372 & ~n7376 ) | ( n7372 & n7430 ) | ( ~n7376 & n7430 ) ;
  assign n7432 = ( n7372 & n7376 ) | ( n7372 & n7430 ) | ( n7376 & n7430 ) ;
  assign n7433 = ( n7376 & n7431 ) | ( n7376 & ~n7432 ) | ( n7431 & ~n7432 ) ;
  assign n7434 = x48 & x52 ;
  assign n7435 = x47 & x53 ;
  assign n7436 = x49 & x51 ;
  assign n7437 = ( ~n7434 & n7435 ) | ( ~n7434 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7438 = ( n7434 & n7435 ) | ( n7434 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7439 = ( n7434 & n7437 ) | ( n7434 & ~n7438 ) | ( n7437 & ~n7438 ) ;
  assign n7440 = ( ~n7417 & n7420 ) | ( ~n7417 & n7439 ) | ( n7420 & n7439 ) ;
  assign n7441 = ( n7417 & n7420 ) | ( n7417 & n7439 ) | ( n7420 & n7439 ) ;
  assign n7442 = ( n7417 & n7440 ) | ( n7417 & ~n7441 ) | ( n7440 & ~n7441 ) ;
  assign n7443 = ( n7382 & n7388 ) | ( n7382 & ~n7414 ) | ( n7388 & ~n7414 ) ;
  assign n7444 = ( n7382 & n7388 ) | ( n7382 & n7414 ) | ( n7388 & n7414 ) ;
  assign n7445 = ( n7414 & n7443 ) | ( n7414 & ~n7444 ) | ( n7443 & ~n7444 ) ;
  assign n7446 = x37 & x63 ;
  assign n7447 = ( n7394 & n7404 ) | ( n7394 & n7446 ) | ( n7404 & n7446 ) ;
  assign n7448 = ( ~n7394 & n7404 ) | ( ~n7394 & n7446 ) | ( n7404 & n7446 ) ;
  assign n7449 = ( n7394 & ~n7447 ) | ( n7394 & n7448 ) | ( ~n7447 & n7448 ) ;
  assign n7450 = ( n7397 & n7445 ) | ( n7397 & n7449 ) | ( n7445 & n7449 ) ;
  assign n7451 = ( ~n7397 & n7445 ) | ( ~n7397 & n7449 ) | ( n7445 & n7449 ) ;
  assign n7452 = ( n7397 & ~n7450 ) | ( n7397 & n7451 ) | ( ~n7450 & n7451 ) ;
  assign n7453 = ( ~n7399 & n7442 ) | ( ~n7399 & n7452 ) | ( n7442 & n7452 ) ;
  assign n7454 = ( n7399 & n7442 ) | ( n7399 & n7452 ) | ( n7442 & n7452 ) ;
  assign n7455 = ( n7399 & n7453 ) | ( n7399 & ~n7454 ) | ( n7453 & ~n7454 ) ;
  assign n7456 = x43 & x57 ;
  assign n7457 = x44 & x56 ;
  assign n7458 = x45 & x55 ;
  assign n7459 = ( ~n7456 & n7457 ) | ( ~n7456 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7460 = ( n7456 & n7457 ) | ( n7456 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7461 = ( n7456 & n7459 ) | ( n7456 & ~n7460 ) | ( n7459 & ~n7460 ) ;
  assign n7462 = x46 & x54 ;
  assign n7463 = x42 & x58 ;
  assign n7464 = x41 & x59 ;
  assign n7465 = ( ~n7462 & n7463 ) | ( ~n7462 & n7464 ) | ( n7463 & n7464 ) ;
  assign n7466 = ( n7462 & n7463 ) | ( n7462 & n7464 ) | ( n7463 & n7464 ) ;
  assign n7467 = ( n7462 & n7465 ) | ( n7462 & ~n7466 ) | ( n7465 & ~n7466 ) ;
  assign n7468 = x40 & x60 ;
  assign n7469 = x38 & x62 ;
  assign n7470 = x39 & x61 ;
  assign n7471 = ( ~n7468 & n7469 ) | ( ~n7468 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7472 = ( n7468 & n7469 ) | ( n7468 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7473 = ( n7468 & n7471 ) | ( n7468 & ~n7472 ) | ( n7471 & ~n7472 ) ;
  assign n7474 = ( ~n7461 & n7467 ) | ( ~n7461 & n7473 ) | ( n7467 & n7473 ) ;
  assign n7475 = ( n7461 & n7467 ) | ( n7461 & n7473 ) | ( n7467 & n7473 ) ;
  assign n7476 = ( n7461 & n7474 ) | ( n7461 & ~n7475 ) | ( n7474 & ~n7475 ) ;
  assign n7477 = ( n7408 & n7423 ) | ( n7408 & n7476 ) | ( n7423 & n7476 ) ;
  assign n7478 = ( n7408 & ~n7423 ) | ( n7408 & n7476 ) | ( ~n7423 & n7476 ) ;
  assign n7479 = ( n7423 & ~n7477 ) | ( n7423 & n7478 ) | ( ~n7477 & n7478 ) ;
  assign n7480 = ( n7425 & n7455 ) | ( n7425 & n7479 ) | ( n7455 & n7479 ) ;
  assign n7481 = ( n7425 & ~n7455 ) | ( n7425 & n7479 ) | ( ~n7455 & n7479 ) ;
  assign n7482 = ( n7455 & ~n7480 ) | ( n7455 & n7481 ) | ( ~n7480 & n7481 ) ;
  assign n7483 = ( n7429 & ~n7432 ) | ( n7429 & n7482 ) | ( ~n7432 & n7482 ) ;
  assign n7484 = ( n7429 & n7432 ) | ( n7429 & n7482 ) | ( n7432 & n7482 ) ;
  assign n7485 = ( n7432 & n7483 ) | ( n7432 & ~n7484 ) | ( n7483 & ~n7484 ) ;
  assign n7486 = ( ~n7460 & n7466 ) | ( ~n7460 & n7472 ) | ( n7466 & n7472 ) ;
  assign n7487 = ( n7460 & n7466 ) | ( n7460 & n7472 ) | ( n7466 & n7472 ) ;
  assign n7488 = ( n7460 & n7486 ) | ( n7460 & ~n7487 ) | ( n7486 & ~n7487 ) ;
  assign n7489 = ( n7444 & n7475 ) | ( n7444 & n7488 ) | ( n7475 & n7488 ) ;
  assign n7490 = ( n7444 & n7475 ) | ( n7444 & ~n7488 ) | ( n7475 & ~n7488 ) ;
  assign n7491 = ( n7488 & ~n7489 ) | ( n7488 & n7490 ) | ( ~n7489 & n7490 ) ;
  assign n7492 = ( n7450 & ~n7477 ) | ( n7450 & n7491 ) | ( ~n7477 & n7491 ) ;
  assign n7493 = ( n7450 & n7477 ) | ( n7450 & n7491 ) | ( n7477 & n7491 ) ;
  assign n7494 = ( n7477 & n7492 ) | ( n7477 & ~n7493 ) | ( n7492 & ~n7493 ) ;
  assign n7495 = x40 & x61 ;
  assign n7496 = x41 & x60 ;
  assign n7497 = ( n7438 & n7495 ) | ( n7438 & n7496 ) | ( n7495 & n7496 ) ;
  assign n7498 = ( ~n7438 & n7495 ) | ( ~n7438 & n7496 ) | ( n7495 & n7496 ) ;
  assign n7499 = ( n7438 & ~n7497 ) | ( n7438 & n7498 ) | ( ~n7497 & n7498 ) ;
  assign n7500 = x39 & x62 ;
  assign n7501 = x50 & x51 ;
  assign n7502 = ( x51 & n7500 ) | ( x51 & n7501 ) | ( n7500 & n7501 ) ;
  assign n7503 = ( x51 & ~n7500 ) | ( x51 & n7501 ) | ( ~n7500 & n7501 ) ;
  assign n7504 = ( n7500 & ~n7502 ) | ( n7500 & n7503 ) | ( ~n7502 & n7503 ) ;
  assign n7505 = ( n7447 & n7499 ) | ( n7447 & n7504 ) | ( n7499 & n7504 ) ;
  assign n7506 = ( n7447 & ~n7499 ) | ( n7447 & n7504 ) | ( ~n7499 & n7504 ) ;
  assign n7507 = ( n7499 & ~n7505 ) | ( n7499 & n7506 ) | ( ~n7505 & n7506 ) ;
  assign n7508 = x48 & x53 ;
  assign n7509 = x44 & x57 ;
  assign n7510 = x49 & x52 ;
  assign n7511 = ( ~n7508 & n7509 ) | ( ~n7508 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = ( n7508 & n7509 ) | ( n7508 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7513 = ( n7508 & n7511 ) | ( n7508 & ~n7512 ) | ( n7511 & ~n7512 ) ;
  assign n7514 = x45 & x56 ;
  assign n7515 = x42 & x59 ;
  assign n7516 = x43 & x58 ;
  assign n7517 = ( ~n7514 & n7515 ) | ( ~n7514 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = ( n7514 & n7515 ) | ( n7514 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7519 = ( n7514 & n7517 ) | ( n7514 & ~n7518 ) | ( n7517 & ~n7518 ) ;
  assign n7520 = x47 & x54 ;
  assign n7521 = x38 & x63 ;
  assign n7522 = x46 & x55 ;
  assign n7523 = ( ~n7520 & n7521 ) | ( ~n7520 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = ( n7520 & n7521 ) | ( n7520 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7525 = ( n7520 & n7523 ) | ( n7520 & ~n7524 ) | ( n7523 & ~n7524 ) ;
  assign n7526 = ( ~n7513 & n7519 ) | ( ~n7513 & n7525 ) | ( n7519 & n7525 ) ;
  assign n7527 = ( n7513 & n7519 ) | ( n7513 & n7525 ) | ( n7519 & n7525 ) ;
  assign n7528 = ( n7513 & n7526 ) | ( n7513 & ~n7527 ) | ( n7526 & ~n7527 ) ;
  assign n7529 = ( n7441 & n7507 ) | ( n7441 & n7528 ) | ( n7507 & n7528 ) ;
  assign n7530 = ( ~n7441 & n7507 ) | ( ~n7441 & n7528 ) | ( n7507 & n7528 ) ;
  assign n7531 = ( n7441 & ~n7529 ) | ( n7441 & n7530 ) | ( ~n7529 & n7530 ) ;
  assign n7532 = ( n7454 & n7494 ) | ( n7454 & n7531 ) | ( n7494 & n7531 ) ;
  assign n7533 = ( ~n7454 & n7494 ) | ( ~n7454 & n7531 ) | ( n7494 & n7531 ) ;
  assign n7534 = ( n7454 & ~n7532 ) | ( n7454 & n7533 ) | ( ~n7532 & n7533 ) ;
  assign n7535 = ( n7480 & ~n7484 ) | ( n7480 & n7534 ) | ( ~n7484 & n7534 ) ;
  assign n7536 = ( n7480 & n7484 ) | ( n7480 & n7534 ) | ( n7484 & n7534 ) ;
  assign n7537 = ( n7484 & n7535 ) | ( n7484 & ~n7536 ) | ( n7535 & ~n7536 ) ;
  assign n7538 = ( n7502 & n7512 ) | ( n7502 & n7524 ) | ( n7512 & n7524 ) ;
  assign n7539 = ( n7502 & n7512 ) | ( n7502 & ~n7524 ) | ( n7512 & ~n7524 ) ;
  assign n7540 = ( n7524 & ~n7538 ) | ( n7524 & n7539 ) | ( ~n7538 & n7539 ) ;
  assign n7541 = ( n7487 & n7527 ) | ( n7487 & n7540 ) | ( n7527 & n7540 ) ;
  assign n7542 = ( n7487 & n7527 ) | ( n7487 & ~n7540 ) | ( n7527 & ~n7540 ) ;
  assign n7543 = ( n7540 & ~n7541 ) | ( n7540 & n7542 ) | ( ~n7541 & n7542 ) ;
  assign n7544 = ( n7489 & ~n7529 ) | ( n7489 & n7543 ) | ( ~n7529 & n7543 ) ;
  assign n7545 = ( n7489 & n7529 ) | ( n7489 & n7543 ) | ( n7529 & n7543 ) ;
  assign n7546 = ( n7529 & n7544 ) | ( n7529 & ~n7545 ) | ( n7544 & ~n7545 ) ;
  assign n7547 = x42 & x60 ;
  assign n7548 = x41 & x61 ;
  assign n7549 = x39 & x63 ;
  assign n7550 = ( ~n7547 & n7548 ) | ( ~n7547 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7551 = ( n7547 & n7548 ) | ( n7547 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7552 = ( n7547 & n7550 ) | ( n7547 & ~n7551 ) | ( n7550 & ~n7551 ) ;
  assign n7553 = ( ~n7497 & n7518 ) | ( ~n7497 & n7552 ) | ( n7518 & n7552 ) ;
  assign n7554 = ( n7497 & n7518 ) | ( n7497 & n7552 ) | ( n7518 & n7552 ) ;
  assign n7555 = ( n7497 & n7553 ) | ( n7497 & ~n7554 ) | ( n7553 & ~n7554 ) ;
  assign n7556 = x49 & x53 ;
  assign n7557 = x50 & x52 ;
  assign n7558 = x48 & x54 ;
  assign n7559 = ( ~n7556 & n7557 ) | ( ~n7556 & n7558 ) | ( n7557 & n7558 ) ;
  assign n7560 = ( n7556 & n7557 ) | ( n7556 & n7558 ) | ( n7557 & n7558 ) ;
  assign n7561 = ( n7556 & n7559 ) | ( n7556 & ~n7560 ) | ( n7559 & ~n7560 ) ;
  assign n7562 = x47 & x55 ;
  assign n7563 = x45 & x57 ;
  assign n7564 = x46 & x56 ;
  assign n7565 = ( ~n7562 & n7563 ) | ( ~n7562 & n7564 ) | ( n7563 & n7564 ) ;
  assign n7566 = ( n7562 & n7563 ) | ( n7562 & n7564 ) | ( n7563 & n7564 ) ;
  assign n7567 = ( n7562 & n7565 ) | ( n7562 & ~n7566 ) | ( n7565 & ~n7566 ) ;
  assign n7568 = x43 & x59 ;
  assign n7569 = x40 & x62 ;
  assign n7570 = x44 & x58 ;
  assign n7571 = ( ~n7568 & n7569 ) | ( ~n7568 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7572 = ( n7568 & n7569 ) | ( n7568 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7573 = ( n7568 & n7571 ) | ( n7568 & ~n7572 ) | ( n7571 & ~n7572 ) ;
  assign n7574 = ( ~n7561 & n7567 ) | ( ~n7561 & n7573 ) | ( n7567 & n7573 ) ;
  assign n7575 = ( n7561 & n7567 ) | ( n7561 & n7573 ) | ( n7567 & n7573 ) ;
  assign n7576 = ( n7561 & n7574 ) | ( n7561 & ~n7575 ) | ( n7574 & ~n7575 ) ;
  assign n7577 = ( n7505 & n7555 ) | ( n7505 & n7576 ) | ( n7555 & n7576 ) ;
  assign n7578 = ( n7505 & ~n7555 ) | ( n7505 & n7576 ) | ( ~n7555 & n7576 ) ;
  assign n7579 = ( n7555 & ~n7577 ) | ( n7555 & n7578 ) | ( ~n7577 & n7578 ) ;
  assign n7580 = ( n7493 & n7546 ) | ( n7493 & n7579 ) | ( n7546 & n7579 ) ;
  assign n7581 = ( ~n7493 & n7546 ) | ( ~n7493 & n7579 ) | ( n7546 & n7579 ) ;
  assign n7582 = ( n7493 & ~n7580 ) | ( n7493 & n7581 ) | ( ~n7580 & n7581 ) ;
  assign n7583 = ( n7532 & n7536 ) | ( n7532 & n7582 ) | ( n7536 & n7582 ) ;
  assign n7584 = ( n7532 & ~n7536 ) | ( n7532 & n7582 ) | ( ~n7536 & n7582 ) ;
  assign n7585 = ( n7536 & ~n7583 ) | ( n7536 & n7584 ) | ( ~n7583 & n7584 ) ;
  assign n7586 = ( n7538 & ~n7554 ) | ( n7538 & n7575 ) | ( ~n7554 & n7575 ) ;
  assign n7587 = ( n7538 & n7554 ) | ( n7538 & n7575 ) | ( n7554 & n7575 ) ;
  assign n7588 = ( n7554 & n7586 ) | ( n7554 & ~n7587 ) | ( n7586 & ~n7587 ) ;
  assign n7589 = ( n7541 & n7577 ) | ( n7541 & n7588 ) | ( n7577 & n7588 ) ;
  assign n7590 = ( n7541 & n7577 ) | ( n7541 & ~n7588 ) | ( n7577 & ~n7588 ) ;
  assign n7591 = ( n7588 & ~n7589 ) | ( n7588 & n7590 ) | ( ~n7589 & n7590 ) ;
  assign n7592 = x46 & x57 ;
  assign n7593 = x47 & x56 ;
  assign n7594 = x43 & x60 ;
  assign n7595 = ( ~n7592 & n7593 ) | ( ~n7592 & n7594 ) | ( n7593 & n7594 ) ;
  assign n7596 = ( n7592 & n7593 ) | ( n7592 & n7594 ) | ( n7593 & n7594 ) ;
  assign n7597 = ( n7592 & n7595 ) | ( n7592 & ~n7596 ) | ( n7595 & ~n7596 ) ;
  assign n7598 = x50 & x53 ;
  assign n7599 = x48 & x55 ;
  assign n7600 = x49 & x54 ;
  assign n7601 = ( ~n7598 & n7599 ) | ( ~n7598 & n7600 ) | ( n7599 & n7600 ) ;
  assign n7602 = ( n7598 & n7599 ) | ( n7598 & n7600 ) | ( n7599 & n7600 ) ;
  assign n7603 = ( n7598 & n7601 ) | ( n7598 & ~n7602 ) | ( n7601 & ~n7602 ) ;
  assign n7604 = x41 & x62 ;
  assign n7605 = x51 & x52 ;
  assign n7606 = ( x52 & n7604 ) | ( x52 & n7605 ) | ( n7604 & n7605 ) ;
  assign n7607 = ( x52 & ~n7604 ) | ( x52 & n7605 ) | ( ~n7604 & n7605 ) ;
  assign n7608 = ( n7604 & ~n7606 ) | ( n7604 & n7607 ) | ( ~n7606 & n7607 ) ;
  assign n7609 = ( ~n7597 & n7603 ) | ( ~n7597 & n7608 ) | ( n7603 & n7608 ) ;
  assign n7610 = ( n7597 & n7603 ) | ( n7597 & n7608 ) | ( n7603 & n7608 ) ;
  assign n7611 = ( n7597 & n7609 ) | ( n7597 & ~n7610 ) | ( n7609 & ~n7610 ) ;
  assign n7612 = x45 & x58 ;
  assign n7613 = x44 & x59 ;
  assign n7614 = x42 & x61 ;
  assign n7615 = ( ~n7612 & n7613 ) | ( ~n7612 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7616 = ( n7612 & n7613 ) | ( n7612 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7617 = ( n7612 & n7615 ) | ( n7612 & ~n7616 ) | ( n7615 & ~n7616 ) ;
  assign n7618 = ( n7551 & n7572 ) | ( n7551 & ~n7617 ) | ( n7572 & ~n7617 ) ;
  assign n7619 = ( n7551 & n7572 ) | ( n7551 & n7617 ) | ( n7572 & n7617 ) ;
  assign n7620 = ( n7617 & n7618 ) | ( n7617 & ~n7619 ) | ( n7618 & ~n7619 ) ;
  assign n7621 = x40 & x63 ;
  assign n7622 = ( n7560 & n7566 ) | ( n7560 & n7621 ) | ( n7566 & n7621 ) ;
  assign n7623 = ( ~n7560 & n7566 ) | ( ~n7560 & n7621 ) | ( n7566 & n7621 ) ;
  assign n7624 = ( n7560 & ~n7622 ) | ( n7560 & n7623 ) | ( ~n7622 & n7623 ) ;
  assign n7625 = ( ~n7611 & n7620 ) | ( ~n7611 & n7624 ) | ( n7620 & n7624 ) ;
  assign n7626 = ( n7611 & n7620 ) | ( n7611 & n7624 ) | ( n7620 & n7624 ) ;
  assign n7627 = ( n7611 & n7625 ) | ( n7611 & ~n7626 ) | ( n7625 & ~n7626 ) ;
  assign n7628 = ( n7545 & n7591 ) | ( n7545 & n7627 ) | ( n7591 & n7627 ) ;
  assign n7629 = ( n7545 & ~n7591 ) | ( n7545 & n7627 ) | ( ~n7591 & n7627 ) ;
  assign n7630 = ( n7591 & ~n7628 ) | ( n7591 & n7629 ) | ( ~n7628 & n7629 ) ;
  assign n7631 = ( n7580 & n7583 ) | ( n7580 & n7630 ) | ( n7583 & n7630 ) ;
  assign n7632 = ( n7580 & ~n7583 ) | ( n7580 & n7630 ) | ( ~n7583 & n7630 ) ;
  assign n7633 = ( n7583 & ~n7631 ) | ( n7583 & n7632 ) | ( ~n7631 & n7632 ) ;
  assign n7634 = x42 & x62 ;
  assign n7635 = x41 & x63 ;
  assign n7636 = ( ~n7606 & n7634 ) | ( ~n7606 & n7635 ) | ( n7634 & n7635 ) ;
  assign n7637 = ( n7606 & n7634 ) | ( n7606 & n7635 ) | ( n7634 & n7635 ) ;
  assign n7638 = ( n7606 & n7636 ) | ( n7606 & ~n7637 ) | ( n7636 & ~n7637 ) ;
  assign n7639 = ( n7619 & n7622 ) | ( n7619 & n7638 ) | ( n7622 & n7638 ) ;
  assign n7640 = ( n7619 & n7622 ) | ( n7619 & ~n7638 ) | ( n7622 & ~n7638 ) ;
  assign n7641 = ( n7638 & ~n7639 ) | ( n7638 & n7640 ) | ( ~n7639 & n7640 ) ;
  assign n7642 = ( n7587 & ~n7626 ) | ( n7587 & n7641 ) | ( ~n7626 & n7641 ) ;
  assign n7643 = ( n7587 & n7626 ) | ( n7587 & n7641 ) | ( n7626 & n7641 ) ;
  assign n7644 = ( n7626 & n7642 ) | ( n7626 & ~n7643 ) | ( n7642 & ~n7643 ) ;
  assign n7645 = x48 & x56 ;
  assign n7646 = x47 & x57 ;
  assign n7647 = x46 & x58 ;
  assign n7648 = ( ~n7645 & n7646 ) | ( ~n7645 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7649 = ( n7645 & n7646 ) | ( n7645 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7650 = ( n7645 & n7648 ) | ( n7645 & ~n7649 ) | ( n7648 & ~n7649 ) ;
  assign n7651 = x45 & x59 ;
  assign n7652 = x44 & x60 ;
  assign n7653 = x43 & x61 ;
  assign n7654 = ( ~n7651 & n7652 ) | ( ~n7651 & n7653 ) | ( n7652 & n7653 ) ;
  assign n7655 = ( n7651 & n7652 ) | ( n7651 & n7653 ) | ( n7652 & n7653 ) ;
  assign n7656 = ( n7651 & n7654 ) | ( n7651 & ~n7655 ) | ( n7654 & ~n7655 ) ;
  assign n7657 = x49 & x55 ;
  assign n7658 = x51 & x53 ;
  assign n7659 = x50 & x54 ;
  assign n7660 = ( ~n7657 & n7658 ) | ( ~n7657 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7661 = ( n7657 & n7658 ) | ( n7657 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7662 = ( n7657 & n7660 ) | ( n7657 & ~n7661 ) | ( n7660 & ~n7661 ) ;
  assign n7663 = ( ~n7650 & n7656 ) | ( ~n7650 & n7662 ) | ( n7656 & n7662 ) ;
  assign n7664 = ( n7650 & n7656 ) | ( n7650 & n7662 ) | ( n7656 & n7662 ) ;
  assign n7665 = ( n7650 & n7663 ) | ( n7650 & ~n7664 ) | ( n7663 & ~n7664 ) ;
  assign n7666 = ( ~n7596 & n7602 ) | ( ~n7596 & n7616 ) | ( n7602 & n7616 ) ;
  assign n7667 = ( n7596 & n7602 ) | ( n7596 & n7616 ) | ( n7602 & n7616 ) ;
  assign n7668 = ( n7596 & n7666 ) | ( n7596 & ~n7667 ) | ( n7666 & ~n7667 ) ;
  assign n7669 = ( n7610 & n7665 ) | ( n7610 & n7668 ) | ( n7665 & n7668 ) ;
  assign n7670 = ( n7610 & ~n7665 ) | ( n7610 & n7668 ) | ( ~n7665 & n7668 ) ;
  assign n7671 = ( n7665 & ~n7669 ) | ( n7665 & n7670 ) | ( ~n7669 & n7670 ) ;
  assign n7672 = ( n7589 & n7644 ) | ( n7589 & n7671 ) | ( n7644 & n7671 ) ;
  assign n7673 = ( ~n7589 & n7644 ) | ( ~n7589 & n7671 ) | ( n7644 & n7671 ) ;
  assign n7674 = ( n7589 & ~n7672 ) | ( n7589 & n7673 ) | ( ~n7672 & n7673 ) ;
  assign n7675 = ( n7628 & n7631 ) | ( n7628 & n7674 ) | ( n7631 & n7674 ) ;
  assign n7676 = ( n7628 & ~n7631 ) | ( n7628 & n7674 ) | ( ~n7631 & n7674 ) ;
  assign n7677 = ( n7631 & ~n7675 ) | ( n7631 & n7676 ) | ( ~n7675 & n7676 ) ;
  assign n7678 = x47 & x58 ;
  assign n7679 = x48 & x57 ;
  assign n7680 = x46 & x59 ;
  assign n7681 = ( ~n7678 & n7679 ) | ( ~n7678 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7682 = ( n7678 & n7679 ) | ( n7678 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7683 = ( n7678 & n7681 ) | ( n7678 & ~n7682 ) | ( n7681 & ~n7682 ) ;
  assign n7684 = x45 & x60 ;
  assign n7685 = x42 & x63 ;
  assign n7686 = x44 & x61 ;
  assign n7687 = ( ~n7684 & n7685 ) | ( ~n7684 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7688 = ( n7684 & n7685 ) | ( n7684 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7689 = ( n7684 & n7687 ) | ( n7684 & ~n7688 ) | ( n7687 & ~n7688 ) ;
  assign n7690 = ( ~n7637 & n7683 ) | ( ~n7637 & n7689 ) | ( n7683 & n7689 ) ;
  assign n7691 = ( n7637 & n7683 ) | ( n7637 & n7689 ) | ( n7683 & n7689 ) ;
  assign n7692 = ( n7637 & n7690 ) | ( n7637 & ~n7691 ) | ( n7690 & ~n7691 ) ;
  assign n7693 = x49 & x56 ;
  assign n7694 = x50 & x55 ;
  assign n7695 = x51 & x54 ;
  assign n7696 = ( ~n7693 & n7694 ) | ( ~n7693 & n7695 ) | ( n7694 & n7695 ) ;
  assign n7697 = ( n7693 & n7694 ) | ( n7693 & n7695 ) | ( n7694 & n7695 ) ;
  assign n7698 = ( n7693 & n7696 ) | ( n7693 & ~n7697 ) | ( n7696 & ~n7697 ) ;
  assign n7699 = x43 & x62 ;
  assign n7700 = x52 & x53 ;
  assign n7701 = ( x53 & n7699 ) | ( x53 & n7700 ) | ( n7699 & n7700 ) ;
  assign n7702 = ( x53 & ~n7699 ) | ( x53 & n7700 ) | ( ~n7699 & n7700 ) ;
  assign n7703 = ( n7699 & ~n7701 ) | ( n7699 & n7702 ) | ( ~n7701 & n7702 ) ;
  assign n7704 = ( ~n7667 & n7698 ) | ( ~n7667 & n7703 ) | ( n7698 & n7703 ) ;
  assign n7705 = ( n7667 & n7698 ) | ( n7667 & n7703 ) | ( n7698 & n7703 ) ;
  assign n7706 = ( n7667 & n7704 ) | ( n7667 & ~n7705 ) | ( n7704 & ~n7705 ) ;
  assign n7707 = ( n7669 & n7692 ) | ( n7669 & n7706 ) | ( n7692 & n7706 ) ;
  assign n7708 = ( ~n7669 & n7692 ) | ( ~n7669 & n7706 ) | ( n7692 & n7706 ) ;
  assign n7709 = ( n7669 & ~n7707 ) | ( n7669 & n7708 ) | ( ~n7707 & n7708 ) ;
  assign n7710 = ( n7649 & ~n7655 ) | ( n7649 & n7661 ) | ( ~n7655 & n7661 ) ;
  assign n7711 = ( n7649 & n7655 ) | ( n7649 & n7661 ) | ( n7655 & n7661 ) ;
  assign n7712 = ( n7655 & n7710 ) | ( n7655 & ~n7711 ) | ( n7710 & ~n7711 ) ;
  assign n7713 = ( n7639 & n7664 ) | ( n7639 & n7712 ) | ( n7664 & n7712 ) ;
  assign n7714 = ( ~n7639 & n7664 ) | ( ~n7639 & n7712 ) | ( n7664 & n7712 ) ;
  assign n7715 = ( n7639 & ~n7713 ) | ( n7639 & n7714 ) | ( ~n7713 & n7714 ) ;
  assign n7716 = ( n7643 & n7709 ) | ( n7643 & n7715 ) | ( n7709 & n7715 ) ;
  assign n7717 = ( ~n7643 & n7709 ) | ( ~n7643 & n7715 ) | ( n7709 & n7715 ) ;
  assign n7718 = ( n7643 & ~n7716 ) | ( n7643 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7719 = ( n7672 & n7675 ) | ( n7672 & n7718 ) | ( n7675 & n7718 ) ;
  assign n7720 = ( n7672 & ~n7675 ) | ( n7672 & n7718 ) | ( ~n7675 & n7718 ) ;
  assign n7721 = ( n7675 & ~n7719 ) | ( n7675 & n7720 ) | ( ~n7719 & n7720 ) ;
  assign n7722 = x46 & x60 ;
  assign n7723 = x44 & x62 ;
  assign n7724 = x45 & x61 ;
  assign n7725 = ( ~n7722 & n7723 ) | ( ~n7722 & n7724 ) | ( n7723 & n7724 ) ;
  assign n7726 = ( n7722 & n7723 ) | ( n7722 & n7724 ) | ( n7723 & n7724 ) ;
  assign n7727 = ( n7722 & n7725 ) | ( n7722 & ~n7726 ) | ( n7725 & ~n7726 ) ;
  assign n7728 = ( n7682 & n7688 ) | ( n7682 & ~n7727 ) | ( n7688 & ~n7727 ) ;
  assign n7729 = ( n7682 & n7688 ) | ( n7682 & n7727 ) | ( n7688 & n7727 ) ;
  assign n7730 = ( n7727 & n7728 ) | ( n7727 & ~n7729 ) | ( n7728 & ~n7729 ) ;
  assign n7731 = x51 & x55 ;
  assign n7732 = x52 & x54 ;
  assign n7733 = x50 & x56 ;
  assign n7734 = ( ~n7731 & n7732 ) | ( ~n7731 & n7733 ) | ( n7732 & n7733 ) ;
  assign n7735 = ( n7731 & n7732 ) | ( n7731 & n7733 ) | ( n7732 & n7733 ) ;
  assign n7736 = ( n7731 & n7734 ) | ( n7731 & ~n7735 ) | ( n7734 & ~n7735 ) ;
  assign n7737 = x49 & x57 ;
  assign n7738 = x48 & x58 ;
  assign n7739 = x47 & x59 ;
  assign n7740 = ( ~n7737 & n7738 ) | ( ~n7737 & n7739 ) | ( n7738 & n7739 ) ;
  assign n7741 = ( n7737 & n7738 ) | ( n7737 & n7739 ) | ( n7738 & n7739 ) ;
  assign n7742 = ( n7737 & n7740 ) | ( n7737 & ~n7741 ) | ( n7740 & ~n7741 ) ;
  assign n7743 = ( ~n7711 & n7736 ) | ( ~n7711 & n7742 ) | ( n7736 & n7742 ) ;
  assign n7744 = ( n7711 & n7736 ) | ( n7711 & n7742 ) | ( n7736 & n7742 ) ;
  assign n7745 = ( n7711 & n7743 ) | ( n7711 & ~n7744 ) | ( n7743 & ~n7744 ) ;
  assign n7746 = ( n7713 & n7730 ) | ( n7713 & n7745 ) | ( n7730 & n7745 ) ;
  assign n7747 = ( ~n7713 & n7730 ) | ( ~n7713 & n7745 ) | ( n7730 & n7745 ) ;
  assign n7748 = ( n7713 & ~n7746 ) | ( n7713 & n7747 ) | ( ~n7746 & n7747 ) ;
  assign n7749 = x43 & x63 ;
  assign n7750 = ( n7697 & n7701 ) | ( n7697 & n7749 ) | ( n7701 & n7749 ) ;
  assign n7751 = ( ~n7697 & n7701 ) | ( ~n7697 & n7749 ) | ( n7701 & n7749 ) ;
  assign n7752 = ( n7697 & ~n7750 ) | ( n7697 & n7751 ) | ( ~n7750 & n7751 ) ;
  assign n7753 = ( n7691 & n7705 ) | ( n7691 & n7752 ) | ( n7705 & n7752 ) ;
  assign n7754 = ( n7691 & ~n7705 ) | ( n7691 & n7752 ) | ( ~n7705 & n7752 ) ;
  assign n7755 = ( n7705 & ~n7753 ) | ( n7705 & n7754 ) | ( ~n7753 & n7754 ) ;
  assign n7756 = ( n7707 & n7748 ) | ( n7707 & n7755 ) | ( n7748 & n7755 ) ;
  assign n7757 = ( n7707 & ~n7748 ) | ( n7707 & n7755 ) | ( ~n7748 & n7755 ) ;
  assign n7758 = ( n7748 & ~n7756 ) | ( n7748 & n7757 ) | ( ~n7756 & n7757 ) ;
  assign n7759 = ( n7716 & n7719 ) | ( n7716 & n7758 ) | ( n7719 & n7758 ) ;
  assign n7760 = ( n7716 & ~n7719 ) | ( n7716 & n7758 ) | ( ~n7719 & n7758 ) ;
  assign n7761 = ( n7719 & ~n7759 ) | ( n7719 & n7760 ) | ( ~n7759 & n7760 ) ;
  assign n7762 = ( n7729 & n7744 ) | ( n7729 & n7750 ) | ( n7744 & n7750 ) ;
  assign n7763 = ( n7729 & ~n7744 ) | ( n7729 & n7750 ) | ( ~n7744 & n7750 ) ;
  assign n7764 = ( n7744 & ~n7762 ) | ( n7744 & n7763 ) | ( ~n7762 & n7763 ) ;
  assign n7765 = x47 & x60 ;
  assign n7766 = x46 & x61 ;
  assign n7767 = ( n7735 & n7765 ) | ( n7735 & n7766 ) | ( n7765 & n7766 ) ;
  assign n7768 = ( ~n7735 & n7765 ) | ( ~n7735 & n7766 ) | ( n7765 & n7766 ) ;
  assign n7769 = ( n7735 & ~n7767 ) | ( n7735 & n7768 ) | ( ~n7767 & n7768 ) ;
  assign n7770 = x50 & x57 ;
  assign n7771 = x51 & x56 ;
  assign n7772 = x52 & x55 ;
  assign n7773 = ( ~n7770 & n7771 ) | ( ~n7770 & n7772 ) | ( n7771 & n7772 ) ;
  assign n7774 = ( n7770 & n7771 ) | ( n7770 & n7772 ) | ( n7771 & n7772 ) ;
  assign n7775 = ( n7770 & n7773 ) | ( n7770 & ~n7774 ) | ( n7773 & ~n7774 ) ;
  assign n7776 = x45 & x62 ;
  assign n7777 = x53 & x54 ;
  assign n7778 = ( x54 & n7776 ) | ( x54 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7779 = ( x54 & ~n7776 ) | ( x54 & n7777 ) | ( ~n7776 & n7777 ) ;
  assign n7780 = ( n7776 & ~n7778 ) | ( n7776 & n7779 ) | ( ~n7778 & n7779 ) ;
  assign n7781 = ( n7769 & n7775 ) | ( n7769 & n7780 ) | ( n7775 & n7780 ) ;
  assign n7782 = ( ~n7769 & n7775 ) | ( ~n7769 & n7780 ) | ( n7775 & n7780 ) ;
  assign n7783 = ( n7769 & ~n7781 ) | ( n7769 & n7782 ) | ( ~n7781 & n7782 ) ;
  assign n7784 = x48 & x59 ;
  assign n7785 = x49 & x58 ;
  assign n7786 = ( ~n6675 & n7784 ) | ( ~n6675 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7787 = ( n6675 & n7784 ) | ( n6675 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7788 = ( n6675 & n7786 ) | ( n6675 & ~n7787 ) | ( n7786 & ~n7787 ) ;
  assign n7789 = ( n7726 & n7741 ) | ( n7726 & ~n7788 ) | ( n7741 & ~n7788 ) ;
  assign n7790 = ( n7726 & n7741 ) | ( n7726 & n7788 ) | ( n7741 & n7788 ) ;
  assign n7791 = ( n7788 & n7789 ) | ( n7788 & ~n7790 ) | ( n7789 & ~n7790 ) ;
  assign n7792 = ( n7753 & n7783 ) | ( n7753 & n7791 ) | ( n7783 & n7791 ) ;
  assign n7793 = ( ~n7753 & n7783 ) | ( ~n7753 & n7791 ) | ( n7783 & n7791 ) ;
  assign n7794 = ( n7753 & ~n7792 ) | ( n7753 & n7793 ) | ( ~n7792 & n7793 ) ;
  assign n7795 = ( n7746 & n7764 ) | ( n7746 & n7794 ) | ( n7764 & n7794 ) ;
  assign n7796 = ( n7746 & ~n7764 ) | ( n7746 & n7794 ) | ( ~n7764 & n7794 ) ;
  assign n7797 = ( n7764 & ~n7795 ) | ( n7764 & n7796 ) | ( ~n7795 & n7796 ) ;
  assign n7798 = ( n7756 & ~n7759 ) | ( n7756 & n7797 ) | ( ~n7759 & n7797 ) ;
  assign n7799 = ( n7756 & n7759 ) | ( n7756 & n7797 ) | ( n7759 & n7797 ) ;
  assign n7800 = ( n7759 & n7798 ) | ( n7759 & ~n7799 ) | ( n7798 & ~n7799 ) ;
  assign n7801 = x50 & x58 ;
  assign n7802 = x49 & x59 ;
  assign n7803 = x48 & x60 ;
  assign n7804 = ( ~n7801 & n7802 ) | ( ~n7801 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7805 = ( n7801 & n7802 ) | ( n7801 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7806 = ( n7801 & n7804 ) | ( n7801 & ~n7805 ) | ( n7804 & ~n7805 ) ;
  assign n7807 = x45 & x63 ;
  assign n7808 = x46 & x62 ;
  assign n7809 = x47 & x61 ;
  assign n7810 = ( ~n7807 & n7808 ) | ( ~n7807 & n7809 ) | ( n7808 & n7809 ) ;
  assign n7811 = ( n7807 & n7808 ) | ( n7807 & n7809 ) | ( n7808 & n7809 ) ;
  assign n7812 = ( n7807 & n7810 ) | ( n7807 & ~n7811 ) | ( n7810 & ~n7811 ) ;
  assign n7813 = ( ~n7767 & n7806 ) | ( ~n7767 & n7812 ) | ( n7806 & n7812 ) ;
  assign n7814 = ( n7767 & n7806 ) | ( n7767 & n7812 ) | ( n7806 & n7812 ) ;
  assign n7815 = ( n7767 & n7813 ) | ( n7767 & ~n7814 ) | ( n7813 & ~n7814 ) ;
  assign n7816 = ( n7774 & n7778 ) | ( n7774 & n7787 ) | ( n7778 & n7787 ) ;
  assign n7817 = ( n7774 & ~n7778 ) | ( n7774 & n7787 ) | ( ~n7778 & n7787 ) ;
  assign n7818 = ( n7778 & ~n7816 ) | ( n7778 & n7817 ) | ( ~n7816 & n7817 ) ;
  assign n7819 = ( n7762 & n7815 ) | ( n7762 & n7818 ) | ( n7815 & n7818 ) ;
  assign n7820 = ( ~n7762 & n7815 ) | ( ~n7762 & n7818 ) | ( n7815 & n7818 ) ;
  assign n7821 = ( n7762 & ~n7819 ) | ( n7762 & n7820 ) | ( ~n7819 & n7820 ) ;
  assign n7822 = x53 & x55 ;
  assign n7823 = x52 & x56 ;
  assign n7824 = x51 & x57 ;
  assign n7825 = ( ~n7822 & n7823 ) | ( ~n7822 & n7824 ) | ( n7823 & n7824 ) ;
  assign n7826 = ( n7822 & n7823 ) | ( n7822 & n7824 ) | ( n7823 & n7824 ) ;
  assign n7827 = ( n7822 & n7825 ) | ( n7822 & ~n7826 ) | ( n7825 & ~n7826 ) ;
  assign n7828 = ( n7781 & n7790 ) | ( n7781 & n7827 ) | ( n7790 & n7827 ) ;
  assign n7829 = ( ~n7781 & n7790 ) | ( ~n7781 & n7827 ) | ( n7790 & n7827 ) ;
  assign n7830 = ( n7781 & ~n7828 ) | ( n7781 & n7829 ) | ( ~n7828 & n7829 ) ;
  assign n7831 = ( ~n7792 & n7821 ) | ( ~n7792 & n7830 ) | ( n7821 & n7830 ) ;
  assign n7832 = ( n7792 & n7821 ) | ( n7792 & n7830 ) | ( n7821 & n7830 ) ;
  assign n7833 = ( n7792 & n7831 ) | ( n7792 & ~n7832 ) | ( n7831 & ~n7832 ) ;
  assign n7834 = ( n7795 & ~n7799 ) | ( n7795 & n7833 ) | ( ~n7799 & n7833 ) ;
  assign n7835 = ( n7795 & n7799 ) | ( n7795 & n7833 ) | ( n7799 & n7833 ) ;
  assign n7836 = ( n7799 & n7834 ) | ( n7799 & ~n7835 ) | ( n7834 & ~n7835 ) ;
  assign n7837 = x48 & x61 ;
  assign n7838 = x50 & x59 ;
  assign n7839 = x49 & x60 ;
  assign n7840 = ( ~n7837 & n7838 ) | ( ~n7837 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7841 = ( n7837 & n7838 ) | ( n7837 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7842 = ( n7837 & n7840 ) | ( n7837 & ~n7841 ) | ( n7840 & ~n7841 ) ;
  assign n7843 = x51 & x58 ;
  assign n7844 = x53 & x56 ;
  assign n7845 = x52 & x57 ;
  assign n7846 = ( ~n7843 & n7844 ) | ( ~n7843 & n7845 ) | ( n7844 & n7845 ) ;
  assign n7847 = ( n7843 & n7844 ) | ( n7843 & n7845 ) | ( n7844 & n7845 ) ;
  assign n7848 = ( n7843 & n7846 ) | ( n7843 & ~n7847 ) | ( n7846 & ~n7847 ) ;
  assign n7849 = ( n7811 & ~n7842 ) | ( n7811 & n7848 ) | ( ~n7842 & n7848 ) ;
  assign n7850 = ( n7811 & n7842 ) | ( n7811 & n7848 ) | ( n7842 & n7848 ) ;
  assign n7851 = ( n7842 & n7849 ) | ( n7842 & ~n7850 ) | ( n7849 & ~n7850 ) ;
  assign n7852 = x46 & x63 ;
  assign n7853 = ( n7805 & n7826 ) | ( n7805 & n7852 ) | ( n7826 & n7852 ) ;
  assign n7854 = ( ~n7805 & n7826 ) | ( ~n7805 & n7852 ) | ( n7826 & n7852 ) ;
  assign n7855 = ( n7805 & ~n7853 ) | ( n7805 & n7854 ) | ( ~n7853 & n7854 ) ;
  assign n7856 = ( n7828 & n7851 ) | ( n7828 & n7855 ) | ( n7851 & n7855 ) ;
  assign n7857 = ( ~n7828 & n7851 ) | ( ~n7828 & n7855 ) | ( n7851 & n7855 ) ;
  assign n7858 = ( n7828 & ~n7856 ) | ( n7828 & n7857 ) | ( ~n7856 & n7857 ) ;
  assign n7859 = x47 & x62 ;
  assign n7860 = x54 & x55 ;
  assign n7861 = ( x55 & n7859 ) | ( x55 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7862 = ( x55 & ~n7859 ) | ( x55 & n7860 ) | ( ~n7859 & n7860 ) ;
  assign n7863 = ( n7859 & ~n7861 ) | ( n7859 & n7862 ) | ( ~n7861 & n7862 ) ;
  assign n7864 = ( ~n7814 & n7816 ) | ( ~n7814 & n7863 ) | ( n7816 & n7863 ) ;
  assign n7865 = ( n7814 & n7816 ) | ( n7814 & n7863 ) | ( n7816 & n7863 ) ;
  assign n7866 = ( n7814 & n7864 ) | ( n7814 & ~n7865 ) | ( n7864 & ~n7865 ) ;
  assign n7867 = ( n7819 & n7858 ) | ( n7819 & n7866 ) | ( n7858 & n7866 ) ;
  assign n7868 = ( n7819 & ~n7858 ) | ( n7819 & n7866 ) | ( ~n7858 & n7866 ) ;
  assign n7869 = ( n7858 & ~n7867 ) | ( n7858 & n7868 ) | ( ~n7867 & n7868 ) ;
  assign n7870 = ( n7832 & ~n7835 ) | ( n7832 & n7869 ) | ( ~n7835 & n7869 ) ;
  assign n7871 = ( n7832 & n7835 ) | ( n7832 & n7869 ) | ( n7835 & n7869 ) ;
  assign n7872 = ( n7835 & n7870 ) | ( n7835 & ~n7871 ) | ( n7870 & ~n7871 ) ;
  assign n7873 = x51 & x59 ;
  assign n7874 = x50 & x60 ;
  assign n7875 = x49 & x61 ;
  assign n7876 = ( ~n7873 & n7874 ) | ( ~n7873 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7877 = ( n7873 & n7874 ) | ( n7873 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7878 = ( n7873 & n7876 ) | ( n7873 & ~n7877 ) | ( n7876 & ~n7877 ) ;
  assign n7879 = ( n7841 & n7847 ) | ( n7841 & ~n7878 ) | ( n7847 & ~n7878 ) ;
  assign n7880 = ( n7841 & n7847 ) | ( n7841 & n7878 ) | ( n7847 & n7878 ) ;
  assign n7881 = ( n7878 & n7879 ) | ( n7878 & ~n7880 ) | ( n7879 & ~n7880 ) ;
  assign n7882 = ( n7850 & n7865 ) | ( n7850 & n7881 ) | ( n7865 & n7881 ) ;
  assign n7883 = ( n7850 & n7865 ) | ( n7850 & ~n7881 ) | ( n7865 & ~n7881 ) ;
  assign n7884 = ( n7881 & ~n7882 ) | ( n7881 & n7883 ) | ( ~n7882 & n7883 ) ;
  assign n7885 = x48 & x62 ;
  assign n7886 = x47 & x63 ;
  assign n7887 = ( ~n7861 & n7885 ) | ( ~n7861 & n7886 ) | ( n7885 & n7886 ) ;
  assign n7888 = ( n7861 & n7885 ) | ( n7861 & n7886 ) | ( n7885 & n7886 ) ;
  assign n7889 = ( n7861 & n7887 ) | ( n7861 & ~n7888 ) | ( n7887 & ~n7888 ) ;
  assign n7890 = x53 & x57 ;
  assign n7891 = x54 & x56 ;
  assign n7892 = x52 & x58 ;
  assign n7893 = ( ~n7890 & n7891 ) | ( ~n7890 & n7892 ) | ( n7891 & n7892 ) ;
  assign n7894 = ( n7890 & n7891 ) | ( n7890 & n7892 ) | ( n7891 & n7892 ) ;
  assign n7895 = ( n7890 & n7893 ) | ( n7890 & ~n7894 ) | ( n7893 & ~n7894 ) ;
  assign n7896 = ( ~n7853 & n7889 ) | ( ~n7853 & n7895 ) | ( n7889 & n7895 ) ;
  assign n7897 = ( n7853 & n7889 ) | ( n7853 & n7895 ) | ( n7889 & n7895 ) ;
  assign n7898 = ( n7853 & n7896 ) | ( n7853 & ~n7897 ) | ( n7896 & ~n7897 ) ;
  assign n7899 = ( n7856 & ~n7884 ) | ( n7856 & n7898 ) | ( ~n7884 & n7898 ) ;
  assign n7900 = ( n7856 & n7884 ) | ( n7856 & n7898 ) | ( n7884 & n7898 ) ;
  assign n7901 = ( n7884 & n7899 ) | ( n7884 & ~n7900 ) | ( n7899 & ~n7900 ) ;
  assign n7902 = ( n7867 & n7871 ) | ( n7867 & n7901 ) | ( n7871 & n7901 ) ;
  assign n7903 = ( n7867 & ~n7871 ) | ( n7867 & n7901 ) | ( ~n7871 & n7901 ) ;
  assign n7904 = ( n7871 & ~n7902 ) | ( n7871 & n7903 ) | ( ~n7902 & n7903 ) ;
  assign n7905 = x49 & x62 ;
  assign n7906 = x55 & x56 ;
  assign n7907 = ( x56 & n7905 ) | ( x56 & n7906 ) | ( n7905 & n7906 ) ;
  assign n7908 = ( x56 & ~n7905 ) | ( x56 & n7906 ) | ( ~n7905 & n7906 ) ;
  assign n7909 = ( n7905 & ~n7907 ) | ( n7905 & n7908 ) | ( ~n7907 & n7908 ) ;
  assign n7910 = x50 & x61 ;
  assign n7911 = x48 & x63 ;
  assign n7912 = x51 & x60 ;
  assign n7913 = ( ~n7910 & n7911 ) | ( ~n7910 & n7912 ) | ( n7911 & n7912 ) ;
  assign n7914 = ( n7910 & n7911 ) | ( n7910 & n7912 ) | ( n7911 & n7912 ) ;
  assign n7915 = ( n7910 & n7913 ) | ( n7910 & ~n7914 ) | ( n7913 & ~n7914 ) ;
  assign n7916 = x54 & x57 ;
  assign n7917 = x53 & x58 ;
  assign n7918 = x52 & x59 ;
  assign n7919 = ( ~n7916 & n7917 ) | ( ~n7916 & n7918 ) | ( n7917 & n7918 ) ;
  assign n7920 = ( n7916 & n7917 ) | ( n7916 & n7918 ) | ( n7917 & n7918 ) ;
  assign n7921 = ( n7916 & n7919 ) | ( n7916 & ~n7920 ) | ( n7919 & ~n7920 ) ;
  assign n7922 = ( ~n7909 & n7915 ) | ( ~n7909 & n7921 ) | ( n7915 & n7921 ) ;
  assign n7923 = ( n7909 & n7915 ) | ( n7909 & n7921 ) | ( n7915 & n7921 ) ;
  assign n7924 = ( n7909 & n7922 ) | ( n7909 & ~n7923 ) | ( n7922 & ~n7923 ) ;
  assign n7925 = ( n7877 & ~n7888 ) | ( n7877 & n7894 ) | ( ~n7888 & n7894 ) ;
  assign n7926 = ( n7877 & n7888 ) | ( n7877 & n7894 ) | ( n7888 & n7894 ) ;
  assign n7927 = ( n7888 & n7925 ) | ( n7888 & ~n7926 ) | ( n7925 & ~n7926 ) ;
  assign n7928 = ( n7880 & n7897 ) | ( n7880 & n7927 ) | ( n7897 & n7927 ) ;
  assign n7929 = ( n7880 & n7897 ) | ( n7880 & ~n7927 ) | ( n7897 & ~n7927 ) ;
  assign n7930 = ( n7927 & ~n7928 ) | ( n7927 & n7929 ) | ( ~n7928 & n7929 ) ;
  assign n7931 = ( n7882 & n7924 ) | ( n7882 & n7930 ) | ( n7924 & n7930 ) ;
  assign n7932 = ( ~n7882 & n7924 ) | ( ~n7882 & n7930 ) | ( n7924 & n7930 ) ;
  assign n7933 = ( n7882 & ~n7931 ) | ( n7882 & n7932 ) | ( ~n7931 & n7932 ) ;
  assign n7934 = ( n7900 & n7902 ) | ( n7900 & n7933 ) | ( n7902 & n7933 ) ;
  assign n7935 = ( n7900 & ~n7902 ) | ( n7900 & n7933 ) | ( ~n7902 & n7933 ) ;
  assign n7936 = ( n7902 & ~n7934 ) | ( n7902 & n7935 ) | ( ~n7934 & n7935 ) ;
  assign n7937 = x55 & x57 ;
  assign n7938 = x53 & x59 ;
  assign n7939 = x54 & x58 ;
  assign n7940 = ( ~n7937 & n7938 ) | ( ~n7937 & n7939 ) | ( n7938 & n7939 ) ;
  assign n7941 = ( n7937 & n7938 ) | ( n7937 & n7939 ) | ( n7938 & n7939 ) ;
  assign n7942 = ( n7937 & n7940 ) | ( n7937 & ~n7941 ) | ( n7940 & ~n7941 ) ;
  assign n7943 = x51 & x61 ;
  assign n7944 = x49 & x63 ;
  assign n7945 = x52 & x60 ;
  assign n7946 = ( ~n7943 & n7944 ) | ( ~n7943 & n7945 ) | ( n7944 & n7945 ) ;
  assign n7947 = ( n7943 & n7944 ) | ( n7943 & n7945 ) | ( n7944 & n7945 ) ;
  assign n7948 = ( n7943 & n7946 ) | ( n7943 & ~n7947 ) | ( n7946 & ~n7947 ) ;
  assign n7949 = ( ~n7914 & n7942 ) | ( ~n7914 & n7948 ) | ( n7942 & n7948 ) ;
  assign n7950 = ( n7914 & n7942 ) | ( n7914 & n7948 ) | ( n7942 & n7948 ) ;
  assign n7951 = ( n7914 & n7949 ) | ( n7914 & ~n7950 ) | ( n7949 & ~n7950 ) ;
  assign n7952 = x50 & x62 ;
  assign n7953 = ( n7907 & n7920 ) | ( n7907 & n7952 ) | ( n7920 & n7952 ) ;
  assign n7954 = ( n7907 & ~n7920 ) | ( n7907 & n7952 ) | ( ~n7920 & n7952 ) ;
  assign n7955 = ( n7920 & ~n7953 ) | ( n7920 & n7954 ) | ( ~n7953 & n7954 ) ;
  assign n7956 = ( n7923 & n7926 ) | ( n7923 & n7955 ) | ( n7926 & n7955 ) ;
  assign n7957 = ( n7923 & ~n7926 ) | ( n7923 & n7955 ) | ( ~n7926 & n7955 ) ;
  assign n7958 = ( n7926 & ~n7956 ) | ( n7926 & n7957 ) | ( ~n7956 & n7957 ) ;
  assign n7959 = ( n7928 & n7951 ) | ( n7928 & n7958 ) | ( n7951 & n7958 ) ;
  assign n7960 = ( ~n7928 & n7951 ) | ( ~n7928 & n7958 ) | ( n7951 & n7958 ) ;
  assign n7961 = ( n7928 & ~n7959 ) | ( n7928 & n7960 ) | ( ~n7959 & n7960 ) ;
  assign n7962 = ( n7931 & n7934 ) | ( n7931 & n7961 ) | ( n7934 & n7961 ) ;
  assign n7963 = ( n7931 & ~n7934 ) | ( n7931 & n7961 ) | ( ~n7934 & n7961 ) ;
  assign n7964 = ( n7934 & ~n7962 ) | ( n7934 & n7963 ) | ( ~n7962 & n7963 ) ;
  assign n7965 = x53 & x60 ;
  assign n7966 = x52 & x61 ;
  assign n7967 = ( n7941 & n7965 ) | ( n7941 & n7966 ) | ( n7965 & n7966 ) ;
  assign n7968 = ( ~n7941 & n7965 ) | ( ~n7941 & n7966 ) | ( n7965 & n7966 ) ;
  assign n7969 = ( n7941 & ~n7967 ) | ( n7941 & n7968 ) | ( ~n7967 & n7968 ) ;
  assign n7970 = ( n7950 & n7953 ) | ( n7950 & n7969 ) | ( n7953 & n7969 ) ;
  assign n7971 = ( n7950 & n7953 ) | ( n7950 & ~n7969 ) | ( n7953 & ~n7969 ) ;
  assign n7972 = ( n7969 & ~n7970 ) | ( n7969 & n7971 ) | ( ~n7970 & n7971 ) ;
  assign n7973 = x50 & x63 ;
  assign n7974 = x55 & x58 ;
  assign n7975 = x54 & x59 ;
  assign n7976 = ( ~n7973 & n7974 ) | ( ~n7973 & n7975 ) | ( n7974 & n7975 ) ;
  assign n7977 = ( n7973 & n7974 ) | ( n7973 & n7975 ) | ( n7974 & n7975 ) ;
  assign n7978 = ( n7973 & n7976 ) | ( n7973 & ~n7977 ) | ( n7976 & ~n7977 ) ;
  assign n7979 = x51 & x62 ;
  assign n7980 = x56 & x57 ;
  assign n7981 = ( x57 & n7979 ) | ( x57 & n7980 ) | ( n7979 & n7980 ) ;
  assign n7982 = ( x57 & ~n7979 ) | ( x57 & n7980 ) | ( ~n7979 & n7980 ) ;
  assign n7983 = ( n7979 & ~n7981 ) | ( n7979 & n7982 ) | ( ~n7981 & n7982 ) ;
  assign n7984 = ( n7947 & ~n7978 ) | ( n7947 & n7983 ) | ( ~n7978 & n7983 ) ;
  assign n7985 = ( n7947 & n7978 ) | ( n7947 & n7983 ) | ( n7978 & n7983 ) ;
  assign n7986 = ( n7978 & n7984 ) | ( n7978 & ~n7985 ) | ( n7984 & ~n7985 ) ;
  assign n7987 = ( n7956 & ~n7972 ) | ( n7956 & n7986 ) | ( ~n7972 & n7986 ) ;
  assign n7988 = ( n7956 & n7972 ) | ( n7956 & n7986 ) | ( n7972 & n7986 ) ;
  assign n7989 = ( n7972 & n7987 ) | ( n7972 & ~n7988 ) | ( n7987 & ~n7988 ) ;
  assign n7990 = ( n7959 & n7962 ) | ( n7959 & n7989 ) | ( n7962 & n7989 ) ;
  assign n7991 = ( n7959 & ~n7962 ) | ( n7959 & n7989 ) | ( ~n7962 & n7989 ) ;
  assign n7992 = ( n7962 & ~n7990 ) | ( n7962 & n7991 ) | ( ~n7990 & n7991 ) ;
  assign n7993 = x56 & x58 ;
  assign n7994 = x55 & x59 ;
  assign n7995 = x54 & x60 ;
  assign n7996 = ( ~n7993 & n7994 ) | ( ~n7993 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7997 = ( n7993 & n7994 ) | ( n7993 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7998 = ( n7993 & n7996 ) | ( n7993 & ~n7997 ) | ( n7996 & ~n7997 ) ;
  assign n7999 = x51 & x63 ;
  assign n8000 = x52 & x62 ;
  assign n8001 = x53 & x61 ;
  assign n8002 = ( ~n7999 & n8000 ) | ( ~n7999 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8003 = ( n7999 & n8000 ) | ( n7999 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8004 = ( n7999 & n8002 ) | ( n7999 & ~n8003 ) | ( n8002 & ~n8003 ) ;
  assign n8005 = ( ~n7985 & n7998 ) | ( ~n7985 & n8004 ) | ( n7998 & n8004 ) ;
  assign n8006 = ( n7985 & n7998 ) | ( n7985 & n8004 ) | ( n7998 & n8004 ) ;
  assign n8007 = ( n7985 & n8005 ) | ( n7985 & ~n8006 ) | ( n8005 & ~n8006 ) ;
  assign n8008 = ( n7967 & n7977 ) | ( n7967 & n7981 ) | ( n7977 & n7981 ) ;
  assign n8009 = ( ~n7967 & n7977 ) | ( ~n7967 & n7981 ) | ( n7977 & n7981 ) ;
  assign n8010 = ( n7967 & ~n8008 ) | ( n7967 & n8009 ) | ( ~n8008 & n8009 ) ;
  assign n8011 = ( n7970 & n8007 ) | ( n7970 & n8010 ) | ( n8007 & n8010 ) ;
  assign n8012 = ( n7970 & ~n8007 ) | ( n7970 & n8010 ) | ( ~n8007 & n8010 ) ;
  assign n8013 = ( n8007 & ~n8011 ) | ( n8007 & n8012 ) | ( ~n8011 & n8012 ) ;
  assign n8014 = ( n7988 & ~n7990 ) | ( n7988 & n8013 ) | ( ~n7990 & n8013 ) ;
  assign n8015 = ( n7988 & n7990 ) | ( n7988 & n8013 ) | ( n7990 & n8013 ) ;
  assign n8016 = ( n7990 & n8014 ) | ( n7990 & ~n8015 ) | ( n8014 & ~n8015 ) ;
  assign n8017 = x56 & x59 ;
  assign n8018 = x55 & x60 ;
  assign n8019 = x54 & x61 ;
  assign n8020 = ( ~n8017 & n8018 ) | ( ~n8017 & n8019 ) | ( n8018 & n8019 ) ;
  assign n8021 = ( n8017 & n8018 ) | ( n8017 & n8019 ) | ( n8018 & n8019 ) ;
  assign n8022 = ( n8017 & n8020 ) | ( n8017 & ~n8021 ) | ( n8020 & ~n8021 ) ;
  assign n8023 = x53 & x62 ;
  assign n8024 = x57 & x58 ;
  assign n8025 = ( x58 & n8023 ) | ( x58 & n8024 ) | ( n8023 & n8024 ) ;
  assign n8026 = ( x58 & ~n8023 ) | ( x58 & n8024 ) | ( ~n8023 & n8024 ) ;
  assign n8027 = ( n8023 & ~n8025 ) | ( n8023 & n8026 ) | ( ~n8025 & n8026 ) ;
  assign n8028 = ( ~n8008 & n8022 ) | ( ~n8008 & n8027 ) | ( n8022 & n8027 ) ;
  assign n8029 = ( n8008 & n8022 ) | ( n8008 & n8027 ) | ( n8022 & n8027 ) ;
  assign n8030 = ( n8008 & n8028 ) | ( n8008 & ~n8029 ) | ( n8028 & ~n8029 ) ;
  assign n8031 = x52 & x63 ;
  assign n8032 = ( n7997 & n8003 ) | ( n7997 & n8031 ) | ( n8003 & n8031 ) ;
  assign n8033 = ( ~n7997 & n8003 ) | ( ~n7997 & n8031 ) | ( n8003 & n8031 ) ;
  assign n8034 = ( n7997 & ~n8032 ) | ( n7997 & n8033 ) | ( ~n8032 & n8033 ) ;
  assign n8035 = ( n8006 & n8030 ) | ( n8006 & n8034 ) | ( n8030 & n8034 ) ;
  assign n8036 = ( n8006 & ~n8030 ) | ( n8006 & n8034 ) | ( ~n8030 & n8034 ) ;
  assign n8037 = ( n8030 & ~n8035 ) | ( n8030 & n8036 ) | ( ~n8035 & n8036 ) ;
  assign n8038 = ( n8011 & ~n8015 ) | ( n8011 & n8037 ) | ( ~n8015 & n8037 ) ;
  assign n8039 = ( n8011 & n8015 ) | ( n8011 & n8037 ) | ( n8015 & n8037 ) ;
  assign n8040 = ( n8015 & n8038 ) | ( n8015 & ~n8039 ) | ( n8038 & ~n8039 ) ;
  assign n8041 = x54 & x62 ;
  assign n8042 = x53 & x63 ;
  assign n8043 = ( ~n8025 & n8041 ) | ( ~n8025 & n8042 ) | ( n8041 & n8042 ) ;
  assign n8044 = ( n8025 & n8041 ) | ( n8025 & n8042 ) | ( n8041 & n8042 ) ;
  assign n8045 = ( n8025 & n8043 ) | ( n8025 & ~n8044 ) | ( n8043 & ~n8044 ) ;
  assign n8046 = x57 & x59 ;
  assign n8047 = x56 & x60 ;
  assign n8048 = x55 & x61 ;
  assign n8049 = ( ~n8046 & n8047 ) | ( ~n8046 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8050 = ( n8046 & n8047 ) | ( n8046 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8051 = ( n8046 & n8049 ) | ( n8046 & ~n8050 ) | ( n8049 & ~n8050 ) ;
  assign n8052 = ( n8021 & ~n8045 ) | ( n8021 & n8051 ) | ( ~n8045 & n8051 ) ;
  assign n8053 = ( n8021 & n8045 ) | ( n8021 & n8051 ) | ( n8045 & n8051 ) ;
  assign n8054 = ( n8045 & n8052 ) | ( n8045 & ~n8053 ) | ( n8052 & ~n8053 ) ;
  assign n8055 = ( ~n8029 & n8032 ) | ( ~n8029 & n8054 ) | ( n8032 & n8054 ) ;
  assign n8056 = ( n8029 & n8032 ) | ( n8029 & n8054 ) | ( n8032 & n8054 ) ;
  assign n8057 = ( n8029 & n8055 ) | ( n8029 & ~n8056 ) | ( n8055 & ~n8056 ) ;
  assign n8058 = ( n8035 & n8039 ) | ( n8035 & n8057 ) | ( n8039 & n8057 ) ;
  assign n8059 = ( n8035 & ~n8039 ) | ( n8035 & n8057 ) | ( ~n8039 & n8057 ) ;
  assign n8060 = ( n8039 & ~n8058 ) | ( n8039 & n8059 ) | ( ~n8058 & n8059 ) ;
  assign n8061 = x54 & x63 ;
  assign n8062 = x57 & x60 ;
  assign n8063 = x56 & x61 ;
  assign n8064 = ( ~n8061 & n8062 ) | ( ~n8061 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8065 = ( n8061 & n8062 ) | ( n8061 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8066 = ( n8061 & n8064 ) | ( n8061 & ~n8065 ) | ( n8064 & ~n8065 ) ;
  assign n8067 = ( ~n8044 & n8050 ) | ( ~n8044 & n8066 ) | ( n8050 & n8066 ) ;
  assign n8068 = ( n8044 & n8050 ) | ( n8044 & n8066 ) | ( n8050 & n8066 ) ;
  assign n8069 = ( n8044 & n8067 ) | ( n8044 & ~n8068 ) | ( n8067 & ~n8068 ) ;
  assign n8070 = x55 & x62 ;
  assign n8071 = x58 & x59 ;
  assign n8072 = ( x59 & n8070 ) | ( x59 & n8071 ) | ( n8070 & n8071 ) ;
  assign n8073 = ( x59 & ~n8070 ) | ( x59 & n8071 ) | ( ~n8070 & n8071 ) ;
  assign n8074 = ( n8070 & ~n8072 ) | ( n8070 & n8073 ) | ( ~n8072 & n8073 ) ;
  assign n8075 = ( ~n8053 & n8069 ) | ( ~n8053 & n8074 ) | ( n8069 & n8074 ) ;
  assign n8076 = ( n8053 & n8069 ) | ( n8053 & n8074 ) | ( n8069 & n8074 ) ;
  assign n8077 = ( n8053 & n8075 ) | ( n8053 & ~n8076 ) | ( n8075 & ~n8076 ) ;
  assign n8078 = ( n8056 & ~n8058 ) | ( n8056 & n8077 ) | ( ~n8058 & n8077 ) ;
  assign n8079 = ( n8056 & n8058 ) | ( n8056 & n8077 ) | ( n8058 & n8077 ) ;
  assign n8080 = ( n8058 & n8078 ) | ( n8058 & ~n8079 ) | ( n8078 & ~n8079 ) ;
  assign n8081 = x55 & x63 ;
  assign n8082 = ( n8065 & n8072 ) | ( n8065 & n8081 ) | ( n8072 & n8081 ) ;
  assign n8083 = ( ~n8065 & n8072 ) | ( ~n8065 & n8081 ) | ( n8072 & n8081 ) ;
  assign n8084 = ( n8065 & ~n8082 ) | ( n8065 & n8083 ) | ( ~n8082 & n8083 ) ;
  assign n8085 = x58 & x60 ;
  assign n8086 = x56 & x62 ;
  assign n8087 = x57 & x61 ;
  assign n8088 = ( ~n8085 & n8086 ) | ( ~n8085 & n8087 ) | ( n8086 & n8087 ) ;
  assign n8089 = ( n8085 & n8086 ) | ( n8085 & n8087 ) | ( n8086 & n8087 ) ;
  assign n8090 = ( n8085 & n8088 ) | ( n8085 & ~n8089 ) | ( n8088 & ~n8089 ) ;
  assign n8091 = ( n8068 & n8084 ) | ( n8068 & n8090 ) | ( n8084 & n8090 ) ;
  assign n8092 = ( ~n8068 & n8084 ) | ( ~n8068 & n8090 ) | ( n8084 & n8090 ) ;
  assign n8093 = ( n8068 & ~n8091 ) | ( n8068 & n8092 ) | ( ~n8091 & n8092 ) ;
  assign n8094 = ( n8076 & ~n8079 ) | ( n8076 & n8093 ) | ( ~n8079 & n8093 ) ;
  assign n8095 = ( n8076 & n8079 ) | ( n8076 & n8093 ) | ( n8079 & n8093 ) ;
  assign n8096 = ( n8079 & n8094 ) | ( n8079 & ~n8095 ) | ( n8094 & ~n8095 ) ;
  assign n8097 = n8062 & ~n8086 ;
  assign n8098 = x58 & x61 ;
  assign n8099 = ~n8097 & n8098 ;
  assign n8100 = x56 & x63 ;
  assign n8101 = n8086 & n8089 ;
  assign n8102 = ( ~n8099 & n8100 ) | ( ~n8099 & n8101 ) | ( n8100 & n8101 ) ;
  assign n8103 = ( n8099 & n8100 ) | ( n8099 & n8101 ) | ( n8100 & n8101 ) ;
  assign n8104 = ( n8099 & n8102 ) | ( n8099 & ~n8103 ) | ( n8102 & ~n8103 ) ;
  assign n8105 = x57 & x62 ;
  assign n8106 = x59 & x60 ;
  assign n8107 = ( x60 & n8105 ) | ( x60 & n8106 ) | ( n8105 & n8106 ) ;
  assign n8108 = ( x60 & ~n8105 ) | ( x60 & n8106 ) | ( ~n8105 & n8106 ) ;
  assign n8109 = ( n8105 & ~n8107 ) | ( n8105 & n8108 ) | ( ~n8107 & n8108 ) ;
  assign n8110 = ( n8082 & ~n8104 ) | ( n8082 & n8109 ) | ( ~n8104 & n8109 ) ;
  assign n8111 = ( n8082 & n8104 ) | ( n8082 & n8109 ) | ( n8104 & n8109 ) ;
  assign n8112 = ( n8104 & n8110 ) | ( n8104 & ~n8111 ) | ( n8110 & ~n8111 ) ;
  assign n8113 = ( n8091 & ~n8095 ) | ( n8091 & n8112 ) | ( ~n8095 & n8112 ) ;
  assign n8114 = ( n8091 & n8095 ) | ( n8091 & n8112 ) | ( n8095 & n8112 ) ;
  assign n8115 = ( n8095 & n8113 ) | ( n8095 & ~n8114 ) | ( n8113 & ~n8114 ) ;
  assign n8116 = n8085 & n8087 ;
  assign n8117 = n8103 | n8116 ;
  assign n8118 = x59 & x61 ;
  assign n8119 = x58 & x62 ;
  assign n8120 = x57 & x63 ;
  assign n8121 = ( ~n8118 & n8119 ) | ( ~n8118 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8122 = ( n8118 & n8119 ) | ( n8118 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8123 = ( n8118 & n8121 ) | ( n8118 & ~n8122 ) | ( n8121 & ~n8122 ) ;
  assign n8124 = ( n8107 & n8117 ) | ( n8107 & n8123 ) | ( n8117 & n8123 ) ;
  assign n8125 = ( n8107 & ~n8117 ) | ( n8107 & n8123 ) | ( ~n8117 & n8123 ) ;
  assign n8126 = ( n8117 & ~n8124 ) | ( n8117 & n8125 ) | ( ~n8124 & n8125 ) ;
  assign n8127 = ( n8111 & n8114 ) | ( n8111 & n8126 ) | ( n8114 & n8126 ) ;
  assign n8128 = ( n8111 & ~n8114 ) | ( n8111 & n8126 ) | ( ~n8114 & n8126 ) ;
  assign n8129 = ( n8114 & ~n8127 ) | ( n8114 & n8128 ) | ( ~n8127 & n8128 ) ;
  assign n8130 = x58 & x63 ;
  assign n8131 = x61 & x62 ;
  assign n8132 = x59 & n8131 ;
  assign n8133 = ~x61 & x62 ;
  assign n8134 = ( x60 & n8132 ) | ( x60 & ~n8133 ) | ( n8132 & ~n8133 ) ;
  assign n8135 = x59 & x62 ;
  assign n8136 = ( ~x61 & n8106 ) | ( ~x61 & n8135 ) | ( n8106 & n8135 ) ;
  assign n8137 = ( x61 & ~n8134 ) | ( x61 & n8136 ) | ( ~n8134 & n8136 ) ;
  assign n8138 = ( n8122 & ~n8130 ) | ( n8122 & n8137 ) | ( ~n8130 & n8137 ) ;
  assign n8139 = ( n8122 & n8130 ) | ( n8122 & n8137 ) | ( n8130 & n8137 ) ;
  assign n8140 = ( n8130 & n8138 ) | ( n8130 & ~n8139 ) | ( n8138 & ~n8139 ) ;
  assign n8141 = ( n8124 & n8127 ) | ( n8124 & n8140 ) | ( n8127 & n8140 ) ;
  assign n8142 = ( n8124 & ~n8127 ) | ( n8124 & n8140 ) | ( ~n8127 & n8140 ) ;
  assign n8143 = ( n8127 & ~n8141 ) | ( n8127 & n8142 ) | ( ~n8141 & n8142 ) ;
  assign n8144 = x59 & x63 ;
  assign n8145 = x61 | x62 ;
  assign n8146 = x60 & n8145 ;
  assign n8147 = ( n8131 & n8144 ) | ( n8131 & n8146 ) | ( n8144 & n8146 ) ;
  assign n8148 = ( ~n8131 & n8144 ) | ( ~n8131 & n8146 ) | ( n8144 & n8146 ) ;
  assign n8149 = ( n8132 & ~n8147 ) | ( n8132 & n8148 ) | ( ~n8147 & n8148 ) ;
  assign n8150 = ( n8139 & n8141 ) | ( n8139 & ~n8149 ) | ( n8141 & ~n8149 ) ;
  assign n8151 = ( n8139 & n8141 ) | ( n8139 & n8149 ) | ( n8141 & n8149 ) ;
  assign n8152 = ( n8149 & n8150 ) | ( n8149 & ~n8151 ) | ( n8150 & ~n8151 ) ;
  assign n8153 = x60 & x63 ;
  assign n8154 = n8133 & n8153 ;
  assign n8155 = n8133 | n8153 ;
  assign n8156 = ~n8154 & n8155 ;
  assign n8157 = ( n8147 & ~n8151 ) | ( n8147 & n8156 ) | ( ~n8151 & n8156 ) ;
  assign n8158 = ( n8147 & n8151 ) | ( n8147 & n8156 ) | ( n8151 & n8156 ) ;
  assign n8159 = ( n8151 & n8157 ) | ( n8151 & ~n8158 ) | ( n8157 & ~n8158 ) ;
  assign n8160 = x61 & x63 ;
  assign n8161 = ( x63 & n8146 ) | ( x63 & n8160 ) | ( n8146 & n8160 ) ;
  assign n8162 = ( n8131 & ~n8158 ) | ( n8131 & n8161 ) | ( ~n8158 & n8161 ) ;
  assign n8163 = ( n8158 & n8160 ) | ( n8158 & n8161 ) | ( n8160 & n8161 ) ;
  assign n8164 = ( x62 & n8145 ) | ( x62 & n8158 ) | ( n8145 & n8158 ) ;
  assign n8165 = x63 & n8164 ;
  assign n8166 = ( ~n8145 & n8163 ) | ( ~n8145 & n8165 ) | ( n8163 & n8165 ) ;
  assign n8167 = ( n8158 & n8162 ) | ( n8158 & ~n8166 ) | ( n8162 & ~n8166 ) ;
  assign n8168 = ( ~x61 & x63 ) | ( ~x61 & n8162 ) | ( x63 & n8162 ) ;
  assign n8169 = ( ~n8145 & n8163 ) | ( ~n8145 & n8168 ) | ( n8163 & n8168 ) ;
  assign y0 = x0 ;
  assign y1 = 1'b0 ;
  assign y2 = n65 ;
  assign y3 = n68 ;
  assign y4 = n73 ;
  assign y5 = n80 ;
  assign y6 = n88 ;
  assign y7 = n103 ;
  assign y8 = n123 ;
  assign y9 = n141 ;
  assign y10 = n161 ;
  assign y11 = n183 ;
  assign y12 = n209 ;
  assign y13 = n235 ;
  assign y14 = n260 ;
  assign y15 = n291 ;
  assign y16 = n320 ;
  assign y17 = n354 ;
  assign y18 = n389 ;
  assign y19 = n425 ;
  assign y20 = n465 ;
  assign y21 = n506 ;
  assign y22 = n553 ;
  assign y23 = n599 ;
  assign y24 = n647 ;
  assign y25 = n694 ;
  assign y26 = n744 ;
  assign y27 = n799 ;
  assign y28 = n852 ;
  assign y29 = n909 ;
  assign y30 = n969 ;
  assign y31 = n1030 ;
  assign y32 = n1091 ;
  assign y33 = n1157 ;
  assign y34 = n1230 ;
  assign y35 = n1299 ;
  assign y36 = n1371 ;
  assign y37 = n1445 ;
  assign y38 = n1518 ;
  assign y39 = n1597 ;
  assign y40 = n1676 ;
  assign y41 = n1758 ;
  assign y42 = n1845 ;
  assign y43 = n1934 ;
  assign y44 = n2022 ;
  assign y45 = n2111 ;
  assign y46 = n2200 ;
  assign y47 = n2293 ;
  assign y48 = n2389 ;
  assign y49 = n2487 ;
  assign y50 = n2585 ;
  assign y51 = n2688 ;
  assign y52 = n2793 ;
  assign y53 = n2897 ;
  assign y54 = n3005 ;
  assign y55 = n3115 ;
  assign y56 = n3224 ;
  assign y57 = n3339 ;
  assign y58 = n3457 ;
  assign y59 = n3574 ;
  assign y60 = n3694 ;
  assign y61 = n3815 ;
  assign y62 = n3938 ;
  assign y63 = n4063 ;
  assign y64 = n4196 ;
  assign y65 = n4324 ;
  assign y66 = n4451 ;
  assign y67 = n4570 ;
  assign y68 = n4690 ;
  assign y69 = n4806 ;
  assign y70 = n4922 ;
  assign y71 = n5033 ;
  assign y72 = n5145 ;
  assign y73 = n5252 ;
  assign y74 = n5360 ;
  assign y75 = n5464 ;
  assign y76 = n5567 ;
  assign y77 = n5666 ;
  assign y78 = n5766 ;
  assign y79 = n5861 ;
  assign y80 = n5956 ;
  assign y81 = n6048 ;
  assign y82 = n6139 ;
  assign y83 = n6227 ;
  assign y84 = n6315 ;
  assign y85 = n6398 ;
  assign y86 = n6481 ;
  assign y87 = n6561 ;
  assign y88 = n6640 ;
  assign y89 = n6720 ;
  assign y90 = n6797 ;
  assign y91 = n6868 ;
  assign y92 = n6939 ;
  assign y93 = n7007 ;
  assign y94 = n7075 ;
  assign y95 = n7138 ;
  assign y96 = n7201 ;
  assign y97 = n7261 ;
  assign y98 = n7321 ;
  assign y99 = n7377 ;
  assign y100 = n7433 ;
  assign y101 = n7485 ;
  assign y102 = n7537 ;
  assign y103 = n7585 ;
  assign y104 = n7633 ;
  assign y105 = n7677 ;
  assign y106 = n7721 ;
  assign y107 = n7761 ;
  assign y108 = n7800 ;
  assign y109 = n7836 ;
  assign y110 = n7872 ;
  assign y111 = n7904 ;
  assign y112 = n7936 ;
  assign y113 = n7964 ;
  assign y114 = n7992 ;
  assign y115 = n8016 ;
  assign y116 = n8040 ;
  assign y117 = n8060 ;
  assign y118 = n8080 ;
  assign y119 = n8096 ;
  assign y120 = n8115 ;
  assign y121 = n8129 ;
  assign y122 = n8143 ;
  assign y123 = n8152 ;
  assign y124 = n8159 ;
  assign y125 = n8167 ;
  assign y126 = n8169 ;
  assign y127 = n8165 ;
endmodule
