module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 ;
  assign n148 = x3 | x129 ;
  assign n149 = x54 & ~n148 ;
  assign n150 = ~x4 & n149 ;
  assign n151 = ~x17 & n150 ;
  assign n152 = x11 | x22 ;
  assign n153 = x19 | n152 ;
  assign n154 = n151 & ~n153 ;
  assign n155 = x16 | x18 ;
  assign n156 = n154 & ~n155 ;
  assign n157 = x14 | x21 ;
  assign n158 = ( x8 & x10 ) | ( x8 & n157 ) | ( x10 & n157 ) ;
  assign n159 = x14 & x21 ;
  assign n160 = n158 | n159 ;
  assign n161 = x9 | x12 ;
  assign n162 = x5 | x6 ;
  assign n163 = n161 | n162 ;
  assign n164 = x7 | x13 ;
  assign n165 = n163 | n164 ;
  assign n166 = ( x7 & x13 ) | ( x7 & n163 ) | ( x13 & n163 ) ;
  assign n167 = ( n163 & n165 ) | ( n163 & n166 ) | ( n165 & n166 ) ;
  assign n168 = n160 | n167 ;
  assign n169 = x8 | x10 ;
  assign n170 = n157 | n169 ;
  assign n171 = n164 & n170 ;
  assign n172 = n168 | n171 ;
  assign n173 = n156 & ~n172 ;
  assign n174 = x5 | x22 ;
  assign n175 = x9 | x11 ;
  assign n176 = ( x56 & n174 ) | ( x56 & n175 ) | ( n174 & n175 ) ;
  assign n177 = ( n149 & n174 ) | ( n149 & n175 ) | ( n174 & n175 ) ;
  assign n178 = ~n176 & n177 ;
  assign n179 = n173 | n178 ;
  assign n180 = x54 | n148 ;
  assign n181 = x0 | n180 ;
  assign n182 = n165 | n170 ;
  assign n183 = n155 | n182 ;
  assign n184 = n153 | n183 ;
  assign n185 = x0 & ~n184 ;
  assign n186 = ( ~n179 & n181 ) | ( ~n179 & n185 ) | ( n181 & n185 ) ;
  assign n187 = ( x5 & x9 ) | ( x5 & n161 ) | ( x9 & n161 ) ;
  assign n188 = x5 | x12 ;
  assign n189 = ( x6 & n187 ) | ( x6 & n188 ) | ( n187 & n188 ) ;
  assign n190 = n170 | n189 ;
  assign n191 = n166 | n190 ;
  assign n192 = n156 & ~n191 ;
  assign n193 = ( ~x17 & n148 ) | ( ~x17 & n180 ) | ( n148 & n180 ) ;
  assign n194 = x1 | n193 ;
  assign n195 = x1 & ~n165 ;
  assign n196 = ( ~n192 & n194 ) | ( ~n192 & n195 ) | ( n194 & n195 ) ;
  assign n197 = ~x44 & x82 ;
  assign n198 = ~x42 & n197 ;
  assign n199 = ~x40 & n198 ;
  assign n200 = ~x38 & n199 ;
  assign n201 = ~x50 & n200 ;
  assign n202 = ~x46 & n201 ;
  assign n203 = ~x41 & n202 ;
  assign n204 = ~x43 & n203 ;
  assign n205 = ~x47 & n204 ;
  assign n206 = ~x48 & n205 ;
  assign n207 = ~x45 & n206 ;
  assign n208 = ~x24 & n207 ;
  assign n209 = ~x49 & n208 ;
  assign n210 = ~x15 & n209 ;
  assign n211 = x2 | x20 ;
  assign n212 = n210 & ~n211 ;
  assign n213 = x82 & ~n212 ;
  assign n214 = x122 & x127 ;
  assign n215 = n213 | n214 ;
  assign n216 = x65 | n215 ;
  assign n217 = x20 & n210 ;
  assign n218 = ( ~n210 & n215 ) | ( ~n210 & n217 ) | ( n215 & n217 ) ;
  assign n219 = x2 & n218 ;
  assign n220 = ( x129 & n216 ) | ( x129 & ~n219 ) | ( n216 & ~n219 ) ;
  assign n221 = x123 | x129 ;
  assign n222 = x0 & ~x113 ;
  assign n223 = ~n221 & n222 ;
  assign n224 = x4 | x17 ;
  assign n225 = n184 | n224 ;
  assign n226 = x61 | x118 ;
  assign n227 = x129 | n226 ;
  assign n228 = ~n223 & n227 ;
  assign n229 = ( n223 & n225 ) | ( n223 & ~n228 ) | ( n225 & ~n228 ) ;
  assign n230 = x4 & ~n180 ;
  assign n231 = x10 | n230 ;
  assign n232 = ( n173 & n230 ) | ( n173 & n231 ) | ( n230 & n231 ) ;
  assign n233 = n156 & ~n182 ;
  assign n234 = ~x29 & n233 ;
  assign n235 = x5 & ~n180 ;
  assign n236 = x25 | x59 ;
  assign n237 = x28 & ~n236 ;
  assign n238 = n235 | n237 ;
  assign n239 = ( n234 & n235 ) | ( n234 & n238 ) | ( n235 & n238 ) ;
  assign n240 = ~x28 & n234 ;
  assign n241 = x6 & ~n180 ;
  assign n242 = x25 & ~x59 ;
  assign n243 = n241 | n242 ;
  assign n244 = ( n240 & n241 ) | ( n240 & n243 ) | ( n241 & n243 ) ;
  assign n245 = x7 & ~n180 ;
  assign n246 = x8 | n245 ;
  assign n247 = ( n173 & n245 ) | ( n173 & n246 ) | ( n245 & n246 ) ;
  assign n248 = x8 & ~n180 ;
  assign n249 = x21 | n248 ;
  assign n250 = ( n173 & n248 ) | ( n173 & n249 ) | ( n248 & n249 ) ;
  assign n251 = n151 & ~n183 ;
  assign n252 = ~x19 & n251 ;
  assign n253 = x9 & ~n180 ;
  assign n254 = x11 & ~x22 ;
  assign n255 = n253 | n254 ;
  assign n256 = ( n252 & n253 ) | ( n252 & n255 ) | ( n253 & n255 ) ;
  assign n257 = x10 & ~n180 ;
  assign n258 = x14 | n257 ;
  assign n259 = ( n173 & n257 ) | ( n173 & n258 ) | ( n257 & n258 ) ;
  assign n260 = ~x11 & n252 ;
  assign n261 = x11 & ~n180 ;
  assign n262 = ( n152 & n260 ) | ( n152 & n261 ) | ( n260 & n261 ) ;
  assign n263 = n154 & ~n182 ;
  assign n264 = x12 & ~n180 ;
  assign n265 = ( ~x16 & n155 ) | ( ~x16 & n264 ) | ( n155 & n264 ) ;
  assign n266 = ( n263 & n264 ) | ( n263 & n265 ) | ( n264 & n265 ) ;
  assign n267 = x13 & ~n180 ;
  assign n268 = ~x28 & x29 ;
  assign n269 = ~n236 & n268 ;
  assign n270 = n267 | n269 ;
  assign n271 = ( n233 & n267 ) | ( n233 & n270 ) | ( n267 & n270 ) ;
  assign n272 = x14 & ~n180 ;
  assign n273 = x13 | n272 ;
  assign n274 = ( n192 & n272 ) | ( n192 & n273 ) | ( n272 & n273 ) ;
  assign n275 = ( x15 & n209 ) | ( x15 & n212 ) | ( n209 & n212 ) ;
  assign n276 = ( x15 & n210 ) | ( x15 & ~n275 ) | ( n210 & ~n275 ) ;
  assign n277 = n215 & n276 ;
  assign n278 = x70 | n215 ;
  assign n279 = ( x129 & ~n277 ) | ( x129 & n278 ) | ( ~n277 & n278 ) ;
  assign n280 = x16 & ~n180 ;
  assign n281 = x6 | n280 ;
  assign n282 = ( n192 & n280 ) | ( n192 & n281 ) | ( n280 & n281 ) ;
  assign n283 = x17 & ~n180 ;
  assign n284 = ( ~x25 & n236 ) | ( ~x25 & n283 ) | ( n236 & n283 ) ;
  assign n285 = ( n240 & n283 ) | ( n240 & n284 ) | ( n283 & n284 ) ;
  assign n286 = ~x18 & n263 ;
  assign n287 = x18 & ~n180 ;
  assign n288 = ( n155 & n286 ) | ( n155 & n287 ) | ( n286 & n287 ) ;
  assign n289 = x19 & ~n180 ;
  assign n290 = ( n150 & ~n151 ) | ( n150 & n289 ) | ( ~n151 & n289 ) ;
  assign n291 = ( ~n184 & n289 ) | ( ~n184 & n290 ) | ( n289 & n290 ) ;
  assign n292 = x129 | n215 ;
  assign n293 = x71 | n292 ;
  assign n294 = ~x129 & n215 ;
  assign n295 = ~n212 & n294 ;
  assign n296 = ( x20 & n210 ) | ( x20 & n295 ) | ( n210 & n295 ) ;
  assign n297 = ( n217 & n293 ) | ( n217 & ~n296 ) | ( n293 & ~n296 ) ;
  assign n298 = x21 & ~n180 ;
  assign n299 = ( ~n152 & n153 ) | ( ~n152 & n298 ) | ( n153 & n298 ) ;
  assign n300 = ( n251 & n298 ) | ( n251 & n299 ) | ( n298 & n299 ) ;
  assign n301 = x22 & ~n180 ;
  assign n302 = x5 | n301 ;
  assign n303 = ( n192 & n301 ) | ( n192 & n302 ) | ( n301 & n302 ) ;
  assign n304 = ~x23 & x55 ;
  assign n305 = x61 & ~x129 ;
  assign n306 = ~n304 & n305 ;
  assign n307 = x63 | n292 ;
  assign n308 = ( x24 & n207 ) | ( x24 & n295 ) | ( n207 & n295 ) ;
  assign n309 = x24 & n207 ;
  assign n310 = ( n307 & ~n308 ) | ( n307 & n309 ) | ( ~n308 & n309 ) ;
  assign n311 = x116 & ~n148 ;
  assign n312 = x85 & n311 ;
  assign n313 = x53 | x58 ;
  assign n314 = x26 | x27 ;
  assign n315 = x85 | n313 ;
  assign n316 = x53 & x58 ;
  assign n317 = ( x85 & n315 ) | ( x85 & n316 ) | ( n315 & n316 ) ;
  assign n318 = ( n313 & n314 ) | ( n313 & n317 ) | ( n314 & n317 ) ;
  assign n319 = n312 & ~n318 ;
  assign n320 = n314 | n315 ;
  assign n321 = x110 | n148 ;
  assign n322 = n320 | n321 ;
  assign n323 = x96 | n322 ;
  assign n324 = ~n319 & n323 ;
  assign n325 = x26 & x27 ;
  assign n326 = n148 | n325 ;
  assign n327 = n318 | n326 ;
  assign n328 = x51 | x52 ;
  assign n329 = ~x39 & x116 ;
  assign n330 = ~n328 & n329 ;
  assign n331 = x26 & ~n330 ;
  assign n332 = ~n327 & n331 ;
  assign n333 = x100 | n332 ;
  assign n334 = ( ~n324 & n332 ) | ( ~n324 & n333 ) | ( n332 & n333 ) ;
  assign n335 = x95 | x100 ;
  assign n336 = x97 | n335 ;
  assign n337 = ~n322 & n336 ;
  assign n338 = x116 | n327 ;
  assign n339 = ( n320 & n327 ) | ( n320 & n338 ) | ( n327 & n338 ) ;
  assign n340 = n337 | n339 ;
  assign n341 = x27 & n330 ;
  assign n342 = ( n327 & n340 ) | ( n327 & ~n341 ) | ( n340 & ~n341 ) ;
  assign n343 = ~n334 & n342 ;
  assign n344 = x25 | n340 ;
  assign n345 = ~n343 & n344 ;
  assign n346 = x58 & x116 ;
  assign n347 = ~n327 & n346 ;
  assign n348 = n323 | n335 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = x100 | n324 ;
  assign n351 = n349 & ~n350 ;
  assign n352 = x27 & ~n330 ;
  assign n353 = ~n327 & n352 ;
  assign n354 = n351 | n353 ;
  assign n355 = x28 & ~n340 ;
  assign n356 = n318 | n331 ;
  assign n357 = x26 & x116 ;
  assign n358 = ( x116 & n352 ) | ( x116 & n357 ) | ( n352 & n357 ) ;
  assign n359 = ~n326 & n358 ;
  assign n360 = ~n356 & n359 ;
  assign n361 = n355 | n360 ;
  assign n362 = n351 | n361 ;
  assign n363 = x97 & ~n349 ;
  assign n364 = x29 & ~n340 ;
  assign n365 = n363 | n364 ;
  assign n366 = x106 | x129 ;
  assign n367 = x60 & x109 ;
  assign n368 = x30 & ~x109 ;
  assign n369 = ( ~n366 & n367 ) | ( ~n366 & n368 ) | ( n367 & n368 ) ;
  assign n370 = x106 & ~x129 ;
  assign n371 = x88 & n370 ;
  assign n372 = n369 | n371 ;
  assign n373 = x30 & x109 ;
  assign n374 = x31 & ~x109 ;
  assign n375 = ( ~n366 & n373 ) | ( ~n366 & n374 ) | ( n373 & n374 ) ;
  assign n376 = x89 & n370 ;
  assign n377 = n375 | n376 ;
  assign n378 = x31 & x109 ;
  assign n379 = x32 & ~x109 ;
  assign n380 = ( ~n366 & n378 ) | ( ~n366 & n379 ) | ( n378 & n379 ) ;
  assign n381 = x99 & n370 ;
  assign n382 = n380 | n381 ;
  assign n383 = x32 & x109 ;
  assign n384 = x33 & ~x109 ;
  assign n385 = ( ~n366 & n383 ) | ( ~n366 & n384 ) | ( n383 & n384 ) ;
  assign n386 = x90 & n370 ;
  assign n387 = n385 | n386 ;
  assign n388 = x33 & x109 ;
  assign n389 = x34 & ~x109 ;
  assign n390 = ( ~n366 & n388 ) | ( ~n366 & n389 ) | ( n388 & n389 ) ;
  assign n391 = x91 & n370 ;
  assign n392 = n390 | n391 ;
  assign n393 = x34 & x109 ;
  assign n394 = x35 & ~x109 ;
  assign n395 = ( ~n366 & n393 ) | ( ~n366 & n394 ) | ( n393 & n394 ) ;
  assign n396 = x92 & n370 ;
  assign n397 = n395 | n396 ;
  assign n398 = x35 & x109 ;
  assign n399 = x36 & ~x109 ;
  assign n400 = ( ~n366 & n398 ) | ( ~n366 & n399 ) | ( n398 & n399 ) ;
  assign n401 = x98 & n370 ;
  assign n402 = n400 | n401 ;
  assign n403 = x36 & x109 ;
  assign n404 = x37 & ~x109 ;
  assign n405 = ( ~n366 & n403 ) | ( ~n366 & n404 ) | ( n403 & n404 ) ;
  assign n406 = x93 & n370 ;
  assign n407 = n405 | n406 ;
  assign n408 = x74 | n292 ;
  assign n409 = ( x38 & n199 ) | ( x38 & n295 ) | ( n199 & n295 ) ;
  assign n410 = x38 & n199 ;
  assign n411 = ( n408 & ~n409 ) | ( n408 & n410 ) | ( ~n409 & n410 ) ;
  assign n412 = ~x51 & x109 ;
  assign n413 = ~x52 & n412 ;
  assign n414 = ( x39 & x106 ) | ( x39 & ~n413 ) | ( x106 & ~n413 ) ;
  assign n415 = ~x39 & n413 ;
  assign n416 = ( ~x129 & n414 ) | ( ~x129 & n415 ) | ( n414 & n415 ) ;
  assign n417 = x73 | n292 ;
  assign n418 = ( x40 & n198 ) | ( x40 & n295 ) | ( n198 & n295 ) ;
  assign n419 = x40 & n198 ;
  assign n420 = ( n417 & ~n418 ) | ( n417 & n419 ) | ( ~n418 & n419 ) ;
  assign n421 = x76 | n215 ;
  assign n422 = x41 & ~n202 ;
  assign n423 = n203 & n213 ;
  assign n424 = ( n215 & n422 ) | ( n215 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ( x129 & n421 ) | ( x129 & ~n424 ) | ( n421 & ~n424 ) ;
  assign n426 = x72 | n292 ;
  assign n427 = ( x42 & n197 ) | ( x42 & n295 ) | ( n197 & n295 ) ;
  assign n428 = x42 & n197 ;
  assign n429 = ( n426 & ~n427 ) | ( n426 & n428 ) | ( ~n427 & n428 ) ;
  assign n430 = x77 | n292 ;
  assign n431 = ( x43 & n203 ) | ( x43 & n295 ) | ( n203 & n295 ) ;
  assign n432 = x43 & n203 ;
  assign n433 = ( n430 & ~n431 ) | ( n430 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = x67 | n292 ;
  assign n435 = ( x44 & n213 ) | ( x44 & n294 ) | ( n213 & n294 ) ;
  assign n436 = x44 & n213 ;
  assign n437 = ( n434 & ~n435 ) | ( n434 & n436 ) | ( ~n435 & n436 ) ;
  assign n438 = x68 | n292 ;
  assign n439 = ( x45 & n206 ) | ( x45 & n295 ) | ( n206 & n295 ) ;
  assign n440 = x45 & n206 ;
  assign n441 = ( n438 & ~n439 ) | ( n438 & n440 ) | ( ~n439 & n440 ) ;
  assign n442 = x75 | n292 ;
  assign n443 = ( x46 & n201 ) | ( x46 & n295 ) | ( n201 & n295 ) ;
  assign n444 = x46 & n201 ;
  assign n445 = ( n442 & ~n443 ) | ( n442 & n444 ) | ( ~n443 & n444 ) ;
  assign n446 = x64 | n292 ;
  assign n447 = ( x47 & n204 ) | ( x47 & n295 ) | ( n204 & n295 ) ;
  assign n448 = x47 & n204 ;
  assign n449 = ( n446 & ~n447 ) | ( n446 & n448 ) | ( ~n447 & n448 ) ;
  assign n450 = x62 | n292 ;
  assign n451 = ( x48 & n205 ) | ( x48 & n295 ) | ( n205 & n295 ) ;
  assign n452 = x48 & n205 ;
  assign n453 = ( n450 & ~n451 ) | ( n450 & n452 ) | ( ~n451 & n452 ) ;
  assign n454 = x69 | n292 ;
  assign n455 = ( x49 & n208 ) | ( x49 & n295 ) | ( n208 & n295 ) ;
  assign n456 = x49 & n208 ;
  assign n457 = ( n454 & ~n455 ) | ( n454 & n456 ) | ( ~n455 & n456 ) ;
  assign n458 = x66 | n292 ;
  assign n459 = ( x50 & n200 ) | ( x50 & n295 ) | ( n200 & n295 ) ;
  assign n460 = x50 & n200 ;
  assign n461 = ( n458 & ~n459 ) | ( n458 & n460 ) | ( ~n459 & n460 ) ;
  assign n462 = ( x51 & x106 ) | ( x51 & ~x109 ) | ( x106 & ~x109 ) ;
  assign n463 = ( ~x129 & n412 ) | ( ~x129 & n462 ) | ( n412 & n462 ) ;
  assign n464 = ( x52 & x106 ) | ( x52 & ~n412 ) | ( x106 & ~n412 ) ;
  assign n465 = ( ~x129 & n413 ) | ( ~x129 & n464 ) | ( n413 & n464 ) ;
  assign n466 = x53 & ~n338 ;
  assign n467 = n363 | n466 ;
  assign n468 = x114 & ~x122 ;
  assign n469 = ~n221 & n468 ;
  assign n470 = x58 | n357 ;
  assign n471 = ~x94 & n470 ;
  assign n472 = x37 | n470 ;
  assign n473 = ( n346 & ~n471 ) | ( n346 & n472 ) | ( ~n471 & n472 ) ;
  assign n474 = ~n327 & n473 ;
  assign n475 = x57 & ~n346 ;
  assign n476 = x60 & n346 ;
  assign n477 = ( ~n327 & n475 ) | ( ~n327 & n476 ) | ( n475 & n476 ) ;
  assign n478 = x58 | n330 ;
  assign n479 = x116 & ~n314 ;
  assign n480 = n478 & ~n479 ;
  assign n481 = ~n327 & n480 ;
  assign n482 = x59 & ~n340 ;
  assign n483 = x96 & n337 ;
  assign n484 = n482 | n483 ;
  assign n485 = ~x60 & x122 ;
  assign n486 = ( x60 & x117 ) | ( x60 & x122 ) | ( x117 & x122 ) ;
  assign n487 = ~x117 & x123 ;
  assign n488 = ( ~n485 & n486 ) | ( ~n485 & n487 ) | ( n486 & n487 ) ;
  assign n489 = x114 | x122 ;
  assign n490 = x123 & ~x129 ;
  assign n491 = ~n489 & n490 ;
  assign n492 = x136 & ~x137 ;
  assign n493 = ~x138 & n492 ;
  assign n494 = x132 & x133 ;
  assign n495 = x131 & n494 ;
  assign n496 = n493 & n495 ;
  assign n497 = x62 & ~n496 ;
  assign n498 = ~x140 & n496 ;
  assign n499 = ( ~x129 & n497 ) | ( ~x129 & n498 ) | ( n497 & n498 ) ;
  assign n500 = x63 & ~n496 ;
  assign n501 = ~x142 & n496 ;
  assign n502 = ( ~x129 & n500 ) | ( ~x129 & n501 ) | ( n500 & n501 ) ;
  assign n503 = x64 & ~n496 ;
  assign n504 = ~x139 & n496 ;
  assign n505 = ( ~x129 & n503 ) | ( ~x129 & n504 ) | ( n503 & n504 ) ;
  assign n506 = x65 & ~n496 ;
  assign n507 = ~x146 & n496 ;
  assign n508 = ( ~x129 & n506 ) | ( ~x129 & n507 ) | ( n506 & n507 ) ;
  assign n509 = x136 | x137 ;
  assign n510 = x138 | n509 ;
  assign n511 = n495 & ~n510 ;
  assign n512 = x66 & ~n511 ;
  assign n513 = ~x143 & n511 ;
  assign n514 = ( ~x129 & n512 ) | ( ~x129 & n513 ) | ( n512 & n513 ) ;
  assign n515 = x67 & ~n511 ;
  assign n516 = ~x139 & n511 ;
  assign n517 = ( ~x129 & n515 ) | ( ~x129 & n516 ) | ( n515 & n516 ) ;
  assign n518 = x68 & ~n496 ;
  assign n519 = ~x141 & n496 ;
  assign n520 = ( ~x129 & n518 ) | ( ~x129 & n519 ) | ( n518 & n519 ) ;
  assign n521 = x69 & ~n496 ;
  assign n522 = ~x143 & n496 ;
  assign n523 = ( ~x129 & n521 ) | ( ~x129 & n522 ) | ( n521 & n522 ) ;
  assign n524 = x70 & ~n496 ;
  assign n525 = ~x144 & n496 ;
  assign n526 = ( ~x129 & n524 ) | ( ~x129 & n525 ) | ( n524 & n525 ) ;
  assign n527 = x71 & ~n496 ;
  assign n528 = ~x145 & n496 ;
  assign n529 = ( ~x129 & n527 ) | ( ~x129 & n528 ) | ( n527 & n528 ) ;
  assign n530 = x72 & ~n511 ;
  assign n531 = ~x140 & n511 ;
  assign n532 = ( ~x129 & n530 ) | ( ~x129 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x73 & ~n511 ;
  assign n534 = ~x141 & n511 ;
  assign n535 = ( ~x129 & n533 ) | ( ~x129 & n534 ) | ( n533 & n534 ) ;
  assign n536 = x74 & ~n511 ;
  assign n537 = ~x142 & n511 ;
  assign n538 = ( ~x129 & n536 ) | ( ~x129 & n537 ) | ( n536 & n537 ) ;
  assign n539 = x75 & ~n511 ;
  assign n540 = ~x144 & n511 ;
  assign n541 = ( ~x129 & n539 ) | ( ~x129 & n540 ) | ( n539 & n540 ) ;
  assign n542 = x76 & ~n511 ;
  assign n543 = ~x145 & n511 ;
  assign n544 = ( ~x129 & n542 ) | ( ~x129 & n543 ) | ( n542 & n543 ) ;
  assign n545 = x77 & ~n511 ;
  assign n546 = ~x146 & n511 ;
  assign n547 = ( ~x129 & n545 ) | ( ~x129 & n546 ) | ( n545 & n546 ) ;
  assign n548 = ~x136 & x137 ;
  assign n549 = ~x138 & n548 ;
  assign n550 = n495 & n549 ;
  assign n551 = x78 & ~n550 ;
  assign n552 = x142 & n550 ;
  assign n553 = ( ~x129 & n551 ) | ( ~x129 & n552 ) | ( n551 & n552 ) ;
  assign n554 = x79 & ~n550 ;
  assign n555 = x143 & n550 ;
  assign n556 = ( ~x129 & n554 ) | ( ~x129 & n555 ) | ( n554 & n555 ) ;
  assign n557 = x80 & ~n550 ;
  assign n558 = x144 & n550 ;
  assign n559 = ( ~x129 & n557 ) | ( ~x129 & n558 ) | ( n557 & n558 ) ;
  assign n560 = x81 & ~n550 ;
  assign n561 = x145 & n550 ;
  assign n562 = ( ~x129 & n560 ) | ( ~x129 & n561 ) | ( n560 & n561 ) ;
  assign n563 = x82 & ~n550 ;
  assign n564 = x146 & n550 ;
  assign n565 = ( ~x129 & n563 ) | ( ~x129 & n564 ) | ( n563 & n564 ) ;
  assign n566 = ~x62 & n493 ;
  assign n567 = x138 & ~n509 ;
  assign n568 = x119 & n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = x138 & n548 ;
  assign n571 = ~x115 & n570 ;
  assign n572 = n569 | n571 ;
  assign n573 = x136 & x137 ;
  assign n574 = ~x138 & n573 ;
  assign n575 = x31 & n574 ;
  assign n576 = x72 | n510 ;
  assign n577 = ~n575 & n576 ;
  assign n578 = x138 & n492 ;
  assign n579 = x89 & n578 ;
  assign n580 = x87 & n549 ;
  assign n581 = n579 | n580 ;
  assign n582 = n577 & ~n581 ;
  assign n583 = ~n572 & n582 ;
  assign n584 = x84 & ~n550 ;
  assign n585 = x141 & n550 ;
  assign n586 = ( ~x129 & n584 ) | ( ~x129 & n585 ) | ( n584 & n585 ) ;
  assign n587 = x85 & ~n338 ;
  assign n588 = n483 | n587 ;
  assign n589 = x86 & ~n550 ;
  assign n590 = x139 & n550 ;
  assign n591 = ( ~x129 & n589 ) | ( ~x129 & n590 ) | ( n589 & n590 ) ;
  assign n592 = x87 & ~n550 ;
  assign n593 = x140 & n550 ;
  assign n594 = ( ~x129 & n592 ) | ( ~x129 & n593 ) | ( n592 & n593 ) ;
  assign n595 = n495 & n574 ;
  assign n596 = x88 & ~n595 ;
  assign n597 = x139 & n595 ;
  assign n598 = ( ~x129 & n596 ) | ( ~x129 & n597 ) | ( n596 & n597 ) ;
  assign n599 = x89 & ~n595 ;
  assign n600 = x140 & n595 ;
  assign n601 = ( ~x129 & n599 ) | ( ~x129 & n600 ) | ( n599 & n600 ) ;
  assign n602 = x90 & ~n595 ;
  assign n603 = x142 & n595 ;
  assign n604 = ( ~x129 & n602 ) | ( ~x129 & n603 ) | ( n602 & n603 ) ;
  assign n605 = x91 & ~n595 ;
  assign n606 = x143 & n595 ;
  assign n607 = ( ~x129 & n605 ) | ( ~x129 & n606 ) | ( n605 & n606 ) ;
  assign n608 = x92 & ~n595 ;
  assign n609 = x144 & n595 ;
  assign n610 = ( ~x129 & n608 ) | ( ~x129 & n609 ) | ( n608 & n609 ) ;
  assign n611 = x93 & ~n595 ;
  assign n612 = x146 & n595 ;
  assign n613 = ( ~x129 & n611 ) | ( ~x129 & n612 ) | ( n611 & n612 ) ;
  assign n614 = x82 & n567 ;
  assign n615 = n495 & n614 ;
  assign n616 = x94 & ~n615 ;
  assign n617 = x142 & n615 ;
  assign n618 = ( ~x129 & n616 ) | ( ~x129 & n617 ) | ( n616 & n617 ) ;
  assign n619 = ~x129 & n495 ;
  assign n620 = n321 & ~n619 ;
  assign n621 = x95 & ~n615 ;
  assign n622 = x143 & n615 ;
  assign n623 = ( ~n620 & n621 ) | ( ~n620 & n622 ) | ( n621 & n622 ) ;
  assign n624 = x96 & ~n615 ;
  assign n625 = x146 & n615 ;
  assign n626 = ( ~n620 & n624 ) | ( ~n620 & n625 ) | ( n624 & n625 ) ;
  assign n627 = x97 & ~n615 ;
  assign n628 = x145 & n615 ;
  assign n629 = ( ~n620 & n627 ) | ( ~n620 & n628 ) | ( n627 & n628 ) ;
  assign n630 = x98 & ~n595 ;
  assign n631 = x145 & n595 ;
  assign n632 = ( ~x129 & n630 ) | ( ~x129 & n631 ) | ( n630 & n631 ) ;
  assign n633 = x99 & ~n595 ;
  assign n634 = x141 & n595 ;
  assign n635 = ( ~x129 & n633 ) | ( ~x129 & n634 ) | ( n633 & n634 ) ;
  assign n636 = x100 & ~n615 ;
  assign n637 = x144 & n615 ;
  assign n638 = ( ~n620 & n636 ) | ( ~n620 & n637 ) | ( n636 & n637 ) ;
  assign n639 = x93 & n492 ;
  assign n640 = x96 & n548 ;
  assign n641 = n639 | n640 ;
  assign n642 = ( x124 & ~x137 ) | ( x124 & n492 ) | ( ~x137 & n492 ) ;
  assign n643 = ( ~x37 & x136 ) | ( ~x37 & n492 ) | ( x136 & n492 ) ;
  assign n644 = ( x138 & ~n642 ) | ( x138 & n643 ) | ( ~n642 & n643 ) ;
  assign n645 = ~n641 & n644 ;
  assign n646 = x77 & ~n510 ;
  assign n647 = ~x82 & n549 ;
  assign n648 = n646 | n647 ;
  assign n649 = x65 & n493 ;
  assign n650 = n648 | n649 ;
  assign n651 = n645 | n650 ;
  assign n652 = x69 & n493 ;
  assign n653 = ~x34 & n573 ;
  assign n654 = n652 | n653 ;
  assign n655 = ( ~x91 & x136 ) | ( ~x91 & n573 ) | ( x136 & n573 ) ;
  assign n656 = ( x95 & x136 ) | ( x95 & n509 ) | ( x136 & n509 ) ;
  assign n657 = ( x138 & n655 ) | ( x138 & ~n656 ) | ( n655 & ~n656 ) ;
  assign n658 = n654 | n657 ;
  assign n659 = ~x79 & n549 ;
  assign n660 = x66 & ~n509 ;
  assign n661 = n659 | n660 ;
  assign n662 = n658 | n661 ;
  assign n663 = x63 | x137 ;
  assign n664 = x33 & x137 ;
  assign n665 = ( x136 & ~n663 ) | ( x136 & n664 ) | ( ~n663 & n664 ) ;
  assign n666 = x74 | x137 ;
  assign n667 = x78 & x137 ;
  assign n668 = ( x136 & n666 ) | ( x136 & ~n667 ) | ( n666 & ~n667 ) ;
  assign n669 = ~n665 & n668 ;
  assign n670 = x138 | n669 ;
  assign n671 = x94 & n570 ;
  assign n672 = x90 & n578 ;
  assign n673 = n671 | n672 ;
  assign n674 = n670 & ~n673 ;
  assign n675 = x73 | x136 ;
  assign n676 = ~x68 & x136 ;
  assign n677 = ( x137 & n675 ) | ( x137 & ~n676 ) | ( n675 & ~n676 ) ;
  assign n678 = ( x84 & x136 ) | ( x84 & n509 ) | ( x136 & n509 ) ;
  assign n679 = ( ~x32 & x136 ) | ( ~x32 & n492 ) | ( x136 & n492 ) ;
  assign n680 = ( x138 & n678 ) | ( x138 & ~n679 ) | ( n678 & ~n679 ) ;
  assign n681 = n677 & ~n680 ;
  assign n682 = ( ~x99 & x136 ) | ( ~x99 & n573 ) | ( x136 & n573 ) ;
  assign n683 = ( ~x112 & x136 ) | ( ~x112 & n509 ) | ( x136 & n509 ) ;
  assign n684 = ( x138 & n682 ) | ( x138 & ~n683 ) | ( n682 & ~n683 ) ;
  assign n685 = n681 | n684 ;
  assign n686 = x125 & ~x137 ;
  assign n687 = x100 & x137 ;
  assign n688 = ( ~x136 & n686 ) | ( ~x136 & n687 ) | ( n686 & n687 ) ;
  assign n689 = x92 & n492 ;
  assign n690 = n688 | n689 ;
  assign n691 = x35 & ~x138 ;
  assign n692 = ( x138 & n573 ) | ( x138 & ~n691 ) | ( n573 & ~n691 ) ;
  assign n693 = ~n690 & n692 ;
  assign n694 = ~x80 & n549 ;
  assign n695 = x75 & ~n510 ;
  assign n696 = n694 | n695 ;
  assign n697 = x70 & n493 ;
  assign n698 = n696 | n697 ;
  assign n699 = n693 | n698 ;
  assign n700 = n312 | n337 ;
  assign n701 = x81 & n549 ;
  assign n702 = x36 & n574 ;
  assign n703 = n701 | n702 ;
  assign n704 = x23 & n567 ;
  assign n705 = n703 | n704 ;
  assign n706 = x98 & n578 ;
  assign n707 = x97 & n570 ;
  assign n708 = n706 | n707 ;
  assign n709 = ~x71 & n493 ;
  assign n710 = x76 | n510 ;
  assign n711 = ~n709 & n710 ;
  assign n712 = ~n708 & n711 ;
  assign n713 = ~n705 & n712 ;
  assign n714 = x120 & ~x136 ;
  assign n715 = x88 & x136 ;
  assign n716 = ( ~x137 & n714 ) | ( ~x137 & n715 ) | ( n714 & n715 ) ;
  assign n717 = x111 & n548 ;
  assign n718 = n716 | n717 ;
  assign n719 = x30 & ~x138 ;
  assign n720 = ( x138 & n573 ) | ( x138 & ~n719 ) | ( n573 & ~n719 ) ;
  assign n721 = ~n718 & n720 ;
  assign n722 = ~x86 & n549 ;
  assign n723 = x67 & ~n510 ;
  assign n724 = n722 | n723 ;
  assign n725 = x64 & n493 ;
  assign n726 = n724 | n725 ;
  assign n727 = n721 | n726 ;
  assign n728 = ( x53 & x58 ) | ( x53 & n311 ) | ( x58 & n311 ) ;
  assign n729 = ( x58 & x97 ) | ( x58 & n316 ) | ( x97 & n316 ) ;
  assign n730 = n728 & ~n729 ;
  assign n731 = x139 & n614 ;
  assign n732 = x111 & ~n614 ;
  assign n733 = ( n619 & n731 ) | ( n619 & n732 ) | ( n731 & n732 ) ;
  assign n734 = x141 & n614 ;
  assign n735 = x112 | n614 ;
  assign n736 = ( n619 & n734 ) | ( n619 & ~n735 ) | ( n734 & ~n735 ) ;
  assign n737 = x54 & n152 ;
  assign n738 = x54 | x113 ;
  assign n739 = ( n148 & ~n737 ) | ( n148 & n738 ) | ( ~n737 & n738 ) ;
  assign n740 = x140 & n614 ;
  assign n741 = x115 | n614 ;
  assign n742 = ( n619 & n740 ) | ( n619 & ~n741 ) | ( n740 & ~n741 ) ;
  assign n743 = x4 | x7 ;
  assign n744 = n161 | n743 ;
  assign n745 = n149 & n744 ;
  assign n746 = x122 & ~x129 ;
  assign n747 = ~x54 & x118 ;
  assign n748 = x54 & n269 ;
  assign n749 = ( ~x129 & n747 ) | ( ~x129 & n748 ) | ( n747 & n748 ) ;
  assign n750 = ~x129 & n335 ;
  assign n751 = x3 & ~x111 ;
  assign n752 = x110 | x120 ;
  assign n753 = ( ~x111 & n751 ) | ( ~x111 & n752 ) | ( n751 & n752 ) ;
  assign n754 = ~x129 & n753 ;
  assign n755 = x81 & x120 ;
  assign n756 = ~x129 & n755 ;
  assign n757 = x129 | x134 ;
  assign n758 = x129 | x135 ;
  assign n759 = x57 & ~x129 ;
  assign n760 = ~x96 & x125 ;
  assign n761 = x3 & ~x129 ;
  assign n762 = ( ~x129 & n760 ) | ( ~x129 & n761 ) | ( n760 & n761 ) ;
  assign n763 = ~x126 & n494 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = n186 ;
  assign y16 = n196 ;
  assign y17 = ~n220 ;
  assign y18 = n229 ;
  assign y19 = n232 ;
  assign y20 = n239 ;
  assign y21 = n244 ;
  assign y22 = n247 ;
  assign y23 = n250 ;
  assign y24 = n256 ;
  assign y25 = n259 ;
  assign y26 = n262 ;
  assign y27 = n266 ;
  assign y28 = n271 ;
  assign y29 = n274 ;
  assign y30 = ~n279 ;
  assign y31 = n282 ;
  assign y32 = n285 ;
  assign y33 = n288 ;
  assign y34 = n291 ;
  assign y35 = ~n297 ;
  assign y36 = n300 ;
  assign y37 = n303 ;
  assign y38 = n306 ;
  assign y39 = ~n310 ;
  assign y40 = n345 ;
  assign y41 = n334 ;
  assign y42 = n354 ;
  assign y43 = n362 ;
  assign y44 = n365 ;
  assign y45 = n372 ;
  assign y46 = n377 ;
  assign y47 = n382 ;
  assign y48 = n387 ;
  assign y49 = n392 ;
  assign y50 = n397 ;
  assign y51 = n402 ;
  assign y52 = n407 ;
  assign y53 = ~n411 ;
  assign y54 = n416 ;
  assign y55 = ~n420 ;
  assign y56 = ~n425 ;
  assign y57 = ~n429 ;
  assign y58 = ~n433 ;
  assign y59 = ~n437 ;
  assign y60 = ~n441 ;
  assign y61 = ~n445 ;
  assign y62 = ~n449 ;
  assign y63 = ~n453 ;
  assign y64 = ~n457 ;
  assign y65 = ~n461 ;
  assign y66 = n463 ;
  assign y67 = n465 ;
  assign y68 = n467 ;
  assign y69 = ~n294 ;
  assign y70 = n469 ;
  assign y71 = n474 ;
  assign y72 = n477 ;
  assign y73 = n481 ;
  assign y74 = n484 ;
  assign y75 = n488 ;
  assign y76 = n491 ;
  assign y77 = ~n499 ;
  assign y78 = ~n502 ;
  assign y79 = ~n505 ;
  assign y80 = ~n508 ;
  assign y81 = ~n514 ;
  assign y82 = ~n517 ;
  assign y83 = ~n520 ;
  assign y84 = ~n523 ;
  assign y85 = ~n526 ;
  assign y86 = ~n529 ;
  assign y87 = ~n532 ;
  assign y88 = ~n535 ;
  assign y89 = ~n538 ;
  assign y90 = ~n541 ;
  assign y91 = ~n544 ;
  assign y92 = ~n547 ;
  assign y93 = n553 ;
  assign y94 = n556 ;
  assign y95 = n559 ;
  assign y96 = n562 ;
  assign y97 = n565 ;
  assign y98 = ~n583 ;
  assign y99 = n586 ;
  assign y100 = n588 ;
  assign y101 = n591 ;
  assign y102 = n594 ;
  assign y103 = n598 ;
  assign y104 = n601 ;
  assign y105 = n604 ;
  assign y106 = n607 ;
  assign y107 = n610 ;
  assign y108 = n613 ;
  assign y109 = n618 ;
  assign y110 = n623 ;
  assign y111 = n626 ;
  assign y112 = n629 ;
  assign y113 = n632 ;
  assign y114 = n635 ;
  assign y115 = n638 ;
  assign y116 = ~n651 ;
  assign y117 = ~n662 ;
  assign y118 = ~n674 ;
  assign y119 = ~n685 ;
  assign y120 = ~n699 ;
  assign y121 = n700 ;
  assign y122 = ~n713 ;
  assign y123 = ~n727 ;
  assign y124 = n359 ;
  assign y125 = n730 ;
  assign y126 = n733 ;
  assign y127 = n736 ;
  assign y128 = ~n739 ;
  assign y129 = n221 ;
  assign y130 = n742 ;
  assign y131 = n745 ;
  assign y132 = ~n746 ;
  assign y133 = n749 ;
  assign y134 = n750 ;
  assign y135 = n754 ;
  assign y136 = n756 ;
  assign y137 = n757 ;
  assign y138 = n758 ;
  assign y139 = n759 ;
  assign y140 = n762 ;
  assign y141 = n763 ;
endmodule
