module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 ;
  assign n33 = x2 & ~x3 ;
  assign n34 = x2 & x3 ;
  assign n35 = x3 & ~n34 ;
  assign n36 = n33 | n35 ;
  assign n37 = x4 & x5 ;
  assign n38 = x4 | x5 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n36 & ~n39 ;
  assign n41 = ~x0 & x1 ;
  assign n42 = ~x29 & x30 ;
  assign n43 = x27 | x28 ;
  assign n44 = n42 & ~n43 ;
  assign n45 = x25 | x26 ;
  assign n46 = x23 & ~n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = ~x24 & n47 ;
  assign n49 = x29 & x30 ;
  assign n50 = x27 & ~x28 ;
  assign n51 = n49 & n50 ;
  assign n52 = x25 & ~x26 ;
  assign n53 = x23 & ~x24 ;
  assign n54 = n52 & n53 ;
  assign n55 = n51 & n54 ;
  assign n56 = ~x27 & x28 ;
  assign n57 = x29 & ~x30 ;
  assign n58 = n56 & n57 ;
  assign n59 = x23 & x24 ;
  assign n60 = ~x25 & x26 ;
  assign n61 = n59 & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 | n62 ;
  assign n64 = n48 | n63 ;
  assign n65 = x27 & x28 ;
  assign n66 = x29 | x30 ;
  assign n67 = n65 & ~n66 ;
  assign n68 = ~x23 & x24 ;
  assign n69 = ~n45 & n68 ;
  assign n70 = n67 & n69 ;
  assign n71 = n50 & n57 ;
  assign n72 = x23 | x24 ;
  assign n73 = n45 | n72 ;
  assign n74 = n71 & ~n73 ;
  assign n75 = n70 | n74 ;
  assign n76 = n64 | n75 ;
  assign n77 = x25 & x26 ;
  assign n78 = n53 & n77 ;
  assign n79 = n42 & n56 ;
  assign n80 = n78 & n79 ;
  assign n81 = n68 & n77 ;
  assign n82 = n44 & n81 ;
  assign n83 = n80 | n82 ;
  assign n84 = x23 & n52 ;
  assign n85 = n43 | n66 ;
  assign n86 = n84 & ~n85 ;
  assign n87 = x24 & n86 ;
  assign n88 = ~n43 & n57 ;
  assign n89 = n84 & n88 ;
  assign n90 = ~x24 & n89 ;
  assign n91 = n87 | n90 ;
  assign n92 = n83 | n91 ;
  assign n93 = n76 | n92 ;
  assign n94 = n56 & ~n66 ;
  assign n95 = ~x23 & n52 ;
  assign n96 = n94 & n95 ;
  assign n97 = x24 & n96 ;
  assign n98 = ~n43 & n49 ;
  assign n99 = ~n73 & n98 ;
  assign n100 = n97 | n99 ;
  assign n101 = n52 & n59 ;
  assign n102 = n49 & n56 ;
  assign n103 = n101 & n102 ;
  assign n104 = n51 & n69 ;
  assign n105 = n103 | n104 ;
  assign n106 = n100 | n105 ;
  assign n107 = n53 & n60 ;
  assign n108 = n79 & n107 ;
  assign n109 = n52 & ~n72 ;
  assign n110 = n44 & n109 ;
  assign n111 = n108 | n110 ;
  assign n112 = n42 & n50 ;
  assign n113 = n69 & n112 ;
  assign n114 = x23 & n77 ;
  assign n115 = n112 & n114 ;
  assign n116 = n113 | n115 ;
  assign n117 = n111 | n116 ;
  assign n118 = n106 | n117 ;
  assign n119 = n93 | n118 ;
  assign n120 = x25 & n53 ;
  assign n121 = n57 & n65 ;
  assign n122 = n120 & n121 ;
  assign n123 = ~x26 & n122 ;
  assign n124 = n71 & n107 ;
  assign n125 = ~n73 & n94 ;
  assign n126 = n124 | n125 ;
  assign n127 = n123 | n126 ;
  assign n128 = ~n45 & n59 ;
  assign n129 = n98 & n128 ;
  assign n130 = n49 & n65 ;
  assign n131 = n69 & n130 ;
  assign n132 = n129 | n131 ;
  assign n133 = n107 & n112 ;
  assign n134 = n61 & n79 ;
  assign n135 = n133 | n134 ;
  assign n136 = n132 | n135 ;
  assign n137 = n127 | n136 ;
  assign n138 = n119 | n137 ;
  assign n139 = n59 & n77 ;
  assign n140 = n79 & n139 ;
  assign n141 = n61 & n88 ;
  assign n142 = n50 & ~n66 ;
  assign n143 = n60 & n68 ;
  assign n144 = n142 & n143 ;
  assign n145 = n141 | n144 ;
  assign n146 = n140 | n145 ;
  assign n147 = n54 & ~n85 ;
  assign n148 = n78 & n98 ;
  assign n149 = n147 | n148 ;
  assign n150 = n81 & n88 ;
  assign n151 = n61 & n112 ;
  assign n152 = n150 | n151 ;
  assign n153 = n88 & n143 ;
  assign n154 = n152 | n153 ;
  assign n155 = n149 | n154 ;
  assign n156 = n146 | n155 ;
  assign n157 = n52 & n68 ;
  assign n158 = ~x29 & n65 ;
  assign n159 = n157 & n158 ;
  assign n160 = x30 & n159 ;
  assign n161 = n54 & n130 ;
  assign n162 = n160 | n161 ;
  assign n163 = ~n73 & n112 ;
  assign n164 = n61 & n102 ;
  assign n165 = n44 & n101 ;
  assign n166 = n164 | n165 ;
  assign n167 = n163 | n166 ;
  assign n168 = n162 | n167 ;
  assign n169 = n156 | n168 ;
  assign n170 = n138 | n169 ;
  assign n171 = ~x23 & n77 ;
  assign n172 = n102 & n171 ;
  assign n173 = x24 & n172 ;
  assign n174 = n51 & n61 ;
  assign n175 = ~n72 & n77 ;
  assign n176 = n142 & n175 ;
  assign n177 = n174 | n176 ;
  assign n178 = n88 & n157 ;
  assign n179 = n94 & n109 ;
  assign n180 = n178 | n179 ;
  assign n181 = n177 | n180 ;
  assign n182 = n173 | n181 ;
  assign n183 = ~n45 & n53 ;
  assign n184 = n79 & n183 ;
  assign n185 = n71 & n175 ;
  assign n186 = n184 | n185 ;
  assign n187 = n60 & ~n72 ;
  assign n188 = n98 & n187 ;
  assign n189 = n51 & n157 ;
  assign n190 = n188 | n189 ;
  assign n191 = n94 & n107 ;
  assign n192 = n102 & n109 ;
  assign n193 = n191 | n192 ;
  assign n194 = n190 | n193 ;
  assign n195 = n186 | n194 ;
  assign n196 = n182 | n195 ;
  assign n197 = n121 & n139 ;
  assign n198 = n98 & n139 ;
  assign n199 = n197 | n198 ;
  assign n200 = n58 & n81 ;
  assign n201 = ~n73 & n142 ;
  assign n202 = n200 | n201 ;
  assign n203 = n199 | n202 ;
  assign n204 = n196 | n203 ;
  assign n205 = n114 & n130 ;
  assign n206 = x24 & n205 ;
  assign n207 = n51 & n187 ;
  assign n208 = n44 & n157 ;
  assign n209 = n207 | n208 ;
  assign n210 = n69 & n121 ;
  assign n211 = n209 | n210 ;
  assign n212 = n206 | n211 ;
  assign n213 = n204 | n212 ;
  assign n214 = n61 & n94 ;
  assign n215 = n61 & n130 ;
  assign n216 = n214 | n215 ;
  assign n217 = ~n72 & n94 ;
  assign n218 = n60 & n217 ;
  assign n219 = n216 | n218 ;
  assign n220 = n67 & n78 ;
  assign n221 = n107 & n130 ;
  assign n222 = n88 & n107 ;
  assign n223 = n221 | n222 ;
  assign n224 = n220 | n223 ;
  assign n225 = n121 & n187 ;
  assign n226 = ~n85 & n139 ;
  assign n227 = n225 | n226 ;
  assign n228 = n224 | n227 ;
  assign n229 = n219 | n228 ;
  assign n230 = x23 & n121 ;
  assign n231 = x24 & n60 ;
  assign n232 = n230 & n231 ;
  assign n233 = n58 & n157 ;
  assign n234 = n232 | n233 ;
  assign n235 = n42 & n65 ;
  assign n236 = ~x24 & n235 ;
  assign n237 = n95 & n236 ;
  assign n238 = n51 & n81 ;
  assign n239 = n237 | n238 ;
  assign n240 = n234 | n239 ;
  assign n241 = ~n85 & n187 ;
  assign n242 = n54 & n102 ;
  assign n243 = n241 | n242 ;
  assign n244 = n88 & n175 ;
  assign n245 = n69 & n235 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = n240 | n247 ;
  assign n249 = n229 | n248 ;
  assign n250 = n213 | n249 ;
  assign n251 = x24 & n77 ;
  assign n252 = n58 & n251 ;
  assign n253 = x23 & n252 ;
  assign n254 = n101 & n142 ;
  assign n255 = n253 | n254 ;
  assign n256 = n58 & ~n73 ;
  assign n257 = n121 & n171 ;
  assign n258 = n256 | n257 ;
  assign n259 = n255 | n258 ;
  assign n260 = n54 & n79 ;
  assign n261 = n121 & n157 ;
  assign n262 = n260 | n261 ;
  assign n263 = x25 & n59 ;
  assign n264 = n88 & n263 ;
  assign n265 = n128 & n142 ;
  assign n266 = n264 | n265 ;
  assign n267 = n262 | n266 ;
  assign n268 = n71 & n143 ;
  assign n269 = n88 & n128 ;
  assign n270 = ~n73 & n235 ;
  assign n271 = n269 | n270 ;
  assign n272 = n268 | n271 ;
  assign n273 = n267 | n272 ;
  assign n274 = n259 | n273 ;
  assign n275 = n58 & n69 ;
  assign n276 = n69 & n71 ;
  assign n277 = n275 | n276 ;
  assign n278 = n98 & n143 ;
  assign n279 = ~n85 & n157 ;
  assign n280 = n278 | n279 ;
  assign n281 = n277 | n280 ;
  assign n282 = n274 | n281 ;
  assign n283 = n250 | n282 ;
  assign n284 = n71 & n183 ;
  assign n285 = n69 & n94 ;
  assign n286 = n284 | n285 ;
  assign n287 = n58 & n143 ;
  assign n288 = ~x24 & n77 ;
  assign n289 = n130 & n288 ;
  assign n290 = ~x23 & n289 ;
  assign n291 = n287 | n290 ;
  assign n292 = n286 | n291 ;
  assign n293 = n58 & n101 ;
  assign n294 = n88 & n109 ;
  assign n295 = n293 | n294 ;
  assign n296 = n51 & n128 ;
  assign n297 = n54 & n112 ;
  assign n298 = n296 | n297 ;
  assign n299 = n295 | n298 ;
  assign n300 = n292 | n299 ;
  assign n301 = n95 & n130 ;
  assign n302 = ~x24 & n301 ;
  assign n303 = n130 & n183 ;
  assign n304 = n302 | n303 ;
  assign n305 = n88 & n187 ;
  assign n306 = n61 & n235 ;
  assign n307 = ~x24 & n60 ;
  assign n308 = n230 & n307 ;
  assign n309 = n306 | n308 ;
  assign n310 = n305 | n309 ;
  assign n311 = n304 | n310 ;
  assign n312 = n300 | n311 ;
  assign n313 = n60 & n236 ;
  assign n314 = x23 & n313 ;
  assign n315 = n94 & n139 ;
  assign n316 = n314 | n315 ;
  assign n317 = n81 & ~n85 ;
  assign n318 = n67 & n175 ;
  assign n319 = n317 | n318 ;
  assign n320 = n316 | n319 ;
  assign n321 = n61 & n71 ;
  assign n322 = n81 & n94 ;
  assign n323 = n44 & n61 ;
  assign n324 = n322 | n323 ;
  assign n325 = n321 | n324 ;
  assign n326 = n320 | n325 ;
  assign n327 = n312 | n326 ;
  assign n328 = n130 & n187 ;
  assign n329 = n67 & n101 ;
  assign n330 = n102 & n307 ;
  assign n331 = ~x23 & n330 ;
  assign n332 = n329 | n331 ;
  assign n333 = n328 | n332 ;
  assign n334 = n81 & n142 ;
  assign n335 = n51 & ~n73 ;
  assign n336 = n334 | n335 ;
  assign n337 = n142 & n157 ;
  assign n338 = n58 & n183 ;
  assign n339 = n337 | n338 ;
  assign n340 = n336 | n339 ;
  assign n341 = n69 & n98 ;
  assign n342 = n61 & n67 ;
  assign n343 = n341 | n342 ;
  assign n344 = n340 | n343 ;
  assign n345 = n109 & n142 ;
  assign n346 = n107 & n142 ;
  assign n347 = n102 & n183 ;
  assign n348 = n346 | n347 ;
  assign n349 = n345 | n348 ;
  assign n350 = n78 & n235 ;
  assign n351 = ~x30 & n159 ;
  assign n352 = n350 | n351 ;
  assign n353 = n349 | n352 ;
  assign n354 = n344 | n353 ;
  assign n355 = n333 | n354 ;
  assign n356 = n112 & n128 ;
  assign n357 = n79 & n101 ;
  assign n358 = n356 | n357 ;
  assign n359 = n44 & n175 ;
  assign n360 = n44 & n107 ;
  assign n361 = n359 | n360 ;
  assign n362 = n54 & n98 ;
  assign n363 = n78 & n88 ;
  assign n364 = n362 | n363 ;
  assign n365 = n361 | n364 ;
  assign n366 = n358 | n365 ;
  assign n367 = n235 & n251 ;
  assign n368 = ~x23 & n367 ;
  assign n369 = n58 & n120 ;
  assign n370 = ~x26 & n369 ;
  assign n371 = n368 | n370 ;
  assign n372 = n71 & n128 ;
  assign n373 = n98 & n101 ;
  assign n374 = n79 & n128 ;
  assign n375 = n373 | n374 ;
  assign n376 = n372 | n375 ;
  assign n377 = n371 | n376 ;
  assign n378 = n102 & n143 ;
  assign n379 = n94 & n175 ;
  assign n380 = n101 & n112 ;
  assign n381 = n379 | n380 ;
  assign n382 = n378 | n381 ;
  assign n383 = n377 | n382 ;
  assign n384 = n366 | n383 ;
  assign n385 = n355 | n384 ;
  assign n386 = n327 | n385 ;
  assign n387 = n283 | n386 ;
  assign n388 = n170 | n387 ;
  assign n389 = n42 | n57 ;
  assign n390 = x31 & n389 ;
  assign n391 = n133 | n188 ;
  assign n392 = n81 & n98 ;
  assign n393 = n297 | n392 ;
  assign n394 = n335 | n380 ;
  assign n395 = n393 | n394 ;
  assign n396 = n98 & n157 ;
  assign n397 = n94 & n231 ;
  assign n398 = n396 | n397 ;
  assign n399 = n395 | n398 ;
  assign n400 = n391 | n399 ;
  assign n401 = n71 & n251 ;
  assign n402 = ~x23 & n401 ;
  assign n403 = n308 | n402 ;
  assign n404 = n191 | n221 ;
  assign n405 = n88 & n183 ;
  assign n406 = n67 & n251 ;
  assign n407 = ~x23 & n406 ;
  assign n408 = n405 | n407 ;
  assign n409 = n404 | n408 ;
  assign n410 = n403 | n409 ;
  assign n411 = n400 | n410 ;
  assign n412 = n78 & n112 ;
  assign n413 = n109 & n112 ;
  assign n414 = n356 | n413 ;
  assign n415 = n412 | n414 ;
  assign n416 = n78 & n130 ;
  assign n417 = n278 | n416 ;
  assign n418 = n415 | n417 ;
  assign n419 = ~n85 & n107 ;
  assign n420 = n368 | n419 ;
  assign n421 = n418 | n420 ;
  assign n422 = n84 & n121 ;
  assign n423 = n346 | n422 ;
  assign n424 = n232 | n423 ;
  assign n425 = n421 | n424 ;
  assign n426 = n411 | n425 ;
  assign n427 = n99 | n241 ;
  assign n428 = x23 & n401 ;
  assign n429 = n198 | n428 ;
  assign n430 = n427 | n429 ;
  assign n431 = n175 & n235 ;
  assign n432 = n139 & n235 ;
  assign n433 = n431 | n432 ;
  assign n434 = n44 & ~n73 ;
  assign n435 = ~n73 & n79 ;
  assign n436 = n434 | n435 ;
  assign n437 = n433 | n436 ;
  assign n438 = n430 | n437 ;
  assign n439 = n426 | n438 ;
  assign n440 = n61 & n98 ;
  assign n441 = n142 & n187 ;
  assign n442 = n98 & n109 ;
  assign n443 = n206 | n442 ;
  assign n444 = n441 | n443 ;
  assign n445 = n440 | n444 ;
  assign n446 = n112 & n143 ;
  assign n447 = n197 | n446 ;
  assign n448 = n341 | n373 ;
  assign n449 = n121 & n143 ;
  assign n450 = n269 | n449 ;
  assign n451 = n448 | n450 ;
  assign n452 = n447 | n451 ;
  assign n453 = n445 | n452 ;
  assign n454 = n112 & n175 ;
  assign n455 = n69 & n79 ;
  assign n456 = n78 & n121 ;
  assign n457 = n455 | n456 ;
  assign n458 = n215 | n254 ;
  assign n459 = n457 | n458 ;
  assign n460 = n454 | n459 ;
  assign n461 = n453 | n460 ;
  assign n462 = n439 | n461 ;
  assign n463 = n112 & n171 ;
  assign n464 = x24 & n463 ;
  assign n465 = n98 & n183 ;
  assign n466 = n306 | n465 ;
  assign n467 = n464 | n466 ;
  assign n468 = n81 & n130 ;
  assign n469 = n95 & n112 ;
  assign n470 = x24 & n469 ;
  assign n471 = n98 & n175 ;
  assign n472 = n256 | n471 ;
  assign n473 = n470 | n472 ;
  assign n474 = n468 | n473 ;
  assign n475 = n467 | n474 ;
  assign n476 = n184 | n294 ;
  assign n477 = n112 & n139 ;
  assign n478 = n261 | n477 ;
  assign n479 = n476 | n478 ;
  assign n480 = ~n73 & n88 ;
  assign n481 = n148 | n480 ;
  assign n482 = n379 | n481 ;
  assign n483 = n479 | n482 ;
  assign n484 = n475 | n483 ;
  assign n485 = n130 & n143 ;
  assign n486 = n290 | n485 ;
  assign n487 = ~n85 & n143 ;
  assign n488 = n69 & n88 ;
  assign n489 = n338 | n488 ;
  assign n490 = n487 | n489 ;
  assign n491 = n486 | n490 ;
  assign n492 = n484 | n491 ;
  assign n493 = n98 & n107 ;
  assign n494 = n51 & n183 ;
  assign n495 = n493 | n494 ;
  assign n496 = n275 | n495 ;
  assign n497 = n67 & n139 ;
  assign n498 = n350 | n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n112 & n187 ;
  assign n501 = n337 | n500 ;
  assign n502 = n499 | n501 ;
  assign n503 = n129 | n218 ;
  assign n504 = n104 | n362 ;
  assign n505 = n257 | n504 ;
  assign n506 = n52 | n60 ;
  assign n507 = ~n72 & n506 ;
  assign n508 = n121 & n507 ;
  assign n509 = n151 | n508 ;
  assign n510 = n505 | n509 ;
  assign n511 = n503 | n510 ;
  assign n512 = n502 | n511 ;
  assign n513 = n492 | n512 ;
  assign n514 = n462 | n513 ;
  assign n515 = n45 | n85 ;
  assign n516 = x24 & ~n515 ;
  assign n517 = x26 & n264 ;
  assign n518 = ~n85 & n109 ;
  assign n519 = n517 | n518 ;
  assign n520 = n516 | n519 ;
  assign n521 = ~n45 & n142 ;
  assign n522 = ~x24 & n521 ;
  assign n523 = n520 | n522 ;
  assign n524 = n51 & n109 ;
  assign n525 = n293 | n524 ;
  assign n526 = n112 & n183 ;
  assign n527 = n113 | n526 ;
  assign n528 = n143 & n235 ;
  assign n529 = n527 | n528 ;
  assign n530 = n525 | n529 ;
  assign n531 = n70 | n329 ;
  assign n532 = n226 | n531 ;
  assign n533 = n67 & n128 ;
  assign n534 = n67 & n109 ;
  assign n535 = n533 | n534 ;
  assign n536 = n363 | n535 ;
  assign n537 = n532 | n536 ;
  assign n538 = n530 | n537 ;
  assign n539 = n523 | n538 ;
  assign n540 = n150 | n286 ;
  assign n541 = ~n45 & n71 ;
  assign n542 = n142 & n251 ;
  assign n543 = n541 | n542 ;
  assign n544 = n540 | n543 ;
  assign n545 = n94 & n183 ;
  assign n546 = n71 & n109 ;
  assign n547 = n125 | n546 ;
  assign n548 = n545 | n547 ;
  assign n549 = n544 | n548 ;
  assign n550 = n58 & n109 ;
  assign n551 = n296 | n550 ;
  assign n552 = n233 | n351 ;
  assign n553 = n551 | n552 ;
  assign n554 = n54 & n67 ;
  assign n555 = n370 | n554 ;
  assign n556 = n58 & n187 ;
  assign n557 = n58 & n128 ;
  assign n558 = n556 | n557 ;
  assign n559 = n48 | n558 ;
  assign n560 = n555 | n559 ;
  assign n561 = n553 | n560 ;
  assign n562 = n549 | n561 ;
  assign n563 = n539 | n562 ;
  assign n564 = n514 | n563 ;
  assign n565 = n77 & n79 ;
  assign n566 = ~x24 & n565 ;
  assign n567 = n51 & n175 ;
  assign n568 = n147 | n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = n297 | n470 ;
  assign n571 = n569 | n570 ;
  assign n572 = n279 | n465 ;
  assign n573 = n60 & n71 ;
  assign n574 = ~n72 & n573 ;
  assign n575 = n226 | n574 ;
  assign n576 = n572 | n575 ;
  assign n577 = n571 | n576 ;
  assign n578 = n368 | n442 ;
  assign n579 = n362 | n578 ;
  assign n580 = n433 | n579 ;
  assign n581 = n71 & n84 ;
  assign n582 = n480 | n581 ;
  assign n583 = n123 | n582 ;
  assign n584 = n580 | n583 ;
  assign n585 = n577 | n584 ;
  assign n586 = n44 & n187 ;
  assign n587 = n225 | n586 ;
  assign n588 = n209 | n587 ;
  assign n589 = n139 & n142 ;
  assign n590 = n125 | n589 ;
  assign n591 = n51 & n107 ;
  assign n592 = n337 | n591 ;
  assign n593 = n51 & n143 ;
  assign n594 = n99 | n593 ;
  assign n595 = n592 | n594 ;
  assign n596 = n590 | n595 ;
  assign n597 = n588 | n596 ;
  assign n598 = n585 | n597 ;
  assign n599 = n55 | n485 ;
  assign n600 = n44 & n69 ;
  assign n601 = n70 | n600 ;
  assign n602 = n358 | n601 ;
  assign n603 = n599 | n602 ;
  assign n604 = n409 | n603 ;
  assign n605 = n165 | n413 ;
  assign n606 = n134 | n605 ;
  assign n607 = n380 | n534 ;
  assign n608 = n606 | n607 ;
  assign n609 = n604 | n608 ;
  assign n610 = n598 | n609 ;
  assign n611 = x24 & n47 ;
  assign n612 = n503 | n611 ;
  assign n613 = n51 & n101 ;
  assign n614 = n44 & n54 ;
  assign n615 = n613 | n614 ;
  assign n616 = n58 & n107 ;
  assign n617 = n79 & n143 ;
  assign n618 = n73 | n85 ;
  assign n619 = ~n617 & n618 ;
  assign n620 = ~n616 & n619 ;
  assign n621 = ~n615 & n620 ;
  assign n622 = ~n612 & n621 ;
  assign n623 = n51 & n78 ;
  assign n624 = n101 & n121 ;
  assign n625 = n189 | n624 ;
  assign n626 = n623 | n625 ;
  assign n627 = n108 | n124 ;
  assign n628 = n109 & n121 ;
  assign n629 = n305 | n628 ;
  assign n630 = n627 | n629 ;
  assign n631 = n626 | n630 ;
  assign n632 = n622 & ~n631 ;
  assign n633 = n174 | n241 ;
  assign n634 = n261 | n633 ;
  assign n635 = n79 & n157 ;
  assign n636 = n238 | n635 ;
  assign n637 = n133 | n334 ;
  assign n638 = n636 | n637 ;
  assign n639 = n634 | n638 ;
  assign n640 = n71 & n157 ;
  assign n641 = n533 | n640 ;
  assign n642 = n639 | n641 ;
  assign n643 = n110 | n254 ;
  assign n644 = n201 | n363 ;
  assign n645 = n500 | n644 ;
  assign n646 = n643 | n645 ;
  assign n647 = n79 & n187 ;
  assign n648 = n306 | n341 ;
  assign n649 = n647 | n648 ;
  assign n650 = n498 | n649 ;
  assign n651 = n646 | n650 ;
  assign n652 = n642 | n651 ;
  assign n653 = n632 & ~n652 ;
  assign n654 = ~n610 & n653 ;
  assign n655 = n94 & n114 ;
  assign n656 = ~x24 & n655 ;
  assign n657 = n62 | n264 ;
  assign n658 = n656 | n657 ;
  assign n659 = n94 & n128 ;
  assign n660 = n90 | n659 ;
  assign n661 = n58 & n78 ;
  assign n662 = n67 & n107 ;
  assign n663 = n661 | n662 ;
  assign n664 = n449 | n663 ;
  assign n665 = n660 | n664 ;
  assign n666 = n658 | n665 ;
  assign n667 = n69 & n102 ;
  assign n668 = n402 | n667 ;
  assign n669 = n68 & ~n515 ;
  assign n670 = n179 | n308 ;
  assign n671 = n669 | n670 ;
  assign n672 = n668 | n671 ;
  assign n673 = n666 | n672 ;
  assign n674 = n67 & n143 ;
  assign n675 = n256 | n674 ;
  assign n676 = ~n85 & n231 ;
  assign n677 = x23 & n676 ;
  assign n678 = n61 & n142 ;
  assign n679 = ~n85 & n175 ;
  assign n680 = n678 | n679 ;
  assign n681 = n677 | n680 ;
  assign n682 = n675 | n681 ;
  assign n683 = n178 | n416 ;
  assign n684 = n74 | n265 ;
  assign n685 = n683 | n684 ;
  assign n686 = n682 | n685 ;
  assign n687 = n673 | n686 ;
  assign n688 = ~n85 & n128 ;
  assign n689 = n51 & n139 ;
  assign n690 = n347 | n689 ;
  assign n691 = n688 | n690 ;
  assign n692 = n242 | n260 ;
  assign n693 = n338 | n692 ;
  assign n694 = n691 | n693 ;
  assign n695 = n67 & n187 ;
  assign n696 = n419 | n695 ;
  assign n697 = n192 | n696 ;
  assign n698 = n291 | n697 ;
  assign n699 = n694 | n698 ;
  assign n700 = n79 & n109 ;
  assign n701 = n322 | n374 ;
  assign n702 = n700 | n701 ;
  assign n703 = n699 | n702 ;
  assign n704 = ~n73 & n102 ;
  assign n705 = n428 | n704 ;
  assign n706 = n529 | n705 ;
  assign n707 = n102 & n128 ;
  assign n708 = n144 | n707 ;
  assign n709 = n468 | n708 ;
  assign n710 = n706 | n709 ;
  assign n711 = n206 | n215 ;
  assign n712 = n69 & n142 ;
  assign n713 = n150 | n712 ;
  assign n714 = n711 | n713 ;
  assign n715 = n58 & n175 ;
  assign n716 = n275 | n715 ;
  assign n717 = n714 | n716 ;
  assign n718 = n710 | n717 ;
  assign n719 = n703 | n718 ;
  assign n720 = n687 | n719 ;
  assign n721 = n654 & ~n720 ;
  assign n722 = n226 | n345 ;
  assign n723 = ~x24 & n257 ;
  assign n724 = n412 | n723 ;
  assign n725 = n245 | n374 ;
  assign n726 = n724 | n725 ;
  assign n727 = n722 | n726 ;
  assign n728 = n306 | n677 ;
  assign n729 = n110 | n174 ;
  assign n730 = n188 | n729 ;
  assign n731 = n728 | n730 ;
  assign n732 = n727 | n731 ;
  assign n733 = n485 | n554 ;
  assign n734 = n54 & n94 ;
  assign n735 = n153 | n734 ;
  assign n736 = n733 | n735 ;
  assign n737 = n278 | n695 ;
  assign n738 = n70 | n113 ;
  assign n739 = n737 | n738 ;
  assign n740 = n736 | n739 ;
  assign n741 = n732 | n740 ;
  assign n742 = ~x23 & n397 ;
  assign n743 = n151 | n526 ;
  assign n744 = n742 | n743 ;
  assign n745 = n176 | n407 ;
  assign n746 = n744 | n745 ;
  assign n747 = n315 | n318 ;
  assign n748 = n746 | n747 ;
  assign n749 = n102 & n114 ;
  assign n750 = ~x24 & n749 ;
  assign n751 = n67 & ~n73 ;
  assign n752 = n396 | n751 ;
  assign n753 = n750 | n752 ;
  assign n754 = n371 | n753 ;
  assign n755 = n748 | n754 ;
  assign n756 = n321 | n640 ;
  assign n757 = n164 | n756 ;
  assign n758 = n454 | n471 ;
  assign n759 = n757 | n758 ;
  assign n760 = n755 | n759 ;
  assign n761 = n741 | n760 ;
  assign n762 = n567 | n593 ;
  assign n763 = n440 | n762 ;
  assign n764 = n232 | n342 ;
  assign n765 = n276 | n764 ;
  assign n766 = n290 | n635 ;
  assign n767 = n493 | n613 ;
  assign n768 = n140 | n767 ;
  assign n769 = n766 | n768 ;
  assign n770 = n765 | n769 ;
  assign n771 = n763 | n770 ;
  assign n772 = ~x24 & n581 ;
  assign n773 = n207 | n772 ;
  assign n774 = n360 | n446 ;
  assign n775 = n773 | n774 ;
  assign n776 = n413 | n533 ;
  assign n777 = ~n73 & n121 ;
  assign n778 = n150 | n777 ;
  assign n779 = n776 | n778 ;
  assign n780 = n79 & n81 ;
  assign n781 = n102 & n107 ;
  assign n782 = n780 | n781 ;
  assign n783 = n779 | n782 ;
  assign n784 = n775 | n783 ;
  assign n785 = n771 | n784 ;
  assign n786 = n90 | n269 ;
  assign n787 = n222 | n786 ;
  assign n788 = n456 | n497 ;
  assign n789 = ~n45 & n236 ;
  assign n790 = n788 | n789 ;
  assign n791 = n787 | n790 ;
  assign n792 = n785 | n791 ;
  assign n793 = n402 | n628 ;
  assign n794 = n128 & n235 ;
  assign n795 = n557 | n794 ;
  assign n796 = n793 | n795 ;
  assign n797 = n52 & n72 ;
  assign n798 = n121 & n797 ;
  assign n799 = n334 | n798 ;
  assign n800 = n796 | n799 ;
  assign n801 = n221 | n468 ;
  assign n802 = n172 | n416 ;
  assign n803 = n801 | n802 ;
  assign n804 = n800 | n803 ;
  assign n805 = n284 | n550 ;
  assign n806 = n252 | n268 ;
  assign n807 = n805 | n806 ;
  assign n808 = n147 | n656 ;
  assign n809 = n241 | n528 ;
  assign n810 = n545 | n809 ;
  assign n811 = n808 | n810 ;
  assign n812 = n807 | n811 ;
  assign n813 = n804 | n812 ;
  assign n814 = n323 | n464 ;
  assign n815 = n431 | n662 ;
  assign n816 = n814 | n815 ;
  assign n817 = n103 | n712 ;
  assign n818 = n144 | n817 ;
  assign n819 = n358 | n818 ;
  assign n820 = n487 | n647 ;
  assign n821 = n206 | n820 ;
  assign n822 = n819 | n821 ;
  assign n823 = n256 | n591 ;
  assign n824 = n178 | n378 ;
  assign n825 = n611 | n824 ;
  assign n826 = n823 | n825 ;
  assign n827 = n822 | n826 ;
  assign n828 = n816 | n827 ;
  assign n829 = n813 | n828 ;
  assign n830 = n792 | n829 ;
  assign n831 = n337 | n669 ;
  assign n832 = n189 | n432 ;
  assign n833 = n659 | n832 ;
  assign n834 = n831 | n833 ;
  assign n835 = n78 & ~n85 ;
  assign n836 = n600 | n835 ;
  assign n837 = n218 | n836 ;
  assign n838 = n488 | n616 ;
  assign n839 = n837 | n838 ;
  assign n840 = n834 | n839 ;
  assign n841 = n44 & n143 ;
  assign n842 = n287 | n841 ;
  assign n843 = n359 | n842 ;
  assign n844 = n350 | n373 ;
  assign n845 = n428 | n844 ;
  assign n846 = n843 | n845 ;
  assign n847 = n840 | n846 ;
  assign n848 = n215 | n363 ;
  assign n849 = n260 | n848 ;
  assign n850 = n102 & n157 ;
  assign n851 = n441 | n700 ;
  assign n852 = n850 | n851 ;
  assign n853 = n849 | n852 ;
  assign n854 = n148 | n331 ;
  assign n855 = n63 | n854 ;
  assign n856 = n853 | n855 ;
  assign n857 = n847 | n856 ;
  assign n858 = n830 | n857 ;
  assign n859 = n761 | n858 ;
  assign n860 = n121 & n183 ;
  assign n861 = n82 | n860 ;
  assign n862 = n734 | n861 ;
  assign n863 = x24 & n581 ;
  assign n864 = n210 | n617 ;
  assign n865 = n863 | n864 ;
  assign n866 = n87 | n865 ;
  assign n867 = n862 | n866 ;
  assign n868 = n373 | n704 ;
  assign n869 = n108 | n868 ;
  assign n870 = n867 | n869 ;
  assign n871 = n477 | n623 ;
  assign n872 = n351 | n871 ;
  assign n873 = n465 | n557 ;
  assign n874 = n772 | n873 ;
  assign n875 = n872 | n874 ;
  assign n876 = n220 | n284 ;
  assign n877 = n96 | n322 ;
  assign n878 = n876 | n877 ;
  assign n879 = n223 | n878 ;
  assign n880 = n875 | n879 ;
  assign n881 = n360 | n841 ;
  assign n882 = n237 | n881 ;
  assign n883 = n268 | n297 ;
  assign n884 = n882 | n883 ;
  assign n885 = n335 | n468 ;
  assign n886 = n599 | n885 ;
  assign n887 = n264 | n886 ;
  assign n888 = n884 | n887 ;
  assign n889 = n880 | n888 ;
  assign n890 = n870 | n889 ;
  assign n891 = n615 | n831 ;
  assign n892 = n265 | n315 ;
  assign n893 = n188 | n715 ;
  assign n894 = n892 | n893 ;
  assign n895 = n891 | n894 ;
  assign n896 = n103 | n214 ;
  assign n897 = n895 | n896 ;
  assign n898 = n890 | n897 ;
  assign n899 = n270 | n526 ;
  assign n900 = n90 | n700 ;
  assign n901 = n303 | n689 ;
  assign n902 = n446 | n901 ;
  assign n903 = n900 | n902 ;
  assign n904 = n347 | n679 ;
  assign n905 = n903 | n904 ;
  assign n906 = n147 | n742 ;
  assign n907 = n346 | n508 ;
  assign n908 = n906 | n907 ;
  assign n909 = n905 | n908 ;
  assign n910 = n899 | n909 ;
  assign n911 = n898 | n910 ;
  assign n912 = n44 & n78 ;
  assign n913 = n197 | n912 ;
  assign n914 = n198 | n913 ;
  assign n915 = x24 & n257 ;
  assign n916 = ~n73 & n130 ;
  assign n917 = n254 | n916 ;
  assign n918 = n915 | n917 ;
  assign n919 = n554 | n918 ;
  assign n920 = n914 | n919 ;
  assign n921 = n528 | n850 ;
  assign n922 = n142 & n183 ;
  assign n923 = n616 | n922 ;
  assign n924 = n921 | n923 ;
  assign n925 = n99 | n207 ;
  assign n926 = n924 | n925 ;
  assign n927 = n70 | n144 ;
  assign n928 = n380 | n927 ;
  assign n929 = n200 | n208 ;
  assign n930 = n141 | n345 ;
  assign n931 = n929 | n930 ;
  assign n932 = n928 | n931 ;
  assign n933 = n926 | n932 ;
  assign n934 = n920 | n933 ;
  assign n935 = n338 | n574 ;
  assign n936 = n241 | n441 ;
  assign n937 = n470 | n936 ;
  assign n938 = n935 | n937 ;
  assign n939 = n363 | n480 ;
  assign n940 = n938 | n939 ;
  assign n941 = n215 | n372 ;
  assign n942 = ~n85 & n183 ;
  assign n943 = n238 | n942 ;
  assign n944 = n189 | n943 ;
  assign n945 = n941 | n944 ;
  assign n946 = n374 | n416 ;
  assign n947 = n402 | n695 ;
  assign n948 = n946 | n947 ;
  assign n949 = n945 | n948 ;
  assign n950 = n940 | n949 ;
  assign n951 = n934 | n950 ;
  assign n952 = n911 | n951 ;
  assign n953 = n233 | n493 ;
  assign n954 = n232 | n334 ;
  assign n955 = n953 | n954 ;
  assign n956 = n342 | n677 ;
  assign n957 = n260 | n550 ;
  assign n958 = n956 | n957 ;
  assign n959 = n955 | n958 ;
  assign n960 = n600 | n781 ;
  assign n961 = n518 | n589 ;
  assign n962 = n960 | n961 ;
  assign n963 = n959 | n962 ;
  assign n964 = n392 | n678 ;
  assign n965 = n306 | n396 ;
  assign n966 = n964 | n965 ;
  assign n967 = n745 | n966 ;
  assign n968 = x24 & n749 ;
  assign n969 = n113 | n968 ;
  assign n970 = n431 | n780 ;
  assign n971 = n185 | n970 ;
  assign n972 = n969 | n971 ;
  assign n973 = n967 | n972 ;
  assign n974 = n963 | n973 ;
  assign n975 = n123 | n435 ;
  assign n976 = n151 | n835 ;
  assign n977 = n120 & n142 ;
  assign n978 = n378 | n977 ;
  assign n979 = n976 | n978 ;
  assign n980 = n975 | n979 ;
  assign n981 = n253 | n428 ;
  assign n982 = n980 | n981 ;
  assign n983 = n140 | n341 ;
  assign n984 = n131 | n290 ;
  assign n985 = n983 | n984 ;
  assign n986 = n488 | n712 ;
  assign n987 = n54 & n235 ;
  assign n988 = n986 | n987 ;
  assign n989 = n128 & n130 ;
  assign n990 = n331 | n989 ;
  assign n991 = n988 | n990 ;
  assign n992 = n985 | n991 ;
  assign n993 = n982 | n992 ;
  assign n994 = n974 | n993 ;
  assign n995 = n952 | n994 ;
  assign n996 = n206 | n221 ;
  assign n997 = n200 | n640 ;
  assign n998 = n996 | n997 ;
  assign n999 = n164 | n238 ;
  assign n1000 = n103 | n159 ;
  assign n1001 = n999 | n1000 ;
  assign n1002 = n998 | n1001 ;
  assign n1003 = n668 | n844 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = n232 | n534 ;
  assign n1006 = n71 & n78 ;
  assign n1007 = n454 | n1006 ;
  assign n1008 = n546 | n614 ;
  assign n1009 = n1007 | n1008 ;
  assign n1010 = n1005 | n1009 ;
  assign n1011 = n1004 | n1010 ;
  assign n1012 = n317 | n518 ;
  assign n1013 = n90 | n276 ;
  assign n1014 = n129 | n850 ;
  assign n1015 = n334 | n1014 ;
  assign n1016 = n1013 | n1015 ;
  assign n1017 = n1012 | n1016 ;
  assign n1018 = n55 | n237 ;
  assign n1019 = n99 | n396 ;
  assign n1020 = n183 & n235 ;
  assign n1021 = n356 | n1020 ;
  assign n1022 = n1019 | n1021 ;
  assign n1023 = n134 | n285 ;
  assign n1024 = n257 | n1023 ;
  assign n1025 = n1022 | n1024 ;
  assign n1026 = n1018 | n1025 ;
  assign n1027 = n1017 | n1026 ;
  assign n1028 = n1011 | n1027 ;
  assign n1029 = n338 | n591 ;
  assign n1030 = n526 | n1029 ;
  assign n1031 = ( ~n275 & n515 ) | ( ~n275 & n516 ) | ( n515 & n516 ) ;
  assign n1032 = ~n1030 & n1031 ;
  assign n1033 = n261 | n305 ;
  assign n1034 = n214 | n494 ;
  assign n1035 = n1033 | n1034 ;
  assign n1036 = n302 | n589 ;
  assign n1037 = n1035 | n1036 ;
  assign n1038 = n1032 & ~n1037 ;
  assign n1039 = ~n1028 & n1038 ;
  assign n1040 = n97 | n329 ;
  assign n1041 = n102 & n175 ;
  assign n1042 = n297 | n1041 ;
  assign n1043 = n1040 | n1042 ;
  assign n1044 = n67 & n183 ;
  assign n1045 = n374 | n1044 ;
  assign n1046 = n611 | n1045 ;
  assign n1047 = n1043 | n1046 ;
  assign n1048 = n130 & n157 ;
  assign n1049 = n67 & n231 ;
  assign n1050 = n635 | n1049 ;
  assign n1051 = n1048 | n1050 ;
  assign n1052 = n941 | n1051 ;
  assign n1053 = n1047 | n1052 ;
  assign n1054 = n659 | n863 ;
  assign n1055 = n712 | n1054 ;
  assign n1056 = n87 | n278 ;
  assign n1057 = n1055 | n1056 ;
  assign n1058 = n303 | n623 ;
  assign n1059 = n295 | n1058 ;
  assign n1060 = n184 | n360 ;
  assign n1061 = n1059 | n1060 ;
  assign n1062 = n1057 | n1061 ;
  assign n1063 = n1053 | n1062 ;
  assign n1064 = n500 | n677 ;
  assign n1065 = n434 | n777 ;
  assign n1066 = n191 | n628 ;
  assign n1067 = n1065 | n1066 ;
  assign n1068 = n1064 | n1067 ;
  assign n1069 = n79 & n175 ;
  assign n1070 = n442 | n1069 ;
  assign n1071 = n446 | n661 ;
  assign n1072 = n1070 | n1071 ;
  assign n1073 = n1068 | n1072 ;
  assign n1074 = n121 & n128 ;
  assign n1075 = n485 | n1074 ;
  assign n1076 = n656 | n1075 ;
  assign n1077 = n968 | n1076 ;
  assign n1078 = n1073 | n1077 ;
  assign n1079 = n1063 | n1078 ;
  assign n1080 = n1039 & ~n1079 ;
  assign n1081 = n88 & n101 ;
  assign n1082 = n165 | n1081 ;
  assign n1083 = n392 | n440 ;
  assign n1084 = n104 | n1083 ;
  assign n1085 = n1082 | n1084 ;
  assign n1086 = n101 & n235 ;
  assign n1087 = n308 | n1086 ;
  assign n1088 = n497 | n1087 ;
  assign n1089 = n185 | n772 ;
  assign n1090 = n1088 | n1089 ;
  assign n1091 = n1085 | n1090 ;
  assign n1092 = n407 | n916 ;
  assign n1093 = n892 | n1092 ;
  assign n1094 = n44 & n139 ;
  assign n1095 = n323 | n1094 ;
  assign n1096 = n178 | n780 ;
  assign n1097 = n1095 | n1096 ;
  assign n1098 = n1093 | n1097 ;
  assign n1099 = n1091 | n1098 ;
  assign n1100 = x26 & n977 ;
  assign n1101 = n419 | n1100 ;
  assign n1102 = n700 | n707 ;
  assign n1103 = n233 | n528 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = n1101 | n1104 ;
  assign n1106 = n108 | n912 ;
  assign n1107 = n161 | n922 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = n1105 | n1108 ;
  assign n1110 = n287 | n557 ;
  assign n1111 = n189 | n600 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n477 | n593 ;
  assign n1114 = n860 | n1113 ;
  assign n1115 = n1112 | n1114 ;
  assign n1116 = n1109 | n1115 ;
  assign n1117 = n1099 | n1116 ;
  assign n1118 = n1080 & ~n1117 ;
  assign n1119 = n55 | n74 ;
  assign n1120 = n198 | n915 ;
  assign n1121 = n680 | n1120 ;
  assign n1122 = n1119 | n1121 ;
  assign n1123 = n405 | n1006 ;
  assign n1124 = n689 | n860 ;
  assign n1125 = n1123 | n1124 ;
  assign n1126 = n187 & n235 ;
  assign n1127 = n131 | n1126 ;
  assign n1128 = n1125 | n1127 ;
  assign n1129 = n1122 | n1128 ;
  assign n1130 = n82 | n351 ;
  assign n1131 = n470 | n1130 ;
  assign n1132 = n1129 | n1131 ;
  assign n1133 = n323 | n456 ;
  assign n1134 = n331 | n1133 ;
  assign n1135 = n470 | n780 ;
  assign n1136 = n1134 | n1135 ;
  assign n1137 = n392 | n674 ;
  assign n1138 = n160 | n1137 ;
  assign n1139 = n268 | n912 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = n1136 | n1140 ;
  assign n1142 = n1132 | n1141 ;
  assign n1143 = n761 | n1142 ;
  assign n1144 = n134 | n611 ;
  assign n1145 = n46 & n94 ;
  assign n1146 = n141 | n1145 ;
  assign n1147 = n1144 | n1146 ;
  assign n1148 = n244 | n455 ;
  assign n1149 = n99 | n1148 ;
  assign n1150 = n1147 | n1149 ;
  assign n1151 = n302 | n623 ;
  assign n1152 = n91 | n1151 ;
  assign n1153 = n618 & ~n863 ;
  assign n1154 = ~n1152 & n1153 ;
  assign n1155 = ~n1150 & n1154 ;
  assign n1156 = ~n366 & n1155 ;
  assign n1157 = n297 | n850 ;
  assign n1158 = n163 | n1157 ;
  assign n1159 = n586 | n987 ;
  assign n1160 = n1158 | n1159 ;
  assign n1161 = n294 | n968 ;
  assign n1162 = n589 | n616 ;
  assign n1163 = n206 | n1162 ;
  assign n1164 = n1161 | n1163 ;
  assign n1165 = n1160 | n1164 ;
  assign n1166 = n192 | n557 ;
  assign n1167 = n793 | n1166 ;
  assign n1168 = n1165 | n1167 ;
  assign n1169 = n208 | n667 ;
  assign n1170 = n223 | n1169 ;
  assign n1171 = n150 | n296 ;
  assign n1172 = n225 | n916 ;
  assign n1173 = n200 | n688 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = n1171 | n1174 ;
  assign n1176 = n101 & n130 ;
  assign n1177 = n218 | n1176 ;
  assign n1178 = n123 | n140 ;
  assign n1179 = n1177 | n1178 ;
  assign n1180 = n1175 | n1179 ;
  assign n1181 = n1170 | n1180 ;
  assign n1182 = n1168 | n1181 ;
  assign n1183 = n1156 & ~n1182 ;
  assign n1184 = n841 | n942 ;
  assign n1185 = n129 | n1044 ;
  assign n1186 = n480 | n1185 ;
  assign n1187 = n615 | n1186 ;
  assign n1188 = n1184 | n1187 ;
  assign n1189 = n284 | n308 ;
  assign n1190 = n766 | n1189 ;
  assign n1191 = n1188 | n1190 ;
  assign n1192 = n191 | n823 ;
  assign n1193 = ~x26 & n977 ;
  assign n1194 = n715 | n1193 ;
  assign n1195 = n1192 | n1194 ;
  assign n1196 = n494 | n517 ;
  assign n1197 = n605 | n1196 ;
  assign n1198 = n1195 | n1197 ;
  assign n1199 = n293 | n1094 ;
  assign n1200 = n572 | n1199 ;
  assign n1201 = n1107 | n1200 ;
  assign n1202 = n184 | n214 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = n1198 | n1203 ;
  assign n1205 = n1191 | n1204 ;
  assign n1206 = n1183 & ~n1205 ;
  assign n1207 = ~n1143 & n1206 ;
  assign n1208 = n419 | n860 ;
  assign n1209 = n55 | n293 ;
  assign n1210 = n436 | n1209 ;
  assign n1211 = n1208 | n1210 ;
  assign n1212 = n110 | n322 ;
  assign n1213 = n379 | n1212 ;
  assign n1214 = n1211 | n1213 ;
  assign n1215 = n704 | n986 ;
  assign n1216 = n334 | n556 ;
  assign n1217 = n197 | n1216 ;
  assign n1218 = n683 | n722 ;
  assign n1219 = n1217 | n1218 ;
  assign n1220 = n1215 | n1219 ;
  assign n1221 = n290 | n351 ;
  assign n1222 = n1220 | n1221 ;
  assign n1223 = n1214 | n1222 ;
  assign n1224 = n97 | n176 ;
  assign n1225 = n456 | n1224 ;
  assign n1226 = n173 | n441 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = n160 | n613 ;
  assign n1229 = n337 | n412 ;
  assign n1230 = n1228 | n1229 ;
  assign n1231 = n1227 | n1230 ;
  assign n1232 = n1223 | n1231 ;
  assign n1233 = n396 | n989 ;
  assign n1234 = n465 | n1233 ;
  assign n1235 = n1161 | n1234 ;
  assign n1236 = n80 | n1020 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = n524 | n593 ;
  assign n1239 = n218 | n1238 ;
  assign n1240 = n297 | n517 ;
  assign n1241 = n335 | n357 ;
  assign n1242 = n207 | n1241 ;
  assign n1243 = n1240 | n1242 ;
  assign n1244 = n1239 | n1243 ;
  assign n1245 = n1237 | n1244 ;
  assign n1246 = n1232 | n1245 ;
  assign n1247 = n260 | n581 ;
  assign n1248 = n656 | n1247 ;
  assign n1249 = n333 | n1248 ;
  assign n1250 = n210 | n983 ;
  assign n1251 = n944 | n1250 ;
  assign n1252 = n1249 | n1251 ;
  assign n1253 = n174 | n487 ;
  assign n1254 = n550 | n723 ;
  assign n1255 = n1253 | n1254 ;
  assign n1256 = n470 | n844 ;
  assign n1257 = n480 | n528 ;
  assign n1258 = n628 | n1257 ;
  assign n1259 = n1256 | n1258 ;
  assign n1260 = n735 | n1259 ;
  assign n1261 = n1255 | n1260 ;
  assign n1262 = n1252 | n1261 ;
  assign n1263 = n413 | n617 ;
  assign n1264 = n374 | n534 ;
  assign n1265 = n1263 | n1264 ;
  assign n1266 = n953 | n1265 ;
  assign n1267 = n296 | n446 ;
  assign n1268 = n346 | n1267 ;
  assign n1269 = n202 | n1268 ;
  assign n1270 = n1266 | n1269 ;
  assign n1271 = n449 | n927 ;
  assign n1272 = n261 | n321 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = n1270 | n1273 ;
  assign n1275 = n124 | n1012 ;
  assign n1276 = n74 | n614 ;
  assign n1277 = n494 | n922 ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = n1275 | n1278 ;
  assign n1280 = n1274 | n1279 ;
  assign n1281 = n1262 | n1280 ;
  assign n1282 = n1246 | n1281 ;
  assign n1283 = n497 | n1014 ;
  assign n1284 = n1151 | n1283 ;
  assign n1285 = n222 | n254 ;
  assign n1286 = n1284 | n1285 ;
  assign n1287 = n241 | n516 ;
  assign n1288 = n141 | n198 ;
  assign n1289 = n1287 | n1288 ;
  assign n1290 = n1286 | n1289 ;
  assign n1291 = n103 | n225 ;
  assign n1292 = n253 | n284 ;
  assign n1293 = n1291 | n1292 ;
  assign n1294 = n237 | n611 ;
  assign n1295 = n391 | n1294 ;
  assign n1296 = n1293 | n1295 ;
  assign n1297 = n1290 | n1296 ;
  assign n1298 = n402 | n546 ;
  assign n1299 = n1110 | n1298 ;
  assign n1300 = n370 | n616 ;
  assign n1301 = n404 | n1300 ;
  assign n1302 = n275 | n1086 ;
  assign n1303 = n567 | n1044 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = n781 | n1304 ;
  assign n1306 = n1301 | n1305 ;
  assign n1307 = n1299 | n1306 ;
  assign n1308 = n356 | n591 ;
  assign n1309 = n104 | n1308 ;
  assign n1310 = n368 | n679 ;
  assign n1311 = n279 | n689 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = n1309 | n1312 ;
  assign n1314 = n1307 | n1313 ;
  assign n1315 = n1297 | n1314 ;
  assign n1316 = n1282 | n1315 ;
  assign n1317 = n192 | n781 ;
  assign n1318 = n241 | n350 ;
  assign n1319 = n656 | n1318 ;
  assign n1320 = n1163 | n1319 ;
  assign n1321 = n1317 | n1320 ;
  assign n1322 = n880 | n1321 ;
  assign n1323 = n131 | n185 ;
  assign n1324 = n379 | n1323 ;
  assign n1325 = n134 | n396 ;
  assign n1326 = n1324 | n1325 ;
  assign n1327 = n363 | n440 ;
  assign n1328 = n554 | n1327 ;
  assign n1329 = n1326 | n1328 ;
  assign n1330 = n1322 | n1329 ;
  assign n1331 = n245 | n533 ;
  assign n1332 = n94 & n101 ;
  assign n1333 = n586 | n1332 ;
  assign n1334 = n1331 | n1333 ;
  assign n1335 = n756 | n1334 ;
  assign n1336 = n946 | n969 ;
  assign n1337 = n1335 | n1336 ;
  assign n1338 = n1126 | n1177 ;
  assign n1339 = n470 | n695 ;
  assign n1340 = n257 | n1339 ;
  assign n1341 = n1338 | n1340 ;
  assign n1342 = n1337 | n1341 ;
  assign n1343 = n1330 | n1342 ;
  assign n1344 = n663 | n987 ;
  assign n1345 = n197 | n238 ;
  assign n1346 = n1344 | n1345 ;
  assign n1347 = n104 | n742 ;
  assign n1348 = n373 | n487 ;
  assign n1349 = n1347 | n1348 ;
  assign n1350 = n1346 | n1349 ;
  assign n1351 = n419 | n942 ;
  assign n1352 = n275 | n432 ;
  assign n1353 = n144 | n1352 ;
  assign n1354 = n1082 | n1353 ;
  assign n1355 = n1351 | n1354 ;
  assign n1356 = n1350 | n1355 ;
  assign n1357 = n317 | n372 ;
  assign n1358 = n208 | n242 ;
  assign n1359 = n617 | n1358 ;
  assign n1360 = n446 | n494 ;
  assign n1361 = n1074 | n1360 ;
  assign n1362 = n1359 | n1361 ;
  assign n1363 = n1357 | n1362 ;
  assign n1364 = n70 | n712 ;
  assign n1365 = n210 | n480 ;
  assign n1366 = n1148 | n1365 ;
  assign n1367 = n1364 | n1366 ;
  assign n1368 = n1363 | n1367 ;
  assign n1369 = n1356 | n1368 ;
  assign n1370 = n287 | n428 ;
  assign n1371 = n150 | n297 ;
  assign n1372 = n454 | n1371 ;
  assign n1373 = n1370 | n1372 ;
  assign n1374 = n110 | n611 ;
  assign n1375 = n407 | n689 ;
  assign n1376 = n1374 | n1375 ;
  assign n1377 = n1373 | n1376 ;
  assign n1378 = n1020 | n1041 ;
  assign n1379 = n253 | n750 ;
  assign n1380 = n160 | n302 ;
  assign n1381 = n1379 | n1380 ;
  assign n1382 = n1378 | n1381 ;
  assign n1383 = n1377 | n1382 ;
  assign n1384 = n306 | n335 ;
  assign n1385 = n1005 | n1384 ;
  assign n1386 = n254 | n501 ;
  assign n1387 = n1385 | n1386 ;
  assign n1388 = n48 | n215 ;
  assign n1389 = n198 | n278 ;
  assign n1390 = n1388 | n1389 ;
  assign n1391 = n442 | n704 ;
  assign n1392 = n108 | n526 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = n1390 | n1393 ;
  assign n1395 = n1387 | n1394 ;
  assign n1396 = n1383 | n1395 ;
  assign n1397 = n1369 | n1396 ;
  assign n1398 = n1343 | n1397 ;
  assign n1399 = n133 | n206 ;
  assign n1400 = n287 | n1399 ;
  assign n1401 = n173 | n781 ;
  assign n1402 = n1400 | n1401 ;
  assign n1403 = n332 | n1088 ;
  assign n1404 = n1402 | n1403 ;
  assign n1405 = n487 | n1193 ;
  assign n1406 = n218 | n337 ;
  assign n1407 = n1405 | n1406 ;
  assign n1408 = n237 | n469 ;
  assign n1409 = n380 | n434 ;
  assign n1410 = n1408 | n1409 ;
  assign n1411 = n1407 | n1410 ;
  assign n1412 = n1404 | n1411 ;
  assign n1413 = n350 | n678 ;
  assign n1414 = n556 | n715 ;
  assign n1415 = n99 | n1048 ;
  assign n1416 = n1414 | n1415 ;
  assign n1417 = n1413 | n1416 ;
  assign n1418 = n1412 | n1417 ;
  assign n1419 = n454 | n841 ;
  assign n1420 = n278 | n341 ;
  assign n1421 = n197 | n1420 ;
  assign n1422 = n1419 | n1421 ;
  assign n1423 = n131 | n351 ;
  assign n1424 = n1422 | n1423 ;
  assign n1425 = n48 | n368 ;
  assign n1426 = n661 | n1425 ;
  assign n1427 = n71 & n263 ;
  assign n1428 = n708 | n1427 ;
  assign n1429 = n500 | n1081 ;
  assign n1430 = n1428 | n1429 ;
  assign n1431 = n1426 | n1430 ;
  assign n1432 = n1424 | n1431 ;
  assign n1433 = n1418 | n1432 ;
  assign n1434 = n328 | n480 ;
  assign n1435 = ~n163 & n618 ;
  assign n1436 = ~n1434 & n1435 ;
  assign n1437 = n222 | n524 ;
  assign n1438 = n1436 & ~n1437 ;
  assign n1439 = n245 | n674 ;
  assign n1440 = n1094 | n1439 ;
  assign n1441 = n1438 & ~n1440 ;
  assign n1442 = n613 | n628 ;
  assign n1443 = n801 | n1442 ;
  assign n1444 = n140 | n617 ;
  assign n1445 = n1443 | n1444 ;
  assign n1446 = n1441 & ~n1445 ;
  assign n1447 = n178 | n465 ;
  assign n1448 = n113 | n441 ;
  assign n1449 = n1447 | n1448 ;
  assign n1450 = n656 | n1449 ;
  assign n1451 = ~x24 & n573 ;
  assign n1452 = n215 | n1451 ;
  assign n1453 = n1450 | n1452 ;
  assign n1454 = n412 | n1148 ;
  assign n1455 = n364 | n1454 ;
  assign n1456 = n600 | n777 ;
  assign n1457 = n677 | n723 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = n1455 | n1458 ;
  assign n1460 = n1453 | n1459 ;
  assign n1461 = n1446 & ~n1460 ;
  assign n1462 = n370 | n679 ;
  assign n1463 = n207 | n396 ;
  assign n1464 = n210 | n293 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = n1462 | n1465 ;
  assign n1467 = n97 | n976 ;
  assign n1468 = n762 | n1467 ;
  assign n1469 = n1466 | n1468 ;
  assign n1470 = n432 | n772 ;
  assign n1471 = n150 | n1470 ;
  assign n1472 = n1379 | n1471 ;
  assign n1473 = n1469 | n1472 ;
  assign n1474 = n270 | n435 ;
  assign n1475 = n198 | n1474 ;
  assign n1476 = n108 | n208 ;
  assign n1477 = n1475 | n1476 ;
  assign n1478 = n1473 | n1477 ;
  assign n1479 = n1461 & ~n1478 ;
  assign n1480 = ~n1433 & n1479 ;
  assign n1481 = n185 | n700 ;
  assign n1482 = n346 | n1481 ;
  assign n1483 = n87 | n1482 ;
  assign n1484 = n486 | n1483 ;
  assign n1485 = n379 | n518 ;
  assign n1486 = n200 | n591 ;
  assign n1487 = n243 | n1486 ;
  assign n1488 = n1485 | n1487 ;
  assign n1489 = n90 | n123 ;
  assign n1490 = n160 | n1489 ;
  assign n1491 = n1488 | n1490 ;
  assign n1492 = n275 | n751 ;
  assign n1493 = n153 | n1492 ;
  assign n1494 = n550 | n689 ;
  assign n1495 = n614 | n1494 ;
  assign n1496 = n1493 | n1495 ;
  assign n1497 = n1491 | n1496 ;
  assign n1498 = n1484 | n1497 ;
  assign n1499 = n174 | n190 ;
  assign n1500 = n322 | n402 ;
  assign n1501 = n260 | n360 ;
  assign n1502 = n1500 | n1501 ;
  assign n1503 = n1499 | n1502 ;
  assign n1504 = n419 | n922 ;
  assign n1505 = n471 | n1176 ;
  assign n1506 = n1504 | n1505 ;
  assign n1507 = n1503 | n1506 ;
  assign n1508 = n1498 | n1507 ;
  assign n1509 = n265 | n528 ;
  assign n1510 = n1144 | n1509 ;
  assign n1511 = n158 & n175 ;
  assign n1512 = n296 | n1511 ;
  assign n1513 = n164 | n306 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = n334 | n1119 ;
  assign n1516 = n1514 | n1515 ;
  assign n1517 = n1510 | n1516 ;
  assign n1518 = n695 | n704 ;
  assign n1519 = n449 | n1518 ;
  assign n1520 = n342 | n1519 ;
  assign n1521 = n256 | n416 ;
  assign n1522 = n268 | n1521 ;
  assign n1523 = n722 | n1522 ;
  assign n1524 = n303 | n408 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = n1520 | n1525 ;
  assign n1527 = n1517 | n1526 ;
  assign n1528 = n1508 | n1527 ;
  assign n1529 = n1480 & ~n1528 ;
  assign n1530 = n1287 | n1477 ;
  assign n1531 = n453 | n1530 ;
  assign n1532 = n148 | n589 ;
  assign n1533 = n178 | n346 ;
  assign n1534 = n1126 | n1533 ;
  assign n1535 = n1532 | n1534 ;
  assign n1536 = n1215 | n1535 ;
  assign n1537 = n402 | n617 ;
  assign n1538 = n1041 | n1048 ;
  assign n1539 = n1033 | n1538 ;
  assign n1540 = n1537 | n1539 ;
  assign n1541 = n1536 | n1540 ;
  assign n1542 = n150 | n1193 ;
  assign n1543 = n968 | n1020 ;
  assign n1544 = n1542 | n1543 ;
  assign n1545 = n1541 | n1544 ;
  assign n1546 = n1531 | n1545 ;
  assign n1547 = n296 | n359 ;
  assign n1548 = n322 | n1547 ;
  assign n1549 = n1510 | n1548 ;
  assign n1550 = n141 | n244 ;
  assign n1551 = n1291 | n1550 ;
  assign n1552 = n1549 | n1551 ;
  assign n1553 = n1546 | n1552 ;
  assign n1554 = n428 | n667 ;
  assign n1555 = n165 | n644 ;
  assign n1556 = n1554 | n1555 ;
  assign n1557 = n360 | n700 ;
  assign n1558 = n715 | n1176 ;
  assign n1559 = n1557 | n1558 ;
  assign n1560 = n284 | n780 ;
  assign n1561 = n153 | n1560 ;
  assign n1562 = n1559 | n1561 ;
  assign n1563 = n1556 | n1562 ;
  assign n1564 = n188 | n335 ;
  assign n1565 = n337 | n1564 ;
  assign n1566 = n1130 | n1565 ;
  assign n1567 = n1255 | n1566 ;
  assign n1568 = n1563 | n1567 ;
  assign n1569 = n412 | n989 ;
  assign n1570 = n753 | n1569 ;
  assign n1571 = n297 | n777 ;
  assign n1572 = n160 | n1571 ;
  assign n1573 = n695 | n707 ;
  assign n1574 = n1572 | n1573 ;
  assign n1575 = n1570 | n1574 ;
  assign n1576 = n374 | n1332 ;
  assign n1577 = n232 | n1576 ;
  assign n1578 = n659 | n1577 ;
  assign n1579 = n163 | n405 ;
  assign n1580 = n238 | n912 ;
  assign n1581 = n1579 | n1580 ;
  assign n1582 = n1578 | n1581 ;
  assign n1583 = n1575 | n1582 ;
  assign n1584 = n1568 | n1583 ;
  assign n1585 = n677 | n1134 ;
  assign n1586 = n125 | n233 ;
  assign n1587 = n1012 | n1586 ;
  assign n1588 = n1585 | n1587 ;
  assign n1589 = n474 | n601 ;
  assign n1590 = n567 | n635 ;
  assign n1591 = n477 | n554 ;
  assign n1592 = n1590 | n1591 ;
  assign n1593 = n303 | n987 ;
  assign n1594 = n294 | n624 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = n1592 | n1595 ;
  assign n1597 = n1589 | n1596 ;
  assign n1598 = n1588 | n1597 ;
  assign n1599 = n1584 | n1598 ;
  assign n1600 = n1553 | n1599 ;
  assign n1601 = n335 | n661 ;
  assign n1602 = n428 | n617 ;
  assign n1603 = n493 | n556 ;
  assign n1604 = n1602 | n1603 ;
  assign n1605 = n1601 | n1604 ;
  assign n1606 = n338 | n794 ;
  assign n1607 = n125 | n659 ;
  assign n1608 = n1606 | n1607 ;
  assign n1609 = n1605 | n1608 ;
  assign n1610 = n331 | n416 ;
  assign n1611 = n245 | n861 ;
  assign n1612 = n1610 | n1611 ;
  assign n1613 = n1609 | n1612 ;
  assign n1614 = n486 | n928 ;
  assign n1615 = n214 | n306 ;
  assign n1616 = n455 | n1615 ;
  assign n1617 = n328 | n454 ;
  assign n1618 = n1616 | n1617 ;
  assign n1619 = n1614 | n1618 ;
  assign n1620 = n159 | n446 ;
  assign n1621 = n676 | n1123 ;
  assign n1622 = n1620 | n1621 ;
  assign n1623 = n1239 | n1622 ;
  assign n1624 = n1619 | n1623 ;
  assign n1625 = n1613 | n1624 ;
  assign n1626 = n256 | n434 ;
  assign n1627 = n110 | n1626 ;
  assign n1628 = n986 | n1627 ;
  assign n1629 = n899 | n1628 ;
  assign n1630 = n176 | n678 ;
  assign n1631 = n315 | n1630 ;
  assign n1632 = n1542 | n1631 ;
  assign n1633 = n1629 | n1632 ;
  assign n1634 = n606 | n1633 ;
  assign n1635 = n357 | n470 ;
  assign n1636 = n674 | n1635 ;
  assign n1637 = n80 | n302 ;
  assign n1638 = n149 | n667 ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = n1636 | n1639 ;
  assign n1641 = n1634 | n1640 ;
  assign n1642 = n184 | n835 ;
  assign n1643 = n508 | n1642 ;
  assign n1644 = n318 | n567 ;
  assign n1645 = n1643 | n1644 ;
  assign n1646 = n305 | n546 ;
  assign n1647 = n1447 | n1646 ;
  assign n1648 = n1645 | n1647 ;
  assign n1649 = n379 | n449 ;
  assign n1650 = n477 | n1649 ;
  assign n1651 = n346 | n734 ;
  assign n1652 = n1650 | n1651 ;
  assign n1653 = n103 | n1379 ;
  assign n1654 = n1652 | n1653 ;
  assign n1655 = n1648 | n1654 ;
  assign n1656 = n1641 | n1655 ;
  assign n1657 = n1625 | n1656 ;
  assign n1658 = n48 | n208 ;
  assign n1659 = n396 | n780 ;
  assign n1660 = n1658 | n1659 ;
  assign n1661 = n1040 | n1196 ;
  assign n1662 = n1660 | n1661 ;
  assign n1663 = n402 | n533 ;
  assign n1664 = n1294 | n1663 ;
  assign n1665 = n268 | n278 ;
  assign n1666 = n108 | n1048 ;
  assign n1667 = n1665 | n1666 ;
  assign n1668 = n1664 | n1667 ;
  assign n1669 = n1662 | n1668 ;
  assign n1670 = n244 | n407 ;
  assign n1671 = n700 | n1670 ;
  assign n1672 = n233 | n1332 ;
  assign n1673 = n983 | n1672 ;
  assign n1674 = n1671 | n1673 ;
  assign n1675 = n711 | n1119 ;
  assign n1676 = n1674 | n1675 ;
  assign n1677 = n193 | n751 ;
  assign n1678 = n221 | n1100 ;
  assign n1679 = n1677 | n1678 ;
  assign n1680 = n164 | n922 ;
  assign n1681 = n863 | n1680 ;
  assign n1682 = n345 | n362 ;
  assign n1683 = n1681 | n1682 ;
  assign n1684 = n1679 | n1683 ;
  assign n1685 = n1676 | n1684 ;
  assign n1686 = n1669 | n1685 ;
  assign n1687 = n1657 | n1686 ;
  assign n1688 = n329 | n464 ;
  assign n1689 = n141 | n378 ;
  assign n1690 = n528 | n1689 ;
  assign n1691 = n431 | n989 ;
  assign n1692 = n1690 | n1691 ;
  assign n1693 = n1688 | n1692 ;
  assign n1694 = n134 | n574 ;
  assign n1695 = n80 | n493 ;
  assign n1696 = n1694 | n1695 ;
  assign n1697 = n1693 | n1696 ;
  assign n1698 = n179 | n777 ;
  assign n1699 = n277 | n1698 ;
  assign n1700 = n899 | n1699 ;
  assign n1701 = n1697 | n1700 ;
  assign n1702 = n163 | n644 ;
  assign n1703 = n517 | n591 ;
  assign n1704 = n87 | n1703 ;
  assign n1705 = n189 | n1094 ;
  assign n1706 = n173 | n1705 ;
  assign n1707 = n1704 | n1706 ;
  assign n1708 = n1702 | n1707 ;
  assign n1709 = n1701 | n1708 ;
  assign n1710 = n524 | n616 ;
  assign n1711 = n265 | n321 ;
  assign n1712 = n1710 | n1711 ;
  assign n1713 = n214 | n964 ;
  assign n1714 = n70 | n1713 ;
  assign n1715 = n1712 | n1714 ;
  assign n1716 = n1439 | n1658 ;
  assign n1717 = n545 | n1074 ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = n1715 | n1718 ;
  assign n1720 = n226 | n656 ;
  assign n1721 = n165 | n342 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n256 | n338 ;
  assign n1724 = n197 | n1723 ;
  assign n1725 = n1533 | n1724 ;
  assign n1726 = n1722 | n1725 ;
  assign n1727 = n108 | n1351 ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = n1719 | n1728 ;
  assign n1730 = n1709 | n1729 ;
  assign n1731 = n103 | n113 ;
  assign n1732 = n434 | n1731 ;
  assign n1733 = n465 | n662 ;
  assign n1734 = n379 | n446 ;
  assign n1735 = n1733 | n1734 ;
  assign n1736 = n1732 | n1735 ;
  assign n1737 = n62 | n305 ;
  assign n1738 = n129 | n315 ;
  assign n1739 = n1737 | n1738 ;
  assign n1740 = n1736 | n1739 ;
  assign n1741 = n607 | n1148 ;
  assign n1742 = n296 | n442 ;
  assign n1743 = n262 | n1742 ;
  assign n1744 = n1741 | n1743 ;
  assign n1745 = n494 | n554 ;
  assign n1746 = n556 | n1745 ;
  assign n1747 = n403 | n1746 ;
  assign n1748 = n1744 | n1747 ;
  assign n1749 = n1740 | n1748 ;
  assign n1750 = n184 | n416 ;
  assign n1751 = n99 | n1081 ;
  assign n1752 = n1750 | n1751 ;
  assign n1753 = n1588 | n1752 ;
  assign n1754 = n1749 | n1753 ;
  assign n1755 = n480 | n557 ;
  assign n1756 = n546 | n1044 ;
  assign n1757 = n1755 | n1756 ;
  assign n1758 = n200 | n1757 ;
  assign n1759 = n356 | n1332 ;
  assign n1760 = n1758 | n1759 ;
  assign n1761 = n470 | n863 ;
  assign n1762 = n328 | n396 ;
  assign n1763 = n912 | n1762 ;
  assign n1764 = n1761 | n1763 ;
  assign n1765 = n1760 | n1764 ;
  assign n1766 = n412 | n1405 ;
  assign n1767 = n124 | n669 ;
  assign n1768 = n1766 | n1767 ;
  assign n1769 = n735 | n986 ;
  assign n1770 = n279 | n347 ;
  assign n1771 = n1769 | n1770 ;
  assign n1772 = n1768 | n1771 ;
  assign n1773 = n1765 | n1772 ;
  assign n1774 = n628 | n794 ;
  assign n1775 = n373 | n624 ;
  assign n1776 = n1774 | n1775 ;
  assign n1777 = n335 | n1020 ;
  assign n1778 = n176 | n1777 ;
  assign n1779 = n1776 | n1778 ;
  assign n1780 = n471 | n1069 ;
  assign n1781 = n318 | n1780 ;
  assign n1782 = n635 | n751 ;
  assign n1783 = n500 | n623 ;
  assign n1784 = n1782 | n1783 ;
  assign n1785 = n1781 | n1784 ;
  assign n1786 = n237 | n1006 ;
  assign n1787 = n1665 | n1786 ;
  assign n1788 = n1785 | n1787 ;
  assign n1789 = n1779 | n1788 ;
  assign n1790 = n1773 | n1789 ;
  assign n1791 = n1754 | n1790 ;
  assign n1792 = n1730 | n1791 ;
  assign n1793 = n373 | n493 ;
  assign n1794 = n374 | n644 ;
  assign n1795 = n268 | n780 ;
  assign n1796 = n1794 | n1795 ;
  assign n1797 = n1793 | n1796 ;
  assign n1798 = n1446 & ~n1797 ;
  assign n1799 = n44 & n171 ;
  assign n1800 = n1723 | n1799 ;
  assign n1801 = n1364 | n1800 ;
  assign n1802 = n587 | n1074 ;
  assign n1803 = n241 | n407 ;
  assign n1804 = n134 | n148 ;
  assign n1805 = n1803 | n1804 ;
  assign n1806 = n1802 | n1805 ;
  assign n1807 = n1801 | n1806 ;
  assign n1808 = n1798 & ~n1807 ;
  assign n1809 = n179 | n357 ;
  assign n1810 = n1782 | n1809 ;
  assign n1811 = n1484 | n1810 ;
  assign n1812 = n1808 & ~n1811 ;
  assign n1813 = n470 | n1332 ;
  assign n1814 = n1384 | n1813 ;
  assign n1815 = n1036 | n1814 ;
  assign n1816 = n372 | n611 ;
  assign n1817 = n176 | n405 ;
  assign n1818 = n1558 | n1817 ;
  assign n1819 = n643 | n1818 ;
  assign n1820 = n1816 | n1819 ;
  assign n1821 = n1815 | n1820 ;
  assign n1822 = n191 | n334 ;
  assign n1823 = n242 | n487 ;
  assign n1824 = n915 | n1823 ;
  assign n1825 = n220 | n1086 ;
  assign n1826 = n640 | n1825 ;
  assign n1827 = n1824 | n1826 ;
  assign n1828 = n1822 | n1827 ;
  assign n1829 = n1821 | n1828 ;
  assign n1830 = n1812 & ~n1829 ;
  assign n1831 = n488 | n1100 ;
  assign n1832 = n131 | n285 ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = n104 | n557 ;
  assign n1835 = n624 | n1834 ;
  assign n1836 = n1161 | n1835 ;
  assign n1837 = n1833 | n1836 ;
  assign n1838 = n1681 | n1837 ;
  assign n1839 = n1473 | n1838 ;
  assign n1840 = n1754 | n1839 ;
  assign n1841 = n1830 & ~n1840 ;
  assign n1842 = n86 | n428 ;
  assign n1843 = n200 | n497 ;
  assign n1844 = n913 | n1843 ;
  assign n1845 = n1842 | n1844 ;
  assign n1846 = n173 | n1193 ;
  assign n1847 = n1493 | n1846 ;
  assign n1848 = n1845 | n1847 ;
  assign n1849 = n688 | n777 ;
  assign n1850 = n1208 | n1429 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = n1848 | n1851 ;
  assign n1853 = n161 | n1688 ;
  assign n1854 = n148 | n586 ;
  assign n1855 = n864 | n1854 ;
  assign n1856 = n1853 | n1855 ;
  assign n1857 = n108 | n1020 ;
  assign n1858 = n1856 | n1857 ;
  assign n1859 = n125 | n314 ;
  assign n1860 = n306 | n781 ;
  assign n1861 = n1859 | n1860 ;
  assign n1862 = n378 | n667 ;
  assign n1863 = n1110 | n1862 ;
  assign n1864 = n1184 | n1863 ;
  assign n1865 = n1861 | n1864 ;
  assign n1866 = n1858 | n1865 ;
  assign n1867 = n1852 | n1866 ;
  assign n1868 = n742 | n1100 ;
  assign n1869 = n150 | n159 ;
  assign n1870 = n669 | n1869 ;
  assign n1871 = n1868 | n1870 ;
  assign n1872 = n345 | n405 ;
  assign n1873 = n662 | n1872 ;
  assign n1874 = n766 | n1873 ;
  assign n1875 = n1871 | n1874 ;
  assign n1876 = n260 | n1044 ;
  assign n1877 = n412 | n446 ;
  assign n1878 = n1876 | n1877 ;
  assign n1879 = n189 | n488 ;
  assign n1880 = n1878 | n1879 ;
  assign n1881 = n1134 | n1880 ;
  assign n1882 = n1875 | n1881 ;
  assign n1883 = n1867 | n1882 ;
  assign n1884 = n628 | n987 ;
  assign n1885 = n192 | n337 ;
  assign n1886 = n1884 | n1885 ;
  assign n1887 = n124 | n207 ;
  assign n1888 = n1886 | n1887 ;
  assign n1889 = n379 | n1745 ;
  assign n1890 = n174 | n256 ;
  assign n1891 = n342 | n1890 ;
  assign n1892 = n1889 | n1891 ;
  assign n1893 = n1888 | n1892 ;
  assign n1894 = n272 | n1893 ;
  assign n1895 = n278 | n477 ;
  assign n1896 = n393 | n1518 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = n165 | n356 ;
  assign n1899 = n55 | n700 ;
  assign n1900 = n1898 | n1899 ;
  assign n1901 = n1897 | n1900 ;
  assign n1902 = n1894 | n1901 ;
  assign n1903 = n734 | n772 ;
  assign n1904 = n372 | n712 ;
  assign n1905 = n1903 | n1904 ;
  assign n1906 = n261 | n1086 ;
  assign n1907 = n1905 | n1906 ;
  assign n1908 = n370 | n640 ;
  assign n1909 = n465 | n1908 ;
  assign n1910 = n613 | n647 ;
  assign n1911 = n308 | n1041 ;
  assign n1912 = n1910 | n1911 ;
  assign n1913 = n533 | n589 ;
  assign n1914 = n518 | n989 ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = n1912 | n1915 ;
  assign n1917 = n1909 | n1916 ;
  assign n1918 = n1907 | n1917 ;
  assign n1919 = n1902 | n1918 ;
  assign n1920 = n374 | n435 ;
  assign n1921 = n863 | n1920 ;
  assign n1922 = n1742 | n1921 ;
  assign n1923 = n656 | n750 ;
  assign n1924 = n83 | n1923 ;
  assign n1925 = n1922 | n1924 ;
  assign n1926 = n359 | n362 ;
  assign n1927 = n1702 | n1926 ;
  assign n1928 = n1925 | n1927 ;
  assign n1929 = n249 | n1928 ;
  assign n1930 = n1919 | n1929 ;
  assign n1931 = n1883 | n1930 ;
  assign n1932 = n441 | n534 ;
  assign n1933 = n525 | n1932 ;
  assign n1934 = n257 | n1933 ;
  assign n1935 = n454 | n1176 ;
  assign n1936 = n341 | n591 ;
  assign n1937 = n1935 | n1936 ;
  assign n1938 = n1934 | n1937 ;
  assign n1939 = n487 | n546 ;
  assign n1940 = n394 | n1939 ;
  assign n1941 = n1417 | n1940 ;
  assign n1942 = n1938 | n1941 ;
  assign n1943 = n1931 | n1942 ;
  assign n1944 = n1533 | n1745 ;
  assign n1945 = n1774 | n1944 ;
  assign n1946 = n131 | n500 ;
  assign n1947 = n1945 | n1946 ;
  assign n1948 = n90 | n96 ;
  assign n1949 = n448 | n1948 ;
  assign n1950 = n1947 | n1949 ;
  assign n1951 = n270 | n1414 ;
  assign n1952 = n454 | n1951 ;
  assign n1953 = n477 | n751 ;
  assign n1954 = n83 | n1953 ;
  assign n1955 = n347 | n614 ;
  assign n1956 = n1954 | n1955 ;
  assign n1957 = n989 | n1048 ;
  assign n1958 = n704 | n1957 ;
  assign n1959 = n1956 | n1958 ;
  assign n1960 = n1952 | n1959 ;
  assign n1961 = n1950 | n1960 ;
  assign n1962 = n302 | n1762 ;
  assign n1963 = n449 | n456 ;
  assign n1964 = n1962 | n1963 ;
  assign n1965 = n104 | n1822 ;
  assign n1966 = n777 | n1041 ;
  assign n1967 = n1817 | n1966 ;
  assign n1968 = n1965 | n1967 ;
  assign n1969 = n1964 | n1968 ;
  assign n1970 = n186 | n533 ;
  assign n1971 = n173 | n318 ;
  assign n1972 = n1970 | n1971 ;
  assign n1973 = n1969 | n1972 ;
  assign n1974 = n1961 | n1973 ;
  assign n1975 = n215 | n1012 ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = n147 | n232 ;
  assign n1978 = n433 | n1977 ;
  assign n1979 = n205 | n695 ;
  assign n1980 = n1058 | n1979 ;
  assign n1981 = n1978 | n1980 ;
  assign n1982 = n87 | n661 ;
  assign n1983 = n1094 | n1982 ;
  assign n1984 = n480 | n772 ;
  assign n1985 = n1983 | n1984 ;
  assign n1986 = n1981 | n1985 ;
  assign n1987 = n419 | n468 ;
  assign n1988 = n435 | n1987 ;
  assign n1989 = n864 | n1988 ;
  assign n1990 = n441 | n662 ;
  assign n1991 = n1171 | n1990 ;
  assign n1992 = n1989 | n1991 ;
  assign n1993 = n237 | n278 ;
  assign n1994 = n110 | n370 ;
  assign n1995 = n1993 | n1994 ;
  assign n1996 = n1992 | n1995 ;
  assign n1997 = n524 | n545 ;
  assign n1998 = n74 | n220 ;
  assign n1999 = n1997 | n1998 ;
  assign n2000 = n1092 | n1999 ;
  assign n2001 = n1996 | n2000 ;
  assign n2002 = n1986 | n2001 ;
  assign n2003 = n574 | n678 ;
  assign n2004 = n103 | n591 ;
  assign n2005 = n2003 | n2004 ;
  assign n2006 = n188 | n290 ;
  assign n2007 = n148 | n397 ;
  assign n2008 = n357 | n2007 ;
  assign n2009 = n2006 | n2008 ;
  assign n2010 = n226 | n667 ;
  assign n2011 = n284 | n2010 ;
  assign n2012 = n2009 | n2011 ;
  assign n2013 = n2005 | n2012 ;
  assign n2014 = n2002 | n2013 ;
  assign n2015 = n380 | n835 ;
  assign n2016 = n618 & ~n2015 ;
  assign n2017 = ~n987 & n2016 ;
  assign n2018 = n359 | n1193 ;
  assign n2019 = n550 | n586 ;
  assign n2020 = n1332 | n2019 ;
  assign n2021 = n2018 | n2020 ;
  assign n2022 = n1126 | n2021 ;
  assign n2023 = n2017 & ~n2022 ;
  assign n2024 = n546 | n647 ;
  assign n2025 = n1737 | n2024 ;
  assign n2026 = n275 | n999 ;
  assign n2027 = n48 | n2026 ;
  assign n2028 = n2025 | n2027 ;
  assign n2029 = n2023 & ~n2028 ;
  assign n2030 = n464 | n593 ;
  assign n2031 = n590 | n2030 ;
  assign n2032 = n429 | n2031 ;
  assign n2033 = n612 | n2032 ;
  assign n2034 = n372 | n640 ;
  assign n2035 = n323 | n528 ;
  assign n2036 = n2034 | n2035 ;
  assign n2037 = n1455 | n2036 ;
  assign n2038 = n2033 | n2037 ;
  assign n2039 = n2029 & ~n2038 ;
  assign n2040 = ~n2014 & n2039 ;
  assign n2041 = ~n1976 & n2040 ;
  assign n2042 = n140 | n555 ;
  assign n2043 = n449 | n1107 ;
  assign n2044 = n2042 | n2043 ;
  assign n2045 = n669 | n1048 ;
  assign n2046 = n396 | n968 ;
  assign n2047 = n2045 | n2046 ;
  assign n2048 = n2044 | n2047 ;
  assign n2049 = n1377 | n2048 ;
  assign n2050 = n605 | n1100 ;
  assign n2051 = n435 | n1044 ;
  assign n2052 = n293 | n518 ;
  assign n2053 = n756 | n2052 ;
  assign n2054 = n2051 | n2053 ;
  assign n2055 = n2050 | n2054 ;
  assign n2056 = n2049 | n2055 ;
  assign n2057 = n323 | n616 ;
  assign n2058 = n617 | n942 ;
  assign n2059 = n284 | n455 ;
  assign n2060 = n2058 | n2059 ;
  assign n2061 = n2057 | n2060 ;
  assign n2062 = n129 | n534 ;
  assign n2063 = n2024 | n2062 ;
  assign n2064 = n1257 | n1456 ;
  assign n2065 = n2063 | n2064 ;
  assign n2066 = n2061 | n2065 ;
  assign n2067 = n1055 | n1636 ;
  assign n2068 = n2066 | n2067 ;
  assign n2069 = n2056 | n2068 ;
  assign n2070 = n153 | n303 ;
  assign n2071 = n379 | n1123 ;
  assign n2072 = n772 | n841 ;
  assign n2073 = n2071 | n2072 ;
  assign n2074 = n338 | n545 ;
  assign n2075 = n2073 | n2074 ;
  assign n2076 = n2070 | n2075 ;
  assign n2077 = n2022 | n2076 ;
  assign n2078 = n346 | n372 ;
  assign n2079 = n431 | n567 ;
  assign n2080 = n2078 | n2079 ;
  assign n2081 = n471 | n707 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = n101 | n187 ;
  assign n2084 = ( n130 & n989 ) | ( n130 & n2083 ) | ( n989 & n2083 ) ;
  assign n2085 = n852 | n2084 ;
  assign n2086 = n2082 | n2085 ;
  assign n2087 = n46 & n121 ;
  assign n2088 = n488 | n2087 ;
  assign n2089 = n308 | n2088 ;
  assign n2090 = n1953 | n2089 ;
  assign n2091 = n2086 | n2090 ;
  assign n2092 = n141 | n734 ;
  assign n2093 = n1532 | n2092 ;
  assign n2094 = n493 | n794 ;
  assign n2095 = n715 | n2094 ;
  assign n2096 = n2093 | n2095 ;
  assign n2097 = n623 | n742 ;
  assign n2098 = n2096 | n2097 ;
  assign n2099 = n2091 | n2098 ;
  assign n2100 = n2077 | n2099 ;
  assign n2101 = n2069 | n2100 ;
  assign n2102 = n283 | n2101 ;
  assign n2103 = n214 | n574 ;
  assign n2104 = n617 | n2103 ;
  assign n2105 = n163 | n742 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n131 | n468 ;
  assign n2108 = n1659 | n2107 ;
  assign n2109 = n2106 | n2108 ;
  assign n2110 = n113 | n712 ;
  assign n2111 = n192 | n480 ;
  assign n2112 = n2110 | n2111 ;
  assign n2113 = n222 | n667 ;
  assign n2114 = n842 | n2113 ;
  assign n2115 = n2112 | n2114 ;
  assign n2116 = n2109 | n2115 ;
  assign n2117 = n1497 | n2116 ;
  assign n2118 = n405 | n1094 ;
  assign n2119 = n534 | n647 ;
  assign n2120 = n1041 | n1176 ;
  assign n2121 = n2119 | n2120 ;
  assign n2122 = n2118 | n2121 ;
  assign n2123 = n276 | n378 ;
  assign n2124 = n1253 | n2123 ;
  assign n2125 = n2122 | n2124 ;
  assign n2126 = n996 | n1504 ;
  assign n2127 = n2125 | n2126 ;
  assign n2128 = n589 | n914 ;
  assign n2129 = n2127 | n2128 ;
  assign n2130 = n2117 | n2129 ;
  assign n2131 = n306 | n471 ;
  assign n2132 = n1064 | n2131 ;
  assign n2133 = n497 | n1044 ;
  assign n2134 = n321 | n2133 ;
  assign n2135 = n2132 | n2134 ;
  assign n2136 = n941 | n1970 ;
  assign n2137 = n2135 | n2136 ;
  assign n2138 = n161 | n2087 ;
  assign n2139 = n526 | n2138 ;
  assign n2140 = n364 | n470 ;
  assign n2141 = n2139 | n2140 ;
  assign n2142 = n1520 | n2141 ;
  assign n2143 = n2137 | n2142 ;
  assign n2144 = n124 | n777 ;
  assign n2145 = n317 | n2144 ;
  assign n2146 = n108 | n129 ;
  assign n2147 = n643 | n2146 ;
  assign n2148 = n601 | n2147 ;
  assign n2149 = n2145 | n2148 ;
  assign n2150 = n540 | n1134 ;
  assign n2151 = n2149 | n2150 ;
  assign n2152 = n2143 | n2151 ;
  assign n2153 = n302 | n678 ;
  assign n2154 = n335 | n441 ;
  assign n2155 = n2153 | n2154 ;
  assign n2156 = n179 | n794 ;
  assign n2157 = n2155 | n2156 ;
  assign n2158 = n245 | n413 ;
  assign n2159 = n1196 | n2158 ;
  assign n2160 = n2157 | n2159 ;
  assign n2161 = n220 | n661 ;
  assign n2162 = n357 | n2161 ;
  assign n2163 = n435 | n2162 ;
  assign n2164 = n359 | n370 ;
  assign n2165 = n238 | n293 ;
  assign n2166 = n688 | n2165 ;
  assign n2167 = n2164 | n2166 ;
  assign n2168 = n2163 | n2167 ;
  assign n2169 = n2160 | n2168 ;
  assign n2170 = n314 | n442 ;
  assign n2171 = n339 | n2170 ;
  assign n2172 = n201 | n968 ;
  assign n2173 = n2171 | n2172 ;
  assign n2174 = n210 | n1100 ;
  assign n2175 = n586 | n628 ;
  assign n2176 = n48 | n2175 ;
  assign n2177 = n2174 | n2176 ;
  assign n2178 = n635 | n916 ;
  assign n2179 = n656 | n2178 ;
  assign n2180 = n178 | n328 ;
  assign n2181 = n428 | n2180 ;
  assign n2182 = n2179 | n2181 ;
  assign n2183 = n2177 | n2182 ;
  assign n2184 = n2173 | n2183 ;
  assign n2185 = n2169 | n2184 ;
  assign n2186 = n2152 | n2185 ;
  assign n2187 = n2130 | n2186 ;
  assign n2188 = n528 | n916 ;
  assign n2189 = n265 | n2188 ;
  assign n2190 = n346 | n547 ;
  assign n2191 = n2189 | n2190 ;
  assign n2192 = n1475 | n2191 ;
  assign n2193 = n712 | n2058 ;
  assign n2194 = n2192 | n2193 ;
  assign n2195 = n97 | n261 ;
  assign n2196 = n150 | n2195 ;
  assign n2197 = n357 | n456 ;
  assign n2198 = n1672 | n2197 ;
  assign n2199 = n2196 | n2198 ;
  assign n2200 = n2194 | n2199 ;
  assign n2201 = n220 | n322 ;
  assign n2202 = n368 | n2201 ;
  assign n2203 = n1569 | n2202 ;
  assign n2204 = n545 | n860 ;
  assign n2205 = n628 | n2204 ;
  assign n2206 = n471 | n688 ;
  assign n2207 = n123 | n2206 ;
  assign n2208 = n2205 | n2207 ;
  assign n2209 = n2203 | n2208 ;
  assign n2210 = n161 | n468 ;
  assign n2211 = n449 | n1086 ;
  assign n2212 = n151 | n2211 ;
  assign n2213 = n2210 | n2212 ;
  assign n2214 = n134 | n465 ;
  assign n2215 = n1494 | n2214 ;
  assign n2216 = ~n557 & n618 ;
  assign n2217 = ~n2215 & n2216 ;
  assign n2218 = ~n2213 & n2217 ;
  assign n2219 = ~n2209 & n2218 ;
  assign n2220 = ~n771 & n2219 ;
  assign n2221 = ~n2200 & n2220 ;
  assign n2222 = n241 | n329 ;
  assign n2223 = n485 | n614 ;
  assign n2224 = n679 | n2223 ;
  assign n2225 = n1720 | n2224 ;
  assign n2226 = n729 | n1895 ;
  assign n2227 = n2070 | n2226 ;
  assign n2228 = n2225 | n2227 ;
  assign n2229 = n2222 | n2228 ;
  assign n2230 = n2221 & ~n2229 ;
  assign n2231 = n611 | n1095 ;
  assign n2232 = n336 | n1594 ;
  assign n2233 = n2231 | n2232 ;
  assign n2234 = n406 | n587 ;
  assign n2235 = n1437 | n2234 ;
  assign n2236 = n2233 | n2235 ;
  assign n2237 = n82 | n260 ;
  assign n2238 = n535 | n2237 ;
  assign n2239 = n1340 | n2238 ;
  assign n2240 = n2236 | n2239 ;
  assign n2241 = n331 | n431 ;
  assign n2242 = n70 | n835 ;
  assign n2243 = n661 | n2242 ;
  assign n2244 = n1074 | n2243 ;
  assign n2245 = n2241 | n2244 ;
  assign n2246 = n275 | n317 ;
  assign n2247 = n640 | n2246 ;
  assign n2248 = n314 | n2247 ;
  assign n2249 = n360 | n455 ;
  assign n2250 = n219 | n2249 ;
  assign n2251 = n2248 | n2250 ;
  assign n2252 = n2245 | n2251 ;
  assign n2253 = n2240 | n2252 ;
  assign n2254 = n2230 & ~n2253 ;
  assign n2255 = n315 | n566 ;
  assign n2256 = n208 | n210 ;
  assign n2257 = n2255 | n2256 ;
  assign n2258 = n88 & n797 ;
  assign n2259 = n144 | n2258 ;
  assign n2260 = n1045 | n2259 ;
  assign n2261 = n2257 | n2260 ;
  assign n2262 = n2005 | n2261 ;
  assign n2263 = n55 | n378 ;
  assign n2264 = n351 | n442 ;
  assign n2265 = n2263 | n2264 ;
  assign n2266 = n405 | n416 ;
  assign n2267 = n2158 | n2266 ;
  assign n2268 = n2265 | n2267 ;
  assign n2269 = n173 | n363 ;
  assign n2270 = n305 | n623 ;
  assign n2271 = n419 | n526 ;
  assign n2272 = n2270 | n2271 ;
  assign n2273 = n2269 | n2272 ;
  assign n2274 = n2268 | n2273 ;
  assign n2275 = n2262 | n2274 ;
  assign n2276 = n131 | n750 ;
  assign n2277 = n396 | n446 ;
  assign n2278 = n2276 | n2277 ;
  assign n2279 = n74 | n987 ;
  assign n2280 = n2278 | n2279 ;
  assign n2281 = n2275 | n2280 ;
  assign n2282 = n2254 & ~n2281 ;
  assign n2283 = n618 & ~n1193 ;
  assign n2284 = ~n1224 & n2283 ;
  assign n2285 = n723 | n1044 ;
  assign n2286 = n2284 & ~n2285 ;
  assign n2287 = ~n1609 & n2286 ;
  assign n2288 = n667 | n781 ;
  assign n2289 = n198 | n567 ;
  assign n2290 = n123 | n2289 ;
  assign n2291 = n2288 | n2290 ;
  assign n2292 = n341 | n526 ;
  assign n2293 = n134 | n269 ;
  assign n2294 = n2292 | n2293 ;
  assign n2295 = n1058 | n2294 ;
  assign n2296 = n2291 | n2295 ;
  assign n2297 = n2287 & ~n2296 ;
  assign n2298 = n201 | n1042 ;
  assign n2299 = n404 | n722 ;
  assign n2300 = n2298 | n2299 ;
  assign n2301 = n2297 & ~n2300 ;
  assign n2302 = n605 | n2118 ;
  assign n2303 = n161 | n163 ;
  assign n2304 = n264 | n392 ;
  assign n2305 = n2303 | n2304 ;
  assign n2306 = n2302 | n2305 ;
  assign n2307 = n1048 | n1074 ;
  assign n2308 = n1110 | n2307 ;
  assign n2309 = n2306 | n2308 ;
  assign n2310 = n260 | n591 ;
  assign n2311 = n500 | n624 ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = n164 | n480 ;
  assign n2314 = n2312 | n2313 ;
  assign n2315 = n2309 | n2314 ;
  assign n2316 = n1543 | n1627 ;
  assign n2317 = n551 | n1126 ;
  assign n2318 = n2316 | n2317 ;
  assign n2319 = n1017 | n2318 ;
  assign n2320 = n2315 | n2319 ;
  assign n2321 = n185 | n412 ;
  assign n2322 = n2241 | n2321 ;
  assign n2323 = n189 | n285 ;
  assign n2324 = n315 | n2323 ;
  assign n2325 = n467 | n2324 ;
  assign n2326 = n2322 | n2325 ;
  assign n2327 = n1533 | n1913 ;
  assign n2328 = n105 | n2327 ;
  assign n2329 = n2326 | n2328 ;
  assign n2330 = n2320 | n2329 ;
  assign n2331 = n2301 & ~n2330 ;
  assign n2332 = n329 | n468 ;
  assign n2333 = n200 | n488 ;
  assign n2334 = n2263 | n2333 ;
  assign n2335 = n2332 | n2334 ;
  assign n2336 = n254 | n546 ;
  assign n2337 = n347 | n613 ;
  assign n2338 = n2336 | n2337 ;
  assign n2339 = n2335 | n2338 ;
  assign n2340 = n946 | n2205 ;
  assign n2341 = n2339 | n2340 ;
  assign n2342 = n360 | n373 ;
  assign n2343 = n80 | n454 ;
  assign n2344 = n2342 | n2343 ;
  assign n2345 = n427 | n2344 ;
  assign n2346 = n147 | n179 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = n640 | n704 ;
  assign n2349 = n1302 | n2348 ;
  assign n2350 = n1413 | n2349 ;
  assign n2351 = n173 | n380 ;
  assign n2352 = n270 | n2351 ;
  assign n2353 = n2350 | n2352 ;
  assign n2354 = n2347 | n2353 ;
  assign n2355 = n2341 | n2354 ;
  assign n2356 = n788 | n956 ;
  assign n2357 = n153 | n244 ;
  assign n2358 = n586 | n1113 ;
  assign n2359 = n2357 | n2358 ;
  assign n2360 = n2356 | n2359 ;
  assign n2361 = n2355 | n2360 ;
  assign n2362 = n215 | n337 ;
  assign n2363 = n2361 | n2362 ;
  assign n2364 = n2331 & ~n2363 ;
  assign n2365 = n1625 | n1919 ;
  assign n2366 = n133 | n517 ;
  assign n2367 = n153 | n2366 ;
  assign n2368 = n814 | n2207 ;
  assign n2369 = n2367 | n2368 ;
  assign n2370 = n1837 | n2369 ;
  assign n2371 = n87 | n1876 ;
  assign n2372 = n1955 | n2371 ;
  assign n2373 = n574 | n1020 ;
  assign n2374 = n319 | n2373 ;
  assign n2375 = n2372 | n2374 ;
  assign n2376 = n2370 | n2375 ;
  assign n2377 = n161 | n321 ;
  assign n2378 = n134 | n279 ;
  assign n2379 = n2377 | n2378 ;
  assign n2380 = n188 | n1392 ;
  assign n2381 = n413 | n432 ;
  assign n2382 = n2380 | n2381 ;
  assign n2383 = n2379 | n2382 ;
  assign n2384 = n679 | n1094 ;
  assign n2385 = n148 | n707 ;
  assign n2386 = n2384 | n2385 ;
  assign n2387 = n468 | n942 ;
  assign n2388 = n141 | n2387 ;
  assign n2389 = n2386 | n2388 ;
  assign n2390 = n185 | n303 ;
  assign n2391 = n616 | n2390 ;
  assign n2392 = n373 | n440 ;
  assign n2393 = n1659 | n2392 ;
  assign n2394 = n2391 | n2393 ;
  assign n2395 = n2389 | n2394 ;
  assign n2396 = n2383 | n2395 ;
  assign n2397 = n2376 | n2396 ;
  assign n2398 = n2365 | n2397 ;
  assign n2399 = n392 | n517 ;
  assign n2400 = n705 | n2399 ;
  assign n2401 = n328 | n413 ;
  assign n2402 = n435 | n534 ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = n2400 | n2403 ;
  assign n2405 = n104 | n254 ;
  assign n2406 = n308 | n2405 ;
  assign n2407 = n404 | n1193 ;
  assign n2408 = n2406 | n2407 ;
  assign n2409 = n2404 | n2408 ;
  assign n2410 = n983 | n1357 ;
  assign n2411 = n2409 | n2410 ;
  assign n2412 = n545 | n600 ;
  assign n2413 = n256 | n586 ;
  assign n2414 = n265 | n2413 ;
  assign n2415 = n2412 | n2414 ;
  assign n2416 = n707 | n1006 ;
  assign n2417 = n290 | n1069 ;
  assign n2418 = n2416 | n2417 ;
  assign n2419 = n2415 | n2418 ;
  assign n2420 = n82 | n546 ;
  assign n2421 = n90 | n1862 ;
  assign n2422 = n2420 | n2421 ;
  assign n2423 = n842 | n1593 ;
  assign n2424 = n2422 | n2423 ;
  assign n2425 = n2419 | n2424 ;
  assign n2426 = n2411 | n2425 ;
  assign n2427 = n849 | n1533 ;
  assign n2428 = n222 | n777 ;
  assign n2429 = n627 | n2428 ;
  assign n2430 = n2427 | n2429 ;
  assign n2431 = n133 | n689 ;
  assign n2432 = n1793 | n2431 ;
  assign n2433 = n989 | n2432 ;
  assign n2434 = n253 | n296 ;
  assign n2435 = n2433 | n2434 ;
  assign n2436 = n2430 | n2435 ;
  assign n2437 = n2426 | n2436 ;
  assign n2438 = n225 | n233 ;
  assign n2439 = n816 | n2438 ;
  assign n2440 = n285 | n674 ;
  assign n2441 = n1649 | n2440 ;
  assign n2442 = n338 | n1332 ;
  assign n2443 = n515 & ~n2442 ;
  assign n2444 = ~n915 & n2443 ;
  assign n2445 = ~n2441 & n2444 ;
  assign n2446 = ~n2439 & n2445 ;
  assign n2447 = n148 | n1176 ;
  assign n2448 = n635 | n2447 ;
  assign n2449 = n362 | n835 ;
  assign n2450 = n2448 | n2449 ;
  assign n2451 = n276 | n465 ;
  assign n2452 = n659 | n2451 ;
  assign n2453 = n2450 | n2452 ;
  assign n2454 = n2446 & ~n2453 ;
  assign n2455 = n186 | n1317 ;
  assign n2456 = n1560 | n2455 ;
  assign n2457 = ~n238 & n618 ;
  assign n2458 = ~n1620 & n2457 ;
  assign n2459 = ~n2456 & n2458 ;
  assign n2460 = n214 | n500 ;
  assign n2461 = n295 | n2460 ;
  assign n2462 = n1257 | n2461 ;
  assign n2463 = n2459 & ~n2462 ;
  assign n2464 = n2454 & n2463 ;
  assign n2465 = ~n2437 & n2464 ;
  assign n2466 = n100 | n761 ;
  assign n2467 = n2465 & ~n2466 ;
  assign n2468 = n1895 | n2189 ;
  assign n2469 = n2203 | n2468 ;
  assign n2470 = n201 | n915 ;
  assign n2471 = n2469 | n2470 ;
  assign n2472 = n233 | n655 ;
  assign n2473 = n488 | n2472 ;
  assign n2474 = n1007 | n2473 ;
  assign n2475 = n269 | n345 ;
  assign n2476 = n1309 | n2475 ;
  assign n2477 = n2474 | n2476 ;
  assign n2478 = n485 | n863 ;
  assign n2479 = n140 | n487 ;
  assign n2480 = n2478 | n2479 ;
  assign n2481 = n270 | n1041 ;
  assign n2482 = n900 | n2481 ;
  assign n2483 = n2480 | n2482 ;
  assign n2484 = n2477 | n2483 ;
  assign n2485 = n2471 | n2484 ;
  assign n2486 = n2152 | n2485 ;
  assign n2487 = n80 | n1332 ;
  assign n2488 = n151 | n2487 ;
  assign n2489 = n2367 | n2488 ;
  assign n2490 = n62 | n624 ;
  assign n2491 = n2489 | n2490 ;
  assign n2492 = n464 | n554 ;
  assign n2493 = n226 | n290 ;
  assign n2494 = n2492 | n2493 ;
  assign n2495 = n824 | n2494 ;
  assign n2496 = n1194 | n1462 ;
  assign n2497 = n2495 | n2496 ;
  assign n2498 = n2491 | n2497 ;
  assign n2499 = n618 & ~n1157 ;
  assign n2500 = ~n1658 & n2499 ;
  assign n2501 = ~n834 & n2500 ;
  assign n2502 = n302 | n772 ;
  assign n2503 = n408 | n881 ;
  assign n2504 = n2502 | n2503 ;
  assign n2505 = n1793 | n2402 ;
  assign n2506 = n164 | n613 ;
  assign n2507 = n2505 | n2506 ;
  assign n2508 = n2504 | n2507 ;
  assign n2509 = n2501 & ~n2508 ;
  assign n2510 = n674 | n795 ;
  assign n2511 = n318 | n518 ;
  assign n2512 = n2510 | n2511 ;
  assign n2513 = n277 | n2512 ;
  assign n2514 = n188 | n237 ;
  assign n2515 = n2288 | n2514 ;
  assign n2516 = n197 | n200 ;
  assign n2517 = n2515 | n2516 ;
  assign n2518 = n2513 | n2517 ;
  assign n2519 = n2509 & ~n2518 ;
  assign n2520 = ~n2498 & n2519 ;
  assign n2521 = ~n2486 & n2520 ;
  assign n2522 = n1018 | n1317 ;
  assign n2523 = n892 | n1601 ;
  assign n2524 = n2522 | n2523 ;
  assign n2525 = n600 | n2524 ;
  assign n2526 = n164 | n623 ;
  assign n2527 = n1962 | n2526 ;
  assign n2528 = n174 | n1069 ;
  assign n2529 = n1737 | n2528 ;
  assign n2530 = n2527 | n2529 ;
  assign n2531 = n2525 | n2530 ;
  assign n2532 = n432 | n850 ;
  assign n2533 = n742 | n2532 ;
  assign n2534 = n477 | n1126 ;
  assign n2535 = n2533 | n2534 ;
  assign n2536 = n446 | n678 ;
  assign n2537 = n356 | n2536 ;
  assign n2538 = n2535 | n2537 ;
  assign n2539 = n161 | n440 ;
  assign n2540 = n319 | n2539 ;
  assign n2541 = n2104 | n2540 ;
  assign n2542 = n2538 | n2541 ;
  assign n2543 = n2531 | n2542 ;
  assign n2544 = n103 | n176 ;
  assign n2545 = n1064 | n2544 ;
  assign n2546 = n322 | n586 ;
  assign n2547 = n262 | n2546 ;
  assign n2548 = n2545 | n2547 ;
  assign n2549 = n87 | n198 ;
  assign n2550 = n148 | n253 ;
  assign n2551 = n2549 | n2550 ;
  assign n2552 = n407 | n435 ;
  assign n2553 = ~n454 & n618 ;
  assign n2554 = ~n2552 & n2553 ;
  assign n2555 = ~n1178 & n2554 ;
  assign n2556 = ~n2551 & n2555 ;
  assign n2557 = ~n2548 & n2556 ;
  assign n2558 = n659 | n1086 ;
  assign n2559 = n795 | n2558 ;
  assign n2560 = n1254 | n2559 ;
  assign n2561 = n206 | n238 ;
  assign n2562 = n2206 | n2561 ;
  assign n2563 = n2560 | n2562 ;
  assign n2564 = n2557 & ~n2563 ;
  assign n2565 = n365 | n1874 ;
  assign n2566 = n488 | n493 ;
  assign n2567 = n113 | n1074 ;
  assign n2568 = n2566 | n2567 ;
  assign n2569 = n2565 | n2568 ;
  assign n2570 = n2564 & ~n2569 ;
  assign n2571 = ~n2543 & n2570 ;
  assign n2572 = n323 | n441 ;
  assign n2573 = n243 | n2572 ;
  assign n2574 = n707 | n946 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = n110 | n245 ;
  assign n2577 = n279 | n628 ;
  assign n2578 = n2576 | n2577 ;
  assign n2579 = n70 | n232 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = n2575 | n2580 ;
  assign n2582 = n467 | n1572 ;
  assign n2583 = n404 | n733 ;
  assign n2584 = n207 | n220 ;
  assign n2585 = n1756 | n2584 ;
  assign n2586 = n2583 | n2585 ;
  assign n2587 = n2582 | n2586 ;
  assign n2588 = n2581 | n2587 ;
  assign n2589 = n276 | n689 ;
  assign n2590 = n578 | n2589 ;
  assign n2591 = n1409 | n1420 ;
  assign n2592 = n373 | n534 ;
  assign n2593 = n2591 | n2592 ;
  assign n2594 = n2590 | n2593 ;
  assign n2595 = n44 & n120 ;
  assign n2596 = n667 | n2595 ;
  assign n2597 = n1843 | n2596 ;
  assign n2598 = n824 | n2597 ;
  assign n2599 = n2594 | n2598 ;
  assign n2600 = n2588 | n2599 ;
  assign n2601 = n347 | n567 ;
  assign n2602 = n419 | n679 ;
  assign n2603 = n80 | n104 ;
  assign n2604 = n2602 | n2603 ;
  assign n2605 = n401 | n2604 ;
  assign n2606 = n2601 | n2605 ;
  assign n2607 = n2600 | n2606 ;
  assign n2608 = n2571 & ~n2607 ;
  assign n2609 = n486 | n1439 ;
  assign n2610 = n403 | n2609 ;
  assign n2611 = n322 | n1100 ;
  assign n2612 = n189 | n361 ;
  assign n2613 = n2611 | n2612 ;
  assign n2614 = n2610 | n2613 ;
  assign n2615 = n750 | n2131 ;
  assign n2616 = n2379 | n2615 ;
  assign n2617 = n1523 | n2616 ;
  assign n2618 = n2614 | n2617 ;
  assign n2619 = n253 | n337 ;
  assign n2620 = n351 | n2188 ;
  assign n2621 = n960 | n2620 ;
  assign n2622 = n2619 | n2621 ;
  assign n2623 = n1014 | n1253 ;
  assign n2624 = n1876 | n2623 ;
  assign n2625 = n1354 | n2624 ;
  assign n2626 = n2622 | n2625 ;
  assign n2627 = n2618 | n2626 ;
  assign n2628 = n192 | n221 ;
  assign n2629 = n374 | n493 ;
  assign n2630 = n1755 | n2629 ;
  assign n2631 = n2628 | n2630 ;
  assign n2632 = n380 | n677 ;
  assign n2633 = n314 | n2632 ;
  assign n2634 = n2631 | n2633 ;
  assign n2635 = n1907 | n2634 ;
  assign n2636 = n362 | n1069 ;
  assign n2637 = n578 | n2636 ;
  assign n2638 = n2025 | n2389 ;
  assign n2639 = n2637 | n2638 ;
  assign n2640 = n2635 | n2639 ;
  assign n2641 = n2627 | n2640 ;
  assign n2642 = n1976 | n2641 ;
  assign n2643 = n264 | n787 ;
  assign n2644 = n480 | n497 ;
  assign n2645 = n408 | n2644 ;
  assign n2646 = n2643 | n2645 ;
  assign n2647 = n188 | n345 ;
  assign n2648 = n147 | n342 ;
  assign n2649 = n2647 | n2648 ;
  assign n2650 = n447 | n2649 ;
  assign n2651 = n131 | n165 ;
  assign n2652 = n265 | n2651 ;
  assign n2653 = n434 | n704 ;
  assign n2654 = n2652 | n2653 ;
  assign n2655 = n2650 | n2654 ;
  assign n2656 = n2646 | n2655 ;
  assign n2657 = n707 | n1294 ;
  assign n2658 = n220 | n441 ;
  assign n2659 = n110 | n2658 ;
  assign n2660 = n1178 | n2659 ;
  assign n2661 = n2657 | n2660 ;
  assign n2662 = n2656 | n2661 ;
  assign n2663 = n129 | n751 ;
  assign n2664 = n99 | n245 ;
  assign n2665 = n2663 | n2664 ;
  assign n2666 = n70 | n378 ;
  assign n2667 = n2665 | n2666 ;
  assign n2668 = n1094 | n2667 ;
  assign n2669 = n2637 | n2668 ;
  assign n2670 = n184 | n734 ;
  assign n2671 = n2051 | n2670 ;
  assign n2672 = n1113 | n2671 ;
  assign n2673 = n2669 | n2672 ;
  assign n2674 = n428 | n1299 ;
  assign n2675 = n369 | n756 ;
  assign n2676 = n2674 | n2675 ;
  assign n2677 = n574 | n1723 ;
  assign n2678 = n233 | n2677 ;
  assign n2679 = n807 | n2678 ;
  assign n2680 = n2676 | n2679 ;
  assign n2681 = n2673 | n2680 ;
  assign n2682 = n2662 | n2681 ;
  assign n2683 = n189 | n780 ;
  assign n2684 = n341 | n412 ;
  assign n2685 = n2683 | n2684 ;
  assign n2686 = n1485 | n2685 ;
  assign n2687 = n431 | n2686 ;
  assign n2688 = n1145 | n2448 ;
  assign n2689 = n2687 | n2688 ;
  assign n2690 = n290 | n464 ;
  assign n2691 = n419 | n689 ;
  assign n2692 = n134 | n2691 ;
  assign n2693 = n494 | n999 ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = n2690 | n2694 ;
  assign n2696 = n358 | n1783 ;
  assign n2697 = n207 | n613 ;
  assign n2698 = n334 | n600 ;
  assign n2699 = n2697 | n2698 ;
  assign n2700 = n2696 | n2699 ;
  assign n2701 = n1407 | n2700 ;
  assign n2702 = n2695 | n2701 ;
  assign n2703 = n2689 | n2702 ;
  assign n2704 = n103 | n440 ;
  assign n2705 = n359 | n2704 ;
  assign n2706 = n679 | n922 ;
  assign n2707 = n296 | n554 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = n2705 | n2708 ;
  assign n2710 = n174 | n214 ;
  assign n2711 = n380 | n2710 ;
  assign n2712 = n2549 | n2711 ;
  assign n2713 = n2709 | n2712 ;
  assign n2714 = n1779 | n2713 ;
  assign n2715 = n254 | n667 ;
  assign n2716 = n315 | n350 ;
  assign n2717 = n2715 | n2716 ;
  assign n2718 = n2238 | n2717 ;
  assign n2719 = n374 | n1538 ;
  assign n2720 = n2718 | n2719 ;
  assign n2721 = n2714 | n2720 ;
  assign n2722 = n2703 | n2721 ;
  assign n2723 = n2682 | n2722 ;
  assign n2724 = n567 | n1392 ;
  assign n2725 = n392 | n449 ;
  assign n2726 = n2332 | n2725 ;
  assign n2727 = n2724 | n2726 ;
  assign n2728 = n74 | n153 ;
  assign n2729 = n221 | n912 ;
  assign n2730 = n48 | n2729 ;
  assign n2731 = n2728 | n2730 ;
  assign n2732 = n2727 | n2731 ;
  assign n2733 = n1557 | n2732 ;
  assign n2734 = n1871 | n2733 ;
  assign n2735 = n2723 | n2734 ;
  assign n2736 = n788 | n1462 ;
  assign n2737 = n427 | n2333 ;
  assign n2738 = n2736 | n2737 ;
  assign n2739 = n862 | n2738 ;
  assign n2740 = n303 | n528 ;
  assign n2741 = n269 | n294 ;
  assign n2742 = n2740 | n2741 ;
  assign n2743 = n1192 | n2742 ;
  assign n2744 = n245 | n545 ;
  assign n2745 = n1702 | n2744 ;
  assign n2746 = n2743 | n2745 ;
  assign n2747 = n2739 | n2746 ;
  assign n2748 = n165 | n835 ;
  assign n2749 = n97 | n624 ;
  assign n2750 = n2748 | n2749 ;
  assign n2751 = n2006 | n2750 ;
  assign n2752 = n677 | n916 ;
  assign n2753 = n1086 | n2752 ;
  assign n2754 = n222 | n287 ;
  assign n2755 = n2753 | n2754 ;
  assign n2756 = n2751 | n2755 ;
  assign n2757 = n2747 | n2756 ;
  assign n2758 = n314 | n1332 ;
  assign n2759 = n2270 | n2758 ;
  assign n2760 = n144 | n464 ;
  assign n2761 = n2759 | n2760 ;
  assign n2762 = n334 | n662 ;
  assign n2763 = n2119 | n2762 ;
  assign n2764 = n2440 | n2763 ;
  assign n2765 = n550 | n656 ;
  assign n2766 = n1083 | n2765 ;
  assign n2767 = n147 | n749 ;
  assign n2768 = n2766 | n2767 ;
  assign n2769 = n2764 | n2768 ;
  assign n2770 = n2761 | n2769 ;
  assign n2771 = n2757 | n2770 ;
  assign n2772 = n432 | n628 ;
  assign n2773 = n220 | n2772 ;
  assign n2774 = n176 | n1006 ;
  assign n2775 = n589 | n2774 ;
  assign n2776 = n2773 | n2775 ;
  assign n2777 = n350 | n1795 ;
  assign n2778 = n1380 | n2777 ;
  assign n2779 = n2776 | n2778 ;
  assign n2780 = n62 | n1533 ;
  assign n2781 = n208 | n471 ;
  assign n2782 = n447 | n2781 ;
  assign n2783 = n2780 | n2782 ;
  assign n2784 = n2779 | n2783 ;
  assign n2785 = n129 | n494 ;
  assign n2786 = n526 | n2785 ;
  assign n2787 = n345 | n419 ;
  assign n2788 = n2786 | n2787 ;
  assign n2789 = n359 | n407 ;
  assign n2790 = n2401 | n2789 ;
  assign n2791 = n2788 | n2790 ;
  assign n2792 = n372 | n953 ;
  assign n2793 = n635 | n723 ;
  assign n2794 = n2792 | n2793 ;
  assign n2795 = n2628 | n2794 ;
  assign n2796 = n2791 | n2795 ;
  assign n2797 = n2784 | n2796 ;
  assign n2798 = n2771 | n2797 ;
  assign n2799 = n700 | n2057 ;
  assign n2800 = n1732 | n2799 ;
  assign n2801 = n296 | n772 ;
  assign n2802 = n669 | n2801 ;
  assign n2803 = n1423 | n2802 ;
  assign n2804 = n2800 | n2803 ;
  assign n2805 = n781 | n2619 ;
  assign n2806 = n2804 | n2805 ;
  assign n2807 = n733 | n975 ;
  assign n2808 = n179 | n1126 ;
  assign n2809 = n276 | n2808 ;
  assign n2810 = n2807 | n2809 ;
  assign n2811 = n1113 | n1615 ;
  assign n2812 = n2210 | n2811 ;
  assign n2813 = n2810 | n2812 ;
  assign n2814 = n267 | n1426 ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = n2806 | n2815 ;
  assign n2817 = ( x24 & n613 ) | ( x24 & n1499 ) | ( n613 & n1499 ) ;
  assign n2818 = n1952 | n2817 ;
  assign n2819 = n2816 | n2818 ;
  assign n2820 = n2798 | n2819 ;
  assign n2821 = n210 | n780 ;
  assign n2822 = n160 | n2821 ;
  assign n2823 = n1876 | n2822 ;
  assign n2824 = n659 | n2823 ;
  assign n2825 = n98 & n263 ;
  assign n2826 = n841 | n2825 ;
  assign n2827 = n2824 | n2826 ;
  assign n2828 = n125 | n2131 ;
  assign n2829 = n285 | n442 ;
  assign n2830 = n2492 | n2829 ;
  assign n2831 = n1089 | n2830 ;
  assign n2832 = n2828 | n2831 ;
  assign n2833 = n2827 | n2832 ;
  assign n2834 = n363 | n677 ;
  assign n2835 = n2833 | n2834 ;
  assign n2836 = n712 | n1086 ;
  assign n2837 = n215 | n695 ;
  assign n2838 = n2836 | n2837 ;
  assign n2839 = n1048 | n1332 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n188 | n480 ;
  assign n2842 = n618 & ~n674 ;
  assign n2843 = ~n2841 & n2842 ;
  assign n2844 = ~n2840 & n2843 ;
  assign n2845 = n691 | n1732 ;
  assign n2846 = n2844 & ~n2845 ;
  assign n2847 = ~n2835 & n2846 ;
  assign n2848 = ~n2043 & n2847 ;
  assign n2849 = ~n2485 & n2848 ;
  assign n2850 = n574 | n635 ;
  assign n2851 = n835 | n2850 ;
  assign n2852 = n2078 | n2851 ;
  assign n2853 = n287 | n401 ;
  assign n2854 = n860 | n1020 ;
  assign n2855 = n2853 | n2854 ;
  assign n2856 = n96 | n734 ;
  assign n2857 = n1351 | n2856 ;
  assign n2858 = n2855 | n2857 ;
  assign n2859 = n2412 | n2858 ;
  assign n2860 = n2581 | n2859 ;
  assign n2861 = n2852 | n2860 ;
  assign n2862 = n331 | n762 ;
  assign n2863 = n238 | n1081 ;
  assign n2864 = n2862 | n2863 ;
  assign n2865 = n1035 | n2864 ;
  assign n2866 = n87 | n124 ;
  assign n2867 = n968 | n2866 ;
  assign n2868 = n2865 | n2867 ;
  assign n2869 = n2861 | n2868 ;
  assign n2870 = n640 | n669 ;
  assign n2871 = n1170 | n2870 ;
  assign n2872 = n341 | n751 ;
  assign n2873 = n2059 | n2872 ;
  assign n2874 = n2871 | n2873 ;
  assign n2875 = n468 | n613 ;
  assign n2876 = n535 | n2875 ;
  assign n2877 = n62 | n2019 ;
  assign n2878 = n2876 | n2877 ;
  assign n2879 = n2874 | n2878 ;
  assign n2880 = n360 | n556 ;
  assign n2881 = n133 | n2880 ;
  assign n2882 = n1926 | n2881 ;
  assign n2883 = n431 | n526 ;
  assign n2884 = n319 | n2883 ;
  assign n2885 = n2882 | n2884 ;
  assign n2886 = n2879 | n2885 ;
  assign n2887 = n2869 | n2886 ;
  assign n2888 = n2849 & ~n2887 ;
  assign n2889 = n153 | n1040 ;
  assign n2890 = n533 | n863 ;
  assign n2891 = n2697 | n2890 ;
  assign n2892 = n2889 | n2891 ;
  assign n2893 = n808 | n1106 ;
  assign n2894 = n2892 | n2893 ;
  assign n2895 = n253 | n1074 ;
  assign n2896 = n722 | n2895 ;
  assign n2897 = n124 | n591 ;
  assign n2898 = n942 | n2897 ;
  assign n2899 = n2896 | n2898 ;
  assign n2900 = n2894 | n2899 ;
  assign n2901 = n173 | n756 ;
  assign n2902 = n1006 | n2901 ;
  assign n2903 = n2900 | n2902 ;
  assign n2904 = n1549 | n2903 ;
  assign n2905 = n2847 & ~n2904 ;
  assign n2906 = n408 | n2684 ;
  assign n2907 = n2399 | n2906 ;
  assign n2908 = n201 | n334 ;
  assign n2909 = n316 | n2908 ;
  assign n2910 = n2907 | n2909 ;
  assign n2911 = n502 | n2910 ;
  assign n2912 = n440 | n485 ;
  assign n2913 = n351 | n2912 ;
  assign n2914 = n189 | n369 ;
  assign n2915 = n372 | n2914 ;
  assign n2916 = n2913 | n2915 ;
  assign n2917 = n144 | n176 ;
  assign n2918 = n55 | n715 ;
  assign n2919 = n2917 | n2918 ;
  assign n2920 = n2748 | n2919 ;
  assign n2921 = n2916 | n2920 ;
  assign n2922 = n413 | n600 ;
  assign n2923 = n1133 | n2922 ;
  assign n2924 = n2921 | n2923 ;
  assign n2925 = n1168 | n2924 ;
  assign n2926 = n2911 | n2925 ;
  assign n2927 = n99 | n707 ;
  assign n2928 = n338 | n2927 ;
  assign n2929 = n1698 | n2928 ;
  assign n2930 = n781 | n1069 ;
  assign n2931 = n2420 | n2930 ;
  assign n2932 = n2929 | n2931 ;
  assign n2933 = n416 | n1176 ;
  assign n2934 = n1831 | n2933 ;
  assign n2935 = n48 | n1041 ;
  assign n2936 = n1533 | n2935 ;
  assign n2937 = n2934 | n2936 ;
  assign n2938 = n2932 | n2937 ;
  assign n2939 = n1178 | n1542 ;
  assign n2940 = n357 | n572 ;
  assign n2941 = n2939 | n2940 ;
  assign n2942 = n2938 | n2941 ;
  assign n2943 = n2926 | n2942 ;
  assign n2944 = n2905 & ~n2943 ;
  assign n2945 = n916 | n968 ;
  assign n2946 = n214 | n689 ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = n74 | n1374 ;
  assign n2949 = n2947 | n2948 ;
  assign n2950 = n147 | n1006 ;
  assign n2951 = n660 | n2950 ;
  assign n2952 = n2949 | n2951 ;
  assign n2953 = n1391 | n2024 ;
  assign n2954 = n234 | n2953 ;
  assign n2955 = n623 | n999 ;
  assign n2956 = n392 | n850 ;
  assign n2957 = n2955 | n2956 ;
  assign n2958 = n2954 | n2957 ;
  assign n2959 = n2952 | n2958 ;
  assign n2960 = n1812 & ~n2959 ;
  assign n2961 = n191 | n912 ;
  assign n2962 = n2611 | n2961 ;
  assign n2963 = n254 | n734 ;
  assign n2964 = n160 | n2963 ;
  assign n2965 = n2828 | n2964 ;
  assign n2966 = n2962 | n2965 ;
  assign n2967 = n200 | n456 ;
  assign n2968 = n1378 | n2539 ;
  assign n2969 = n2967 | n2968 ;
  assign n2970 = n2966 | n2969 ;
  assign n2971 = n265 | n431 ;
  assign n2972 = n2487 | n2971 ;
  assign n2973 = n319 | n488 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = n2970 | n2974 ;
  assign n2976 = n1433 | n2975 ;
  assign n2977 = n2960 & ~n2976 ;
  assign n2978 = n396 | n1006 ;
  assign n2979 = n321 | n2978 ;
  assign n2980 = n222 | n485 ;
  assign n2981 = n2979 | n2980 ;
  assign n2982 = n322 | n455 ;
  assign n2983 = n197 | n2982 ;
  assign n2984 = n2981 | n2983 ;
  assign n2985 = n1986 | n2984 ;
  assign n2986 = n1637 | n2145 ;
  assign n2987 = n2265 | n2986 ;
  assign n2988 = n176 | n268 ;
  assign n2989 = n144 | n1074 ;
  assign n2990 = n2988 | n2989 ;
  assign n2991 = n1419 | n1586 ;
  assign n2992 = n2990 | n2991 ;
  assign n2993 = n2987 | n2992 ;
  assign n2994 = n2985 | n2993 ;
  assign n2995 = n715 | n750 ;
  assign n2996 = n269 | n794 ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = n316 | n2997 ;
  assign n2999 = n173 | n308 ;
  assign n3000 = n220 | n624 ;
  assign n3001 = n885 | n3000 ;
  assign n3002 = n2999 | n3001 ;
  assign n3003 = n2998 | n3002 ;
  assign n3004 = n362 | n379 ;
  assign n3005 = n2119 | n3004 ;
  assign n3006 = n3003 | n3005 ;
  assign n3007 = n192 | n707 ;
  assign n3008 = n330 | n704 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = n689 | n3009 ;
  assign n3011 = n338 | n1041 ;
  assign n3012 = n1793 | n3011 ;
  assign n3013 = n848 | n2908 ;
  assign n3014 = n3012 | n3013 ;
  assign n3015 = n3010 | n3014 ;
  assign n3016 = n518 | n860 ;
  assign n3017 = n191 | n3016 ;
  assign n3018 = n2321 | n3017 ;
  assign n3019 = n2800 | n3018 ;
  assign n3020 = n3015 | n3019 ;
  assign n3021 = n253 | n487 ;
  assign n3022 = n150 | n2683 ;
  assign n3023 = n3021 | n3022 ;
  assign n3024 = n360 | n497 ;
  assign n3025 = n675 | n3024 ;
  assign n3026 = n640 | n912 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = n3023 | n3027 ;
  assign n3029 = n3020 | n3028 ;
  assign n3030 = n3006 | n3029 ;
  assign n3031 = n2994 | n3030 ;
  assign n3032 = n161 | n915 ;
  assign n3033 = n556 | n751 ;
  assign n3034 = n3032 | n3033 ;
  assign n3035 = n356 | n2601 ;
  assign n3036 = n3034 | n3035 ;
  assign n3037 = n237 | n428 ;
  assign n3038 = n588 | n3037 ;
  assign n3039 = n3036 | n3038 ;
  assign n3040 = n179 | n285 ;
  assign n3041 = n1550 | n3040 ;
  assign n3042 = n1713 | n3041 ;
  assign n3043 = n2017 & ~n3042 ;
  assign n3044 = ~n3039 & n3043 ;
  assign n3045 = n1013 | n1425 ;
  assign n3046 = n1646 | n3045 ;
  assign n3047 = n2791 | n3046 ;
  assign n3048 = n3044 & ~n3047 ;
  assign n3049 = ~n3031 & n3048 ;
  assign n3050 = n97 | n350 ;
  assign n3051 = n1953 | n3050 ;
  assign n3052 = n88 & n507 ;
  assign n3053 = n3051 | n3052 ;
  assign n3054 = n260 | n734 ;
  assign n3055 = n556 | n1086 ;
  assign n3056 = n3054 | n3055 ;
  assign n3057 = n2050 | n3056 ;
  assign n3058 = n3053 | n3057 ;
  assign n3059 = n108 | n380 ;
  assign n3060 = n178 | n3059 ;
  assign n3061 = n131 | n226 ;
  assign n3062 = n3060 | n3061 ;
  assign n3063 = n1761 | n2058 ;
  assign n3064 = n3062 | n3063 ;
  assign n3065 = n408 | n2967 ;
  assign n3066 = n3064 | n3065 ;
  assign n3067 = n3058 | n3066 ;
  assign n3068 = n293 | n723 ;
  assign n3069 = n48 | n917 ;
  assign n3070 = n3068 | n3069 ;
  assign n3071 = n104 | n153 ;
  assign n3072 = n208 | n1069 ;
  assign n3073 = n3071 | n3072 ;
  assign n3074 = n3070 | n3073 ;
  assign n3075 = n3067 | n3074 ;
  assign n3076 = n133 | n659 ;
  assign n3077 = n1338 | n3076 ;
  assign n3078 = n342 | n374 ;
  assign n3079 = n574 | n3078 ;
  assign n3080 = n163 | n488 ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = n221 | n435 ;
  assign n3083 = n160 | n3082 ;
  assign n3084 = n3081 | n3083 ;
  assign n3085 = n3077 | n3084 ;
  assign n3086 = n3075 | n3085 ;
  assign n3087 = n2994 | n3086 ;
  assign n3088 = n1926 | n2042 ;
  assign n3089 = n2298 | n3088 ;
  assign n3090 = n198 | n712 ;
  assign n3091 = ~x25 & n59 ;
  assign n3092 = n58 & n3091 ;
  assign n3093 = n3090 | n3092 ;
  assign n3094 = n789 | n3093 ;
  assign n3095 = n1064 | n1923 ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = n3089 | n3096 ;
  assign n3098 = n422 | n662 ;
  assign n3099 = n151 | n3098 ;
  assign n3100 = n238 | n497 ;
  assign n3101 = n534 | n667 ;
  assign n3102 = n3100 | n3101 ;
  assign n3103 = n3099 | n3102 ;
  assign n3104 = n763 | n3037 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = n253 | n368 ;
  assign n3107 = n669 | n3106 ;
  assign n3108 = n3105 | n3107 ;
  assign n3109 = n3097 | n3108 ;
  assign n3110 = n2441 | n2758 ;
  assign n3111 = n90 | n601 ;
  assign n3112 = n1816 | n3111 ;
  assign n3113 = n3110 | n3112 ;
  assign n3114 = n225 | n287 ;
  assign n3115 = n427 | n3114 ;
  assign n3116 = n74 | n493 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = n679 | n781 ;
  assign n3119 = n356 | n3118 ;
  assign n3120 = n3117 | n3119 ;
  assign n3121 = n3113 | n3120 ;
  assign n3122 = n3109 | n3121 ;
  assign n3123 = n3087 | n3122 ;
  assign n3124 = ~n3049 & n3123 ;
  assign n3125 = n2977 & ~n3124 ;
  assign n3126 = n2944 | n3125 ;
  assign n3127 = n2888 & n3126 ;
  assign n3128 = n2820 & ~n3127 ;
  assign n3129 = n2735 | n3128 ;
  assign n3130 = n2642 & n3129 ;
  assign n3131 = n2608 & ~n3130 ;
  assign n3132 = n2521 | n3131 ;
  assign n3133 = n2467 & n3132 ;
  assign n3134 = n2398 & ~n3133 ;
  assign n3135 = n2364 & ~n3134 ;
  assign n3136 = n2282 | n3135 ;
  assign n3137 = ~n2187 & n3136 ;
  assign n3138 = n2102 & ~n3137 ;
  assign n3139 = n2041 & ~n3138 ;
  assign n3140 = n1943 & ~n3139 ;
  assign n3141 = n1841 & ~n3140 ;
  assign n3142 = n1792 & ~n3141 ;
  assign n3143 = n1687 | n3142 ;
  assign n3144 = n1600 & n3143 ;
  assign n3145 = n1529 & ~n3144 ;
  assign n3146 = n1398 & ~n3145 ;
  assign n3147 = n1316 | n3146 ;
  assign n3148 = ~n1207 & n3147 ;
  assign n3149 = n1118 & ~n3148 ;
  assign n3150 = n995 & ~n3149 ;
  assign n3151 = n859 | n3150 ;
  assign n3152 = ~n721 & n3151 ;
  assign n3153 = n293 | n407 ;
  assign n3154 = n578 | n3153 ;
  assign n3155 = n557 | n589 ;
  assign n3156 = n174 | n269 ;
  assign n3157 = n3155 | n3156 ;
  assign n3158 = n3154 | n3157 ;
  assign n3159 = n1470 | n3158 ;
  assign n3160 = ~n517 & n618 ;
  assign n3161 = ~n2658 & n3160 ;
  assign n3162 = ~n3159 & n3161 ;
  assign n3163 = n286 | n844 ;
  assign n3164 = n1045 | n3163 ;
  assign n3165 = n705 | n3164 ;
  assign n3166 = n842 | n2222 ;
  assign n3167 = n294 | n545 ;
  assign n3168 = n2263 | n3167 ;
  assign n3169 = n3166 | n3168 ;
  assign n3170 = n3165 | n3169 ;
  assign n3171 = n3162 & ~n3170 ;
  assign n3172 = n2164 | n2514 ;
  assign n3173 = n186 | n659 ;
  assign n3174 = n2895 | n3173 ;
  assign n3175 = n3172 | n3174 ;
  assign n3176 = n1069 | n1550 ;
  assign n3177 = n1616 | n3176 ;
  assign n3178 = n3175 | n3177 ;
  assign n3179 = n3171 & ~n3178 ;
  assign n3180 = n89 | n695 ;
  assign n3181 = n1267 | n3180 ;
  assign n3182 = n1217 | n3181 ;
  assign n3183 = n83 | n2690 ;
  assign n3184 = n3182 | n3183 ;
  assign n3185 = n337 | n679 ;
  assign n3186 = n983 | n3185 ;
  assign n3187 = n757 | n3186 ;
  assign n3188 = n3184 | n3187 ;
  assign n3189 = n700 | n794 ;
  assign n3190 = n661 | n3189 ;
  assign n3191 = n1486 | n3190 ;
  assign n3192 = n524 | n1048 ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = n404 | n1005 ;
  assign n3195 = n322 | n342 ;
  assign n3196 = n2180 | n3195 ;
  assign n3197 = n1380 | n3196 ;
  assign n3198 = n3194 | n3197 ;
  assign n3199 = n3193 | n3198 ;
  assign n3200 = n3188 | n3199 ;
  assign n3201 = n3179 & ~n3200 ;
  assign n3202 = n201 | n2416 ;
  assign n3203 = n1399 | n3202 ;
  assign n3204 = n611 | n3203 ;
  assign n3205 = n360 | n624 ;
  assign n3206 = n242 | n850 ;
  assign n3207 = n3205 | n3206 ;
  assign n3208 = n527 | n3207 ;
  assign n3209 = n3204 | n3208 ;
  assign n3210 = n198 | n303 ;
  assign n3211 = n1737 | n3210 ;
  assign n3212 = n3209 | n3211 ;
  assign n3213 = n111 | n207 ;
  assign n3214 = n3004 | n3213 ;
  assign n3215 = n2438 | n2704 ;
  assign n3216 = n1849 | n3215 ;
  assign n3217 = n3214 | n3216 ;
  assign n3218 = n917 | n1224 ;
  assign n3219 = n3217 | n3218 ;
  assign n3220 = n163 | n313 ;
  assign n3221 = n419 | n546 ;
  assign n3222 = n3220 | n3221 ;
  assign n3223 = n351 | n470 ;
  assign n3224 = n1302 | n1777 ;
  assign n3225 = n3223 | n3224 ;
  assign n3226 = n3222 | n3225 ;
  assign n3227 = n3219 | n3226 ;
  assign n3228 = n3212 | n3227 ;
  assign n3229 = n465 | n712 ;
  assign n3230 = n2852 | n3229 ;
  assign n3231 = n3228 | n3230 ;
  assign n3232 = n3201 & ~n3231 ;
  assign n3233 = ~n3049 & n3232 ;
  assign n3234 = ~n3123 & n3233 ;
  assign n3235 = ( n3049 & ~n3123 ) | ( n3049 & n3234 ) | ( ~n3123 & n3234 ) ;
  assign n3236 = n2977 | n3235 ;
  assign n3237 = n2944 & n3236 ;
  assign n3238 = n2888 | n3237 ;
  assign n3239 = ~n2820 & n3238 ;
  assign n3240 = n2735 & ~n3239 ;
  assign n3241 = n2642 | n3240 ;
  assign n3242 = ~n2608 & n3241 ;
  assign n3243 = n2521 & ~n3242 ;
  assign n3244 = n2467 | n3243 ;
  assign n3245 = ~n2364 & n2398 ;
  assign n3246 = ( n2364 & n3244 ) | ( n2364 & ~n3245 ) | ( n3244 & ~n3245 ) ;
  assign n3247 = n2282 & n3246 ;
  assign n3248 = n2187 & ~n3247 ;
  assign n3249 = n2102 | n3248 ;
  assign n3250 = ~n2041 & n3249 ;
  assign n3251 = n1943 | n3250 ;
  assign n3252 = ~n1841 & n3251 ;
  assign n3253 = n1687 & n1792 ;
  assign n3254 = ( n1687 & n3252 ) | ( n1687 & n3253 ) | ( n3252 & n3253 ) ;
  assign n3255 = n1600 | n3254 ;
  assign n3256 = ~n1529 & n3255 ;
  assign n3257 = n1398 | n3256 ;
  assign n3258 = n1316 & n3257 ;
  assign n3259 = n1207 & ~n3258 ;
  assign n3260 = n1118 | n3259 ;
  assign n3261 = ~n995 & n3260 ;
  assign n3262 = n859 & ~n3261 ;
  assign n3263 = n721 & ~n3262 ;
  assign n3264 = n564 & ~n3263 ;
  assign n3265 = ~n3152 & n3264 ;
  assign n3266 = n564 | n3152 ;
  assign n3267 = n3263 | n3266 ;
  assign n3268 = ( ~n564 & n3265 ) | ( ~n564 & n3267 ) | ( n3265 & n3267 ) ;
  assign n3269 = n390 & ~n3268 ;
  assign n3270 = ~x31 & n389 ;
  assign n3271 = n564 & n3270 ;
  assign n3272 = x31 & ~n66 ;
  assign n3273 = x31 & n49 ;
  assign n3274 = ( n49 & n3272 ) | ( n49 & ~n3273 ) | ( n3272 & ~n3273 ) ;
  assign n3275 = ~n721 & n3274 ;
  assign n3276 = n3271 | n3275 ;
  assign n3277 = n859 & n3273 ;
  assign n3278 = n3276 | n3277 ;
  assign n3279 = n3269 | n3278 ;
  assign n3280 = n370 | n647 ;
  assign n3281 = n133 | n256 ;
  assign n3282 = n218 | n3281 ;
  assign n3283 = n3280 | n3282 ;
  assign n3284 = n331 | n3283 ;
  assign n3285 = n80 | n412 ;
  assign n3286 = n2636 | n3285 ;
  assign n3287 = n3284 | n3286 ;
  assign n3288 = n182 | n1769 ;
  assign n3289 = n3287 | n3288 ;
  assign n3290 = n113 | n528 ;
  assign n3291 = n124 | n432 ;
  assign n3292 = n3290 | n3291 ;
  assign n3293 = n244 | n347 ;
  assign n3294 = n3292 | n3293 ;
  assign n3295 = n103 | n593 ;
  assign n3296 = n220 | n3295 ;
  assign n3297 = n2725 | n3026 ;
  assign n3298 = n3296 | n3297 ;
  assign n3299 = n3294 | n3298 ;
  assign n3300 = n3289 | n3299 ;
  assign n3301 = n522 | n851 ;
  assign n3302 = n1221 | n3301 ;
  assign n3303 = n480 | n550 ;
  assign n3304 = ~n85 & n251 ;
  assign n3305 = n275 | n3304 ;
  assign n3306 = n3303 | n3305 ;
  assign n3307 = n3302 | n3306 ;
  assign n3308 = n2204 | n2377 ;
  assign n3309 = n3307 | n3308 ;
  assign n3310 = n3300 | n3309 ;
  assign n3311 = n210 | n915 ;
  assign n3312 = n987 | n3311 ;
  assign n3313 = n546 | n662 ;
  assign n3314 = n2611 | n3313 ;
  assign n3315 = n3312 | n3314 ;
  assign n3316 = n1876 | n2057 ;
  assign n3317 = n508 | n3316 ;
  assign n3318 = n3315 | n3317 ;
  assign n3319 = n276 | n485 ;
  assign n3320 = n605 | n3319 ;
  assign n3321 = n1210 | n3320 ;
  assign n3322 = n3318 | n3321 ;
  assign n3323 = n524 | n841 ;
  assign n3324 = n2664 | n3323 ;
  assign n3325 = n715 | n989 ;
  assign n3326 = n3324 | n3325 ;
  assign n3327 = n850 | n1006 ;
  assign n3328 = n493 | n3327 ;
  assign n3329 = n3326 | n3328 ;
  assign n3330 = n3322 | n3329 ;
  assign n3331 = n3310 | n3330 ;
  assign n3332 = n122 | n574 ;
  assign n3333 = n1202 | n3052 ;
  assign n3334 = n3332 | n3333 ;
  assign n3335 = n74 | n125 ;
  assign n3336 = n342 | n591 ;
  assign n3337 = n82 | n3336 ;
  assign n3338 = n3335 | n3337 ;
  assign n3339 = n3334 | n3338 ;
  assign n3340 = n625 | n3339 ;
  assign n3341 = n1396 | n3340 ;
  assign n3342 = n3331 | n3341 ;
  assign n3343 = ( ~n388 & n3279 ) | ( ~n388 & n3342 ) | ( n3279 & n3342 ) ;
  assign n3344 = n315 | n545 ;
  assign n3345 = n2132 | n3344 ;
  assign n3346 = n257 | n863 ;
  assign n3347 = n244 | n261 ;
  assign n3348 = n3346 | n3347 ;
  assign n3349 = n3345 | n3348 ;
  assign n3350 = n323 | n695 ;
  assign n3351 = n318 | n3350 ;
  assign n3352 = n1199 | n1257 ;
  assign n3353 = n3351 | n3352 ;
  assign n3354 = n271 | n3353 ;
  assign n3355 = n302 | n517 ;
  assign n3356 = n1809 | n3355 ;
  assign n3357 = n2867 | n3356 ;
  assign n3358 = n3354 | n3357 ;
  assign n3359 = n3349 | n3358 ;
  assign n3360 = n613 | n662 ;
  assign n3361 = n317 | n1822 ;
  assign n3362 = n3360 | n3361 ;
  assign n3363 = n788 | n1250 ;
  assign n3364 = n3362 | n3363 ;
  assign n3365 = n129 | n860 ;
  assign n3366 = n147 | n554 ;
  assign n3367 = n3365 | n3366 ;
  assign n3368 = n70 | n667 ;
  assign n3369 = n294 | n3368 ;
  assign n3370 = n3367 | n3369 ;
  assign n3371 = n3364 | n3370 ;
  assign n3372 = n3359 | n3371 ;
  assign n3373 = n192 | n1081 ;
  assign n3374 = n141 | n174 ;
  assign n3375 = n600 | n3374 ;
  assign n3376 = n3373 | n3375 ;
  assign n3377 = n780 | n989 ;
  assign n3378 = n586 | n3377 ;
  assign n3379 = n120 & n130 ;
  assign n3380 = n647 | n3379 ;
  assign n3381 = n3378 | n3380 ;
  assign n3382 = n3376 | n3381 ;
  assign n3383 = n854 | n1184 ;
  assign n3384 = n345 | n678 ;
  assign n3385 = n380 | n435 ;
  assign n3386 = n3384 | n3385 ;
  assign n3387 = n2030 | n3386 ;
  assign n3388 = n3383 | n3387 ;
  assign n3389 = n3382 | n3388 ;
  assign n3390 = n245 | n392 ;
  assign n3391 = n2107 | n3390 ;
  assign n3392 = n3173 | n3391 ;
  assign n3393 = n442 | n1029 ;
  assign n3394 = n3392 | n3393 ;
  assign n3395 = n477 | n715 ;
  assign n3396 = n1998 | n3395 ;
  assign n3397 = n3394 | n3396 ;
  assign n3398 = n3389 | n3397 ;
  assign n3399 = n3372 | n3398 ;
  assign n3400 = n3231 | n3399 ;
  assign n3401 = ( x26 & n388 ) | ( x26 & n3400 ) | ( n388 & n3400 ) ;
  assign n3402 = ( ~x26 & n388 ) | ( ~x26 & n3400 ) | ( n388 & n3400 ) ;
  assign n3403 = ( x26 & ~n3401 ) | ( x26 & n3402 ) | ( ~n3401 & n3402 ) ;
  assign n3404 = n564 & n3274 ;
  assign n3405 = ~n721 & n3273 ;
  assign n3406 = n3404 | n3405 ;
  assign n3407 = n390 | n3406 ;
  assign n3408 = ( n60 & n2083 ) | ( n60 & ~n3091 ) | ( n2083 & ~n3091 ) ;
  assign n3409 = ( n142 & n337 ) | ( n142 & n3408 ) | ( n337 & n3408 ) ;
  assign n3410 = n1193 | n3409 ;
  assign n3411 = n44 | n121 ;
  assign n3412 = ~n777 & n3411 ;
  assign n3413 = n3410 | n3412 ;
  assign n3414 = n163 | n3413 ;
  assign n3415 = n220 | n527 ;
  assign n3416 = n3414 | n3415 ;
  assign n3417 = n112 | n435 ;
  assign n3418 = ( n435 & ~n3416 ) | ( n435 & n3417 ) | ( ~n3416 & n3417 ) ;
  assign n3419 = n184 | n3418 ;
  assign n3420 = n269 | n346 ;
  assign n3421 = n416 | n3420 ;
  assign n3422 = n1301 | n3421 ;
  assign n3423 = n2260 | n3422 ;
  assign n3424 = n486 | n711 ;
  assign n3425 = n214 | n715 ;
  assign n3426 = n2765 | n3425 ;
  assign n3427 = n108 | n287 ;
  assign n3428 = n2333 | n3427 ;
  assign n3429 = n3426 | n3428 ;
  assign n3430 = n3424 | n3429 ;
  assign n3431 = n254 | n357 ;
  assign n3432 = n218 | n3431 ;
  assign n3433 = n305 | n379 ;
  assign n3434 = n3432 | n3433 ;
  assign n3435 = n3430 | n3434 ;
  assign n3436 = n3423 | n3435 ;
  assign n3437 = n635 | n780 ;
  assign n3438 = n134 | n3437 ;
  assign n3439 = n260 | n647 ;
  assign n3440 = n3438 | n3439 ;
  assign n3441 = n1236 | n3440 ;
  assign n3442 = n1069 | n1444 ;
  assign n3443 = n3441 | n3442 ;
  assign n3444 = n3436 | n3443 ;
  assign n3445 = n233 | n742 ;
  assign n3446 = n557 | n661 ;
  assign n3447 = n3445 | n3446 ;
  assign n3448 = n141 | n293 ;
  assign n3449 = n2982 | n3448 ;
  assign n3450 = n315 | n468 ;
  assign n3451 = n3449 | n3450 ;
  assign n3452 = n3447 | n3451 ;
  assign n3453 = n62 | n294 ;
  assign n3454 = n153 | n222 ;
  assign n3455 = n3453 | n3454 ;
  assign n3456 = n246 | n851 ;
  assign n3457 = n3455 | n3456 ;
  assign n3458 = n3452 | n3457 ;
  assign n3459 = n270 | n337 ;
  assign n3460 = n3033 | n3459 ;
  assign n3461 = n3458 | n3460 ;
  assign n3462 = n3444 | n3461 ;
  assign n3463 = n160 | n313 ;
  assign n3464 = n2644 | n3463 ;
  assign n3465 = n777 | n987 ;
  assign n3466 = n2602 | n3465 ;
  assign n3467 = n3464 | n3466 ;
  assign n3468 = n677 | n835 ;
  assign n3469 = n3021 | n3468 ;
  assign n3470 = n3467 | n3469 ;
  assign n3471 = n401 | n794 ;
  assign n3472 = n241 | n3471 ;
  assign n3473 = n527 | n1302 ;
  assign n3474 = n3472 | n3473 ;
  assign n3475 = n317 | n942 ;
  assign n3476 = n3474 | n3475 ;
  assign n3477 = n1723 | n3476 ;
  assign n3478 = n3470 | n3477 ;
  assign n3479 = n1100 | n1630 ;
  assign n3480 = n210 | n2087 ;
  assign n3481 = n618 & ~n3480 ;
  assign n3482 = ~n3479 & n3481 ;
  assign n3483 = ~n3478 & n3482 ;
  assign n3484 = n237 | n408 ;
  assign n3485 = n3483 & ~n3484 ;
  assign n3486 = ~n3462 & n3485 ;
  assign n3487 = ~n3419 & n3486 ;
  assign n3488 = n3266 & ~n3487 ;
  assign n3489 = ~n3264 & n3266 ;
  assign n3490 = n3487 & ~n3489 ;
  assign n3491 = n3264 & ~n3487 ;
  assign n3492 = ( n3488 & n3490 ) | ( n3488 & ~n3491 ) | ( n3490 & ~n3491 ) ;
  assign n3493 = ( n3406 & n3407 ) | ( n3406 & ~n3492 ) | ( n3407 & ~n3492 ) ;
  assign n3494 = n3270 & ~n3487 ;
  assign n3495 = n3493 | n3494 ;
  assign n3496 = ( n3343 & ~n3403 ) | ( n3343 & n3495 ) | ( ~n3403 & n3495 ) ;
  assign n3497 = n50 | n56 ;
  assign n3498 = x26 & x27 ;
  assign n3499 = ~x26 & x27 ;
  assign n3500 = ( x26 & ~n3498 ) | ( x26 & n3499 ) | ( ~n3498 & n3499 ) ;
  assign n3501 = n3497 & ~n3500 ;
  assign n3502 = n85 & ~n521 ;
  assign n3503 = ~n345 & n3502 ;
  assign n3504 = n1044 | n1630 ;
  assign n3505 = n2762 | n3504 ;
  assign n3506 = n94 | n751 ;
  assign n3507 = n1100 | n3506 ;
  assign n3508 = n70 | n589 ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = n3505 | n3509 ;
  assign n3511 = ( n45 & ~n72 ) | ( n45 & n506 ) | ( ~n72 & n506 ) ;
  assign n3512 = ( n67 & n535 ) | ( n67 & n3511 ) | ( n535 & n3511 ) ;
  assign n3513 = n3510 | n3512 ;
  assign n3514 = n220 | n3513 ;
  assign n3515 = n3410 | n3514 ;
  assign n3516 = n3503 & ~n3515 ;
  assign n3517 = n3501 & ~n3516 ;
  assign n3518 = x29 & n3517 ;
  assign n3519 = n581 | n1414 ;
  assign n3520 = n58 | n276 ;
  assign n3521 = n2144 | n3520 ;
  assign n3522 = n77 | n128 ;
  assign n3523 = n3521 | n3522 ;
  assign n3524 = ~n71 & n3522 ;
  assign n3525 = ( n3519 & n3523 ) | ( n3519 & ~n3524 ) | ( n3523 & ~n3524 ) ;
  assign n3526 = n2680 | n3525 ;
  assign n3527 = n88 | n2646 ;
  assign n3528 = n74 | n3527 ;
  assign n3529 = n3526 | n3528 ;
  assign n3530 = n3411 | n3529 ;
  assign n3531 = n163 | n1193 ;
  assign n3532 = n3503 & ~n3531 ;
  assign n3533 = ~n3530 & n3532 ;
  assign n3534 = x26 | n43 ;
  assign n3535 = x26 | x29 ;
  assign n3536 = ( n158 & ~n3534 ) | ( n158 & n3535 ) | ( ~n3534 & n3535 ) ;
  assign n3537 = ~n3533 & n3536 ;
  assign n3538 = x28 & x29 ;
  assign n3539 = x28 | x29 ;
  assign n3540 = ~n3538 & n3539 ;
  assign n3541 = n3500 & n3540 ;
  assign n3542 = n3537 | n3541 ;
  assign n3543 = n236 & n506 ;
  assign n3544 = n725 | n3543 ;
  assign n3545 = n3290 | n3544 ;
  assign n3546 = n160 | n357 ;
  assign n3547 = n455 | n1086 ;
  assign n3548 = n3189 | n3547 ;
  assign n3549 = n3546 | n3548 ;
  assign n3550 = n3545 | n3549 ;
  assign n3551 = n270 | n1392 ;
  assign n3552 = n3550 | n3551 ;
  assign n3553 = n3419 | n3552 ;
  assign n3554 = n3443 | n3553 ;
  assign n3555 = n51 & ~n77 ;
  assign n3556 = n1083 | n3555 ;
  assign n3557 = n1389 | n3556 ;
  assign n3558 = ~n493 & n515 ;
  assign n3559 = ~n3557 & n3558 ;
  assign n3560 = n188 | n593 ;
  assign n3561 = n148 | n613 ;
  assign n3562 = n3560 | n3561 ;
  assign n3563 = n296 | n335 ;
  assign n3564 = n207 | n471 ;
  assign n3565 = n3563 | n3564 ;
  assign n3566 = n3562 | n3565 ;
  assign n3567 = n3559 & ~n3566 ;
  assign n3568 = n129 | n341 ;
  assign n3569 = n1019 | n3568 ;
  assign n3570 = n844 | n3569 ;
  assign n3571 = n466 | n518 ;
  assign n3572 = n3570 | n3571 ;
  assign n3573 = n580 | n3572 ;
  assign n3574 = n3567 & ~n3573 ;
  assign n3575 = n2601 | n2955 ;
  assign n3576 = n3010 | n3575 ;
  assign n3577 = n103 | n3206 ;
  assign n3578 = n1862 | n3577 ;
  assign n3579 = n3576 | n3578 ;
  assign n3580 = n3574 & ~n3579 ;
  assign n3581 = n659 | n2856 ;
  assign n3582 = n3479 | n3581 ;
  assign n3583 = n549 | n3582 ;
  assign n3584 = n3527 | n3583 ;
  assign n3585 = n3580 & ~n3584 ;
  assign n3586 = n161 | n2276 ;
  assign n3587 = n2084 | n2945 ;
  assign n3588 = n3586 | n3587 ;
  assign n3589 = n304 | n3588 ;
  assign n3590 = n87 | n2839 ;
  assign n3591 = n3589 | n3590 ;
  assign n3592 = n185 | n573 ;
  assign n3593 = n1041 | n3592 ;
  assign n3594 = n147 | n279 ;
  assign n3595 = n3593 | n3594 ;
  assign n3596 = n2902 | n3595 ;
  assign n3597 = n581 | n3409 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3591 | n3598 ;
  assign n3600 = n3585 & ~n3599 ;
  assign n3601 = ~n3554 & n3600 ;
  assign n3602 = ~n3488 & n3601 ;
  assign n3603 = n3533 | n3602 ;
  assign n3604 = ~n3264 & n3487 ;
  assign n3605 = n3601 | n3604 ;
  assign n3606 = n3533 & n3605 ;
  assign n3607 = n3516 | n3606 ;
  assign n3608 = ~n3516 & n3606 ;
  assign n3609 = ( ~n3603 & n3607 ) | ( ~n3603 & n3608 ) | ( n3607 & n3608 ) ;
  assign n3610 = ( n3537 & n3542 ) | ( n3537 & n3609 ) | ( n3542 & n3609 ) ;
  assign n3611 = x29 & ~n3610 ;
  assign n3612 = ( ~x29 & n3517 ) | ( ~x29 & n3610 ) | ( n3517 & n3610 ) ;
  assign n3613 = ( ~n3518 & n3611 ) | ( ~n3518 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3614 = n412 | n432 ;
  assign n3615 = n1119 | n1401 ;
  assign n3616 = n3614 | n3615 ;
  assign n3617 = n780 | n2490 ;
  assign n3618 = n1544 | n3617 ;
  assign n3619 = n3616 | n3618 ;
  assign n3620 = n287 | n835 ;
  assign n3621 = n1694 | n3620 ;
  assign n3622 = n164 | n464 ;
  assign n3623 = n144 | n207 ;
  assign n3624 = n3622 | n3623 ;
  assign n3625 = n3621 | n3624 ;
  assign n3626 = n2605 | n3625 ;
  assign n3627 = n3619 | n3626 ;
  assign n3628 = n2818 | n3627 ;
  assign n3629 = n2673 | n3628 ;
  assign n3630 = n509 | n1224 ;
  assign n3631 = n127 | n3630 ;
  assign n3632 = n913 | n1374 ;
  assign n3633 = n303 | n518 ;
  assign n3634 = n82 | n712 ;
  assign n3635 = n3633 | n3634 ;
  assign n3636 = n3632 | n3635 ;
  assign n3637 = n3631 | n3636 ;
  assign n3638 = n695 | n1803 ;
  assign n3639 = n337 | n497 ;
  assign n3640 = n264 | n3639 ;
  assign n3641 = n742 | n3640 ;
  assign n3642 = n3638 | n3641 ;
  assign n3643 = n3637 | n3642 ;
  assign n3644 = n1038 & ~n3643 ;
  assign n3645 = n640 | n2935 ;
  assign n3646 = n939 | n1413 ;
  assign n3647 = n3645 | n3646 ;
  assign n3648 = n296 | n916 ;
  assign n3649 = n163 | n341 ;
  assign n3650 = n3648 | n3649 ;
  assign n3651 = n2412 | n2567 ;
  assign n3652 = n3650 | n3651 ;
  assign n3653 = n3647 | n3652 ;
  assign n3654 = n3644 & ~n3653 ;
  assign n3655 = n178 | n989 ;
  assign n3656 = n317 | n3655 ;
  assign n3657 = n359 | n1626 ;
  assign n3658 = n3656 | n3657 ;
  assign n3659 = n1735 | n3658 ;
  assign n3660 = n431 | n581 ;
  assign n3661 = n147 | n3660 ;
  assign n3662 = n2276 | n3661 ;
  assign n3663 = n1107 | n3662 ;
  assign n3664 = n3659 | n3663 ;
  assign n3665 = n90 | n1710 ;
  assign n3666 = n254 | n329 ;
  assign n3667 = n1444 | n3666 ;
  assign n3668 = n3665 | n3667 ;
  assign n3669 = n3664 | n3668 ;
  assign n3670 = n3654 & ~n3669 ;
  assign n3671 = ~n3629 & n3670 ;
  assign n3672 = ( n3266 & n3490 ) | ( n3266 & n3601 ) | ( n3490 & n3601 ) ;
  assign n3673 = ( ~n3266 & n3490 ) | ( ~n3266 & n3601 ) | ( n3490 & n3601 ) ;
  assign n3674 = ( n3266 & ~n3672 ) | ( n3266 & n3673 ) | ( ~n3672 & n3673 ) ;
  assign n3675 = n3270 & ~n3601 ;
  assign n3676 = n3274 & ~n3487 ;
  assign n3677 = n3675 | n3676 ;
  assign n3678 = n390 | n3677 ;
  assign n3679 = ( n3674 & n3677 ) | ( n3674 & n3678 ) | ( n3677 & n3678 ) ;
  assign n3680 = n564 & n3273 ;
  assign n3681 = n3679 | n3680 ;
  assign n3682 = ( ~n3402 & n3671 ) | ( ~n3402 & n3681 ) | ( n3671 & n3681 ) ;
  assign n3683 = ( n3402 & n3671 ) | ( n3402 & ~n3681 ) | ( n3671 & ~n3681 ) ;
  assign n3684 = ( ~n3671 & n3682 ) | ( ~n3671 & n3683 ) | ( n3682 & n3683 ) ;
  assign n3685 = ( n3496 & n3613 ) | ( n3496 & n3684 ) | ( n3613 & n3684 ) ;
  assign n3686 = n55 | n751 ;
  assign n3687 = n1058 | n3686 ;
  assign n3688 = n90 | n1020 ;
  assign n3689 = n3687 | n3688 ;
  assign n3690 = n221 | n323 ;
  assign n3691 = n232 | n3690 ;
  assign n3692 = n3689 | n3691 ;
  assign n3693 = n2271 | n3692 ;
  assign n3694 = n465 | n688 ;
  assign n3695 = n1994 | n3694 ;
  assign n3696 = n962 | n1176 ;
  assign n3697 = n3695 | n3696 ;
  assign n3698 = n3693 | n3697 ;
  assign n3699 = n351 | n750 ;
  assign n3700 = n756 | n3699 ;
  assign n3701 = n208 | n488 ;
  assign n3702 = n434 | n3701 ;
  assign n3703 = n3344 | n3702 ;
  assign n3704 = n3700 | n3703 ;
  assign n3705 = n402 | n1041 ;
  assign n3706 = n134 | n264 ;
  assign n3707 = n3705 | n3706 ;
  assign n3708 = n487 | n1137 ;
  assign n3709 = n329 | n1044 ;
  assign n3710 = n3708 | n3709 ;
  assign n3711 = n3707 | n3710 ;
  assign n3712 = n3704 | n3711 ;
  assign n3713 = n3698 | n3712 ;
  assign n3714 = n133 | n242 ;
  assign n3715 = n225 | n296 ;
  assign n3716 = n990 | n3715 ;
  assign n3717 = n3714 | n3716 ;
  assign n3718 = n904 | n1993 ;
  assign n3719 = n3717 | n3718 ;
  assign n3720 = n346 | n1074 ;
  assign n3721 = n3064 | n3720 ;
  assign n3722 = n3719 | n3721 ;
  assign n3723 = n3713 | n3722 ;
  assign n3724 = n97 | n338 ;
  assign n3725 = n2828 | n3724 ;
  assign n3726 = n190 | n1630 ;
  assign n3727 = n270 | n3726 ;
  assign n3728 = n3725 | n3727 ;
  assign n3729 = n191 | n284 ;
  assign n3730 = n497 | n500 ;
  assign n3731 = n3729 | n3730 ;
  assign n3732 = n915 | n3731 ;
  assign n3733 = n317 | n362 ;
  assign n3734 = n2019 | n3733 ;
  assign n3735 = n3732 | n3734 ;
  assign n3736 = n3728 | n3735 ;
  assign n3737 = n113 | n485 ;
  assign n3738 = n368 | n3737 ;
  assign n3739 = n1998 | n2420 ;
  assign n3740 = n3738 | n3739 ;
  assign n3741 = n3736 | n3740 ;
  assign n3742 = n129 | n238 ;
  assign n3743 = n328 | n1126 ;
  assign n3744 = n3742 | n3743 ;
  assign n3745 = n1006 | n1069 ;
  assign n3746 = n285 | n3745 ;
  assign n3747 = n3744 | n3746 ;
  assign n3748 = n1893 | n3747 ;
  assign n3749 = n3741 | n3748 ;
  assign n3750 = n3723 | n3749 ;
  assign n3751 = n601 | n2357 ;
  assign n3752 = n116 | n3220 ;
  assign n3753 = n3751 | n3752 ;
  assign n3754 = n256 | n546 ;
  assign n3755 = n370 | n915 ;
  assign n3756 = n3754 | n3755 ;
  assign n3757 = n834 | n3756 ;
  assign n3758 = n3753 | n3757 ;
  assign n3759 = n305 | n1094 ;
  assign n3760 = n265 | n3759 ;
  assign n3761 = x25 & n217 ;
  assign n3762 = n3760 | n3761 ;
  assign n3763 = n210 | n487 ;
  assign n3764 = n578 | n3763 ;
  assign n3765 = n3762 | n3764 ;
  assign n3766 = n518 | n750 ;
  assign n3767 = n332 | n3766 ;
  assign n3768 = n3765 | n3767 ;
  assign n3769 = n3758 | n3768 ;
  assign n3770 = n1419 | n2690 ;
  assign n3771 = n534 | n688 ;
  assign n3772 = n2144 | n3771 ;
  assign n3773 = n1542 | n3772 ;
  assign n3774 = n3770 | n3773 ;
  assign n3775 = n2098 | n3774 ;
  assign n3776 = n164 | n374 ;
  assign n3777 = n268 | n318 ;
  assign n3778 = n3776 | n3777 ;
  assign n3779 = n1110 | n3560 ;
  assign n3780 = n3778 | n3779 ;
  assign n3781 = n3775 | n3780 ;
  assign n3782 = n1172 | n2107 ;
  assign n3783 = n222 | n1060 ;
  assign n3784 = n3782 | n3783 ;
  assign n3785 = n1105 | n3784 ;
  assign n3786 = n270 | n524 ;
  assign n3787 = n3362 | n3786 ;
  assign n3788 = n3785 | n3787 ;
  assign n3789 = n3781 | n3788 ;
  assign n3790 = n3769 | n3789 ;
  assign n3791 = n151 | n346 ;
  assign n3792 = n1505 | n3690 ;
  assign n3793 = n3791 | n3792 ;
  assign n3794 = n1718 | n3793 ;
  assign n3795 = n556 | n635 ;
  assign n3796 = n232 | n3795 ;
  assign n3797 = n677 | n3796 ;
  assign n3798 = n3794 | n3797 ;
  assign n3799 = n99 | n526 ;
  assign n3800 = n655 | n3799 ;
  assign n3801 = n422 | n1020 ;
  assign n3802 = n3800 | n3801 ;
  assign n3803 = n173 | n1014 ;
  assign n3804 = n2707 | n3803 ;
  assign n3805 = n3802 | n3804 ;
  assign n3806 = n457 | n1107 ;
  assign n3807 = n2658 | n3806 ;
  assign n3808 = n3805 | n3807 ;
  assign n3809 = n3798 | n3808 ;
  assign n3810 = n1984 | n2051 ;
  assign n3811 = n285 | n335 ;
  assign n3812 = n125 | n3811 ;
  assign n3813 = n3810 | n3812 ;
  assign n3814 = n357 | n614 ;
  assign n3815 = n446 | n3814 ;
  assign n3816 = n3813 | n3815 ;
  assign n3817 = n449 | n704 ;
  assign n3818 = n363 | n647 ;
  assign n3819 = n3817 | n3818 ;
  assign n3820 = n692 | n1123 ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = n2333 | n3821 ;
  assign n3823 = n3816 | n3822 ;
  assign n3824 = n3809 | n3823 ;
  assign n3825 = n3790 | n3824 ;
  assign n3826 = ( ~x23 & n3750 ) | ( ~x23 & n3825 ) | ( n3750 & n3825 ) ;
  assign n3827 = n3151 & n3263 ;
  assign n3828 = n3152 & ~n3262 ;
  assign n3829 = ( n721 & ~n3827 ) | ( n721 & n3828 ) | ( ~n3827 & n3828 ) ;
  assign n3830 = n995 & n3273 ;
  assign n3831 = ~n721 & n3270 ;
  assign n3832 = n3830 | n3831 ;
  assign n3833 = n859 & n3274 ;
  assign n3834 = n3832 | n3833 ;
  assign n3835 = n390 | n3834 ;
  assign n3836 = ( ~n3829 & n3834 ) | ( ~n3829 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3837 = ( ~n388 & n3826 ) | ( ~n388 & n3836 ) | ( n3826 & n3836 ) ;
  assign n3838 = ~n1118 & n3259 ;
  assign n3839 = ( n1118 & n3148 ) | ( n1118 & n3259 ) | ( n3148 & n3259 ) ;
  assign n3840 = n1118 | n3148 ;
  assign n3841 = ( n3838 & ~n3839 ) | ( n3838 & n3840 ) | ( ~n3839 & n3840 ) ;
  assign n3842 = ~n1118 & n3270 ;
  assign n3843 = ~n1207 & n3274 ;
  assign n3844 = n3842 | n3843 ;
  assign n3845 = n1316 & n3273 ;
  assign n3846 = n3844 | n3845 ;
  assign n3847 = n390 | n3846 ;
  assign n3848 = ( n3841 & n3846 ) | ( n3841 & n3847 ) | ( n3846 & n3847 ) ;
  assign n3849 = n238 | n593 ;
  assign n3850 = n3459 | n3849 ;
  assign n3851 = n3183 | n3850 ;
  assign n3852 = n1331 | n1392 ;
  assign n3853 = n202 | n1166 ;
  assign n3854 = n3852 | n3853 ;
  assign n3855 = n3851 | n3854 ;
  assign n3856 = n2077 | n3855 ;
  assign n3857 = n1537 | n2431 ;
  assign n3858 = n480 | n647 ;
  assign n3859 = n315 | n3858 ;
  assign n3860 = n975 | n3859 ;
  assign n3861 = n3857 | n3860 ;
  assign n3862 = n1715 | n3861 ;
  assign n3863 = n3856 | n3862 ;
  assign n3864 = n528 | n751 ;
  assign n3865 = n285 | n3864 ;
  assign n3866 = n165 | n600 ;
  assign n3867 = n2670 | n3866 ;
  assign n3868 = n3865 | n3867 ;
  assign n3869 = n3025 | n3868 ;
  assign n3870 = n607 | n2307 ;
  assign n3871 = n3869 | n3870 ;
  assign n3872 = n1909 | n2010 ;
  assign n3873 = n3871 | n3872 ;
  assign n3874 = n129 | n2762 ;
  assign n3875 = n750 | n3874 ;
  assign n3876 = n160 | n705 ;
  assign n3877 = n509 | n3876 ;
  assign n3878 = n1689 | n1998 ;
  assign n3879 = n3877 | n3878 ;
  assign n3880 = n3875 | n3879 ;
  assign n3881 = n3873 | n3880 ;
  assign n3882 = n3863 | n3881 ;
  assign n3883 = n314 | n611 ;
  assign n3884 = n2754 | n3883 ;
  assign n3885 = n147 | n163 ;
  assign n3886 = n969 | n3885 ;
  assign n3887 = n3884 | n3886 ;
  assign n3888 = n190 | n2506 ;
  assign n3889 = n3468 | n3888 ;
  assign n3890 = n3887 | n3889 ;
  assign n3891 = n131 | n362 ;
  assign n3892 = n742 | n3891 ;
  assign n3893 = n1325 | n1429 ;
  assign n3894 = n3892 | n3893 ;
  assign n3895 = n1226 | n3021 ;
  assign n3896 = n3894 | n3895 ;
  assign n3897 = n2210 | n3052 ;
  assign n3898 = n431 | n442 ;
  assign n3899 = n3666 | n3898 ;
  assign n3900 = n3897 | n3899 ;
  assign n3901 = n3896 | n3900 ;
  assign n3902 = n2375 | n3901 ;
  assign n3903 = n3890 | n3902 ;
  assign n3904 = n3882 | n3903 ;
  assign n3905 = n294 | n380 ;
  assign n3906 = n2758 | n3905 ;
  assign n3907 = n486 | n935 ;
  assign n3908 = n3906 | n3907 ;
  assign n3909 = n708 | n1166 ;
  assign n3910 = n3908 | n3909 ;
  assign n3911 = n1745 | n1763 ;
  assign n3912 = n1351 | n1399 ;
  assign n3913 = n3911 | n3912 ;
  assign n3914 = n3910 | n3913 ;
  assign n3915 = n550 | n915 ;
  assign n3916 = n3791 | n3915 ;
  assign n3917 = n269 | n279 ;
  assign n3918 = n1590 | n3917 ;
  assign n3919 = n51 & n95 ;
  assign n3920 = n374 | n3919 ;
  assign n3921 = n3918 | n3920 ;
  assign n3922 = n3916 | n3921 ;
  assign n3923 = n242 | n341 ;
  assign n3924 = n134 | n3923 ;
  assign n3925 = n2982 | n3924 ;
  assign n3926 = n3922 | n3925 ;
  assign n3927 = n3914 | n3926 ;
  assign n3928 = n794 | n1291 ;
  assign n3929 = n968 | n3928 ;
  assign n3930 = n110 | n184 ;
  assign n3931 = n987 | n3930 ;
  assign n3932 = n2752 | n3931 ;
  assign n3933 = n3929 | n3932 ;
  assign n3934 = n407 | n781 ;
  assign n3935 = n87 | n1518 ;
  assign n3936 = n3934 | n3935 ;
  assign n3937 = n1113 | n1843 ;
  assign n3938 = n3936 | n3937 ;
  assign n3939 = n3933 | n3938 ;
  assign n3940 = n2055 | n3939 ;
  assign n3941 = n1294 | n3425 ;
  assign n3942 = n308 | n722 ;
  assign n3943 = n3941 | n3942 ;
  assign n3944 = n883 | n1241 ;
  assign n3945 = n74 | n164 ;
  assign n3946 = n315 | n688 ;
  assign n3947 = n3945 | n3946 ;
  assign n3948 = n3944 | n3947 ;
  assign n3949 = n3943 | n3948 ;
  assign n3950 = n3940 | n3949 ;
  assign n3951 = n108 | n586 ;
  assign n3952 = n82 | n402 ;
  assign n3953 = n3951 | n3952 ;
  assign n3954 = n378 | n689 ;
  assign n3955 = n350 | n3954 ;
  assign n3956 = n3953 | n3955 ;
  assign n3957 = n723 | n835 ;
  assign n3958 = n176 | n301 ;
  assign n3959 = n3957 | n3958 ;
  assign n3960 = n971 | n3959 ;
  assign n3961 = n3956 | n3960 ;
  assign n3962 = n666 | n3961 ;
  assign n3963 = n842 | n2935 ;
  assign n3964 = n990 | n3963 ;
  assign n3965 = n364 | n2773 ;
  assign n3966 = n600 | n860 ;
  assign n3967 = n3454 | n3966 ;
  assign n3968 = n3965 | n3967 ;
  assign n3969 = n3964 | n3968 ;
  assign n3970 = n546 | n921 ;
  assign n3971 = n141 | n275 ;
  assign n3972 = n3666 | n3971 ;
  assign n3973 = n3970 | n3972 ;
  assign n3974 = n244 | n405 ;
  assign n3975 = n2897 | n3974 ;
  assign n3976 = n123 | n3975 ;
  assign n3977 = n3973 | n3976 ;
  assign n3978 = n3969 | n3977 ;
  assign n3979 = n3962 | n3978 ;
  assign n3980 = n3950 | n3979 ;
  assign n3981 = n3927 | n3980 ;
  assign n3982 = ( ~x20 & n3904 ) | ( ~x20 & n3981 ) | ( n3904 & n3981 ) ;
  assign n3983 = n2983 | n3883 ;
  assign n3984 = n929 | n3218 ;
  assign n3985 = n3983 | n3984 ;
  assign n3986 = n2842 & ~n3622 ;
  assign n3987 = n419 | n617 ;
  assign n3988 = n3986 & ~n3987 ;
  assign n3989 = ~n3985 & n3988 ;
  assign n3990 = ~n1215 & n3989 ;
  assign n3991 = ~n2819 & n3990 ;
  assign n3992 = n242 | n723 ;
  assign n3993 = n2698 | n3992 ;
  assign n3994 = n104 | n245 ;
  assign n3995 = n335 | n432 ;
  assign n3996 = n3994 | n3995 ;
  assign n3997 = n3993 | n3996 ;
  assign n3998 = n2308 | n3997 ;
  assign n3999 = n237 | n3453 ;
  assign n4000 = n403 | n3999 ;
  assign n4001 = n518 | n922 ;
  assign n4002 = n226 | n4001 ;
  assign n4003 = n1184 | n4002 ;
  assign n4004 = n4000 | n4003 ;
  assign n4005 = n3998 | n4004 ;
  assign n4006 = n129 | n679 ;
  assign n4007 = n221 | n428 ;
  assign n4008 = n178 | n494 ;
  assign n4009 = n1044 | n4008 ;
  assign n4010 = n4007 | n4009 ;
  assign n4011 = n4006 | n4010 ;
  assign n4012 = n3214 | n4011 ;
  assign n4013 = n4005 | n4012 ;
  assign n4014 = n1908 | n3898 ;
  assign n4015 = n338 | n500 ;
  assign n4016 = n80 | n4015 ;
  assign n4017 = n1750 | n4016 ;
  assign n4018 = n4014 | n4017 ;
  assign n4019 = n1399 | n1955 ;
  assign n4020 = n4018 | n4019 ;
  assign n4021 = n1583 | n4020 ;
  assign n4022 = n4013 | n4021 ;
  assign n4023 = n3991 & ~n4022 ;
  assign n4024 = ( n3848 & ~n3982 ) | ( n3848 & n4023 ) | ( ~n3982 & n4023 ) ;
  assign n4025 = ( n3750 & ~n3848 ) | ( n3750 & n4024 ) | ( ~n3848 & n4024 ) ;
  assign n4026 = n859 & n3270 ;
  assign n4027 = ~n1118 & n3273 ;
  assign n4028 = n4026 | n4027 ;
  assign n4029 = n995 & n3274 ;
  assign n4030 = n4028 | n4029 ;
  assign n4031 = n390 | n4030 ;
  assign n4032 = n3151 | n3261 ;
  assign n4033 = ~n3150 & n3262 ;
  assign n4034 = ( ~n859 & n4032 ) | ( ~n859 & n4033 ) | ( n4032 & n4033 ) ;
  assign n4035 = ( n4030 & n4031 ) | ( n4030 & ~n4034 ) | ( n4031 & ~n4034 ) ;
  assign n4036 = ( x23 & n3750 ) | ( x23 & n3825 ) | ( n3750 & n3825 ) ;
  assign n4037 = ( x23 & n3826 ) | ( x23 & ~n4036 ) | ( n3826 & ~n4036 ) ;
  assign n4038 = ( n4025 & ~n4035 ) | ( n4025 & n4037 ) | ( ~n4035 & n4037 ) ;
  assign n4039 = n3500 & ~n3540 ;
  assign n4040 = ~n3601 & n4039 ;
  assign n4041 = n564 & n3536 ;
  assign n4042 = n4040 | n4041 ;
  assign n4043 = ~n3487 & n3501 ;
  assign n4044 = n4042 | n4043 ;
  assign n4045 = n3541 | n4044 ;
  assign n4046 = ( n3674 & n4044 ) | ( n3674 & n4045 ) | ( n4044 & n4045 ) ;
  assign n4047 = x29 & ~n4046 ;
  assign n4048 = ~x29 & n4046 ;
  assign n4049 = n4047 | n4048 ;
  assign n4050 = ( n388 & ~n3826 ) | ( n388 & n3836 ) | ( ~n3826 & n3836 ) ;
  assign n4051 = ( ~n3836 & n3837 ) | ( ~n3836 & n4050 ) | ( n3837 & n4050 ) ;
  assign n4052 = ( n4038 & ~n4049 ) | ( n4038 & n4051 ) | ( ~n4049 & n4051 ) ;
  assign n4053 = ( n388 & n3279 ) | ( n388 & n3342 ) | ( n3279 & n3342 ) ;
  assign n4054 = ( n388 & n3343 ) | ( n388 & ~n4053 ) | ( n3343 & ~n4053 ) ;
  assign n4055 = ( ~n3837 & n4052 ) | ( ~n3837 & n4054 ) | ( n4052 & n4054 ) ;
  assign n4056 = ( n3516 & ~n3603 ) | ( n3516 & n3606 ) | ( ~n3603 & n3606 ) ;
  assign n4057 = ~n3516 & n3603 ;
  assign n4058 = ( ~n3608 & n4056 ) | ( ~n3608 & n4057 ) | ( n4056 & n4057 ) ;
  assign n4059 = n3501 & ~n3533 ;
  assign n4060 = n3516 | n4039 ;
  assign n4061 = n3516 & ~n3536 ;
  assign n4062 = ( n4059 & n4060 ) | ( n4059 & ~n4061 ) | ( n4060 & ~n4061 ) ;
  assign n4063 = n3541 | n4062 ;
  assign n4064 = ( ~n4058 & n4062 ) | ( ~n4058 & n4063 ) | ( n4062 & n4063 ) ;
  assign n4065 = x29 & ~n4064 ;
  assign n4066 = ~x29 & n4064 ;
  assign n4067 = n4065 | n4066 ;
  assign n4068 = ( n3343 & n3403 ) | ( n3343 & ~n3495 ) | ( n3403 & ~n3495 ) ;
  assign n4069 = ( ~n3343 & n3496 ) | ( ~n3343 & n4068 ) | ( n3496 & n4068 ) ;
  assign n4070 = ( n4055 & ~n4067 ) | ( n4055 & n4069 ) | ( ~n4067 & n4069 ) ;
  assign n4071 = n859 & n3501 ;
  assign n4072 = ~n721 & n4039 ;
  assign n4073 = n4071 | n4072 ;
  assign n4074 = n995 & n3536 ;
  assign n4075 = n4073 | n4074 ;
  assign n4076 = n3541 | n4075 ;
  assign n4077 = ( ~n3829 & n4075 ) | ( ~n3829 & n4076 ) | ( n4075 & n4076 ) ;
  assign n4078 = x29 & ~n4077 ;
  assign n4079 = ~x29 & n4077 ;
  assign n4080 = n4078 | n4079 ;
  assign n4081 = n1316 & ~n3257 ;
  assign n4082 = ( n1316 & ~n3146 ) | ( n1316 & n3257 ) | ( ~n3146 & n3257 ) ;
  assign n4083 = n1316 & ~n3146 ;
  assign n4084 = ( n4081 & n4082 ) | ( n4081 & ~n4083 ) | ( n4082 & ~n4083 ) ;
  assign n4085 = n1316 & n3270 ;
  assign n4086 = ~n1529 & n3273 ;
  assign n4087 = n4085 | n4086 ;
  assign n4088 = n1398 & n3274 ;
  assign n4089 = n4087 | n4088 ;
  assign n4090 = n390 | n4089 ;
  assign n4091 = ( n4084 & n4089 ) | ( n4084 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4092 = n500 | n723 ;
  assign n4093 = n583 | n4092 ;
  assign n4094 = n615 | n954 ;
  assign n4095 = n4093 | n4094 ;
  assign n4096 = n1439 | n1601 ;
  assign n4097 = n1169 | n4096 ;
  assign n4098 = n1077 | n4097 ;
  assign n4099 = n4095 | n4098 ;
  assign n4100 = n1020 | n2748 ;
  assign n4101 = n306 | n442 ;
  assign n4102 = n242 | n345 ;
  assign n4103 = n4101 | n4102 ;
  assign n4104 = n4100 | n4103 ;
  assign n4105 = n2995 | n4104 ;
  assign n4106 = n4099 | n4105 ;
  assign n4107 = n1081 | n1799 ;
  assign n4108 = n1287 | n4107 ;
  assign n4109 = n74 | n1762 ;
  assign n4110 = n1737 | n4109 ;
  assign n4111 = n4108 | n4110 ;
  assign n4112 = n214 | n3026 ;
  assign n4113 = n2030 | n4112 ;
  assign n4114 = n4111 | n4113 ;
  assign n4115 = n4106 | n4114 ;
  assign n4116 = n1306 | n4115 ;
  assign n4117 = n147 | n413 ;
  assign n4118 = n677 | n4117 ;
  assign n4119 = n1524 | n4118 ;
  assign n4120 = n547 | n4119 ;
  assign n4121 = n919 | n1551 ;
  assign n4122 = n280 | n1518 ;
  assign n4123 = n456 | n1253 ;
  assign n4124 = n4122 | n4123 ;
  assign n4125 = n124 | n322 ;
  assign n4126 = n851 | n4125 ;
  assign n4127 = n3656 | n4126 ;
  assign n4128 = n4124 | n4127 ;
  assign n4129 = n4121 | n4128 ;
  assign n4130 = n4120 | n4129 ;
  assign n4131 = n104 | n314 ;
  assign n4132 = n215 | n850 ;
  assign n4133 = n308 | n4132 ;
  assign n4134 = n4131 | n4133 ;
  assign n4135 = n253 | n465 ;
  assign n4136 = n1409 | n4135 ;
  assign n4137 = n4134 | n4136 ;
  assign n4138 = n4130 | n4137 ;
  assign n4139 = n153 | n331 ;
  assign n4140 = n1399 | n4139 ;
  assign n4141 = n474 | n4140 ;
  assign n4142 = n201 | n1695 ;
  assign n4143 = n318 | n3686 ;
  assign n4144 = n4142 | n4143 ;
  assign n4145 = n4141 | n4144 ;
  assign n4146 = n2689 | n4145 ;
  assign n4147 = n268 | n440 ;
  assign n4148 = n2458 & ~n4147 ;
  assign n4149 = ~n986 & n4148 ;
  assign n4150 = ~n4146 & n4149 ;
  assign n4151 = ~n4138 & n4150 ;
  assign n4152 = ~n4116 & n4151 ;
  assign n4153 = ( n3904 & ~n4091 ) | ( n3904 & n4152 ) | ( ~n4091 & n4152 ) ;
  assign n4154 = ~n1207 & n3258 ;
  assign n4155 = n1207 & n3258 ;
  assign n4156 = ( n1207 & ~n3147 ) | ( n1207 & n4155 ) | ( ~n3147 & n4155 ) ;
  assign n4157 = ( n3148 & ~n4154 ) | ( n3148 & n4156 ) | ( ~n4154 & n4156 ) ;
  assign n4158 = n1316 & n3274 ;
  assign n4159 = ~n1207 & n3270 ;
  assign n4160 = n1398 & n3273 ;
  assign n4161 = n4159 | n4160 ;
  assign n4162 = n4158 | n4161 ;
  assign n4163 = n390 | n4162 ;
  assign n4164 = ( ~n4157 & n4162 ) | ( ~n4157 & n4163 ) | ( n4162 & n4163 ) ;
  assign n4165 = ( x20 & n3904 ) | ( x20 & n3981 ) | ( n3904 & n3981 ) ;
  assign n4166 = ( x20 & n3982 ) | ( x20 & ~n4165 ) | ( n3982 & ~n4165 ) ;
  assign n4167 = ( n4153 & ~n4164 ) | ( n4153 & n4166 ) | ( ~n4164 & n4166 ) ;
  assign n4168 = ( n3848 & n3982 ) | ( n3848 & ~n4023 ) | ( n3982 & ~n4023 ) ;
  assign n4169 = ( ~n3848 & n4024 ) | ( ~n3848 & n4168 ) | ( n4024 & n4168 ) ;
  assign n4170 = ( n4080 & ~n4167 ) | ( n4080 & n4169 ) | ( ~n4167 & n4169 ) ;
  assign n4171 = n995 & ~n3260 ;
  assign n4172 = ( n995 & ~n3149 ) | ( n995 & n3260 ) | ( ~n3149 & n3260 ) ;
  assign n4173 = ( ~n3150 & n4171 ) | ( ~n3150 & n4172 ) | ( n4171 & n4172 ) ;
  assign n4174 = n995 & n3270 ;
  assign n4175 = ~n1207 & n3273 ;
  assign n4176 = n4174 | n4175 ;
  assign n4177 = ~n1118 & n3274 ;
  assign n4178 = n4176 | n4177 ;
  assign n4179 = n390 | n4178 ;
  assign n4180 = ( n4173 & n4178 ) | ( n4173 & n4179 ) | ( n4178 & n4179 ) ;
  assign n4181 = ( n3750 & n3848 ) | ( n3750 & n4024 ) | ( n3848 & n4024 ) ;
  assign n4182 = ( n3848 & n4025 ) | ( n3848 & ~n4181 ) | ( n4025 & ~n4181 ) ;
  assign n4183 = ( n4170 & n4180 ) | ( n4170 & n4182 ) | ( n4180 & n4182 ) ;
  assign n4184 = ( n4025 & n4035 ) | ( n4025 & ~n4037 ) | ( n4035 & ~n4037 ) ;
  assign n4185 = ( ~n4025 & n4038 ) | ( ~n4025 & n4184 ) | ( n4038 & n4184 ) ;
  assign n4186 = n564 & n3501 ;
  assign n4187 = ~n721 & n3536 ;
  assign n4188 = n4186 | n4187 ;
  assign n4189 = ~n3487 & n4039 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = n3541 | n4190 ;
  assign n4192 = ( ~n3492 & n4190 ) | ( ~n3492 & n4191 ) | ( n4190 & n4191 ) ;
  assign n4193 = x29 & ~n4192 ;
  assign n4194 = ~x29 & n4192 ;
  assign n4195 = n4193 | n4194 ;
  assign n4196 = ( n4183 & n4185 ) | ( n4183 & n4195 ) | ( n4185 & n4195 ) ;
  assign n4197 = n2083 & ~n3533 ;
  assign n4198 = x26 & n4197 ;
  assign n4199 = x25 | n59 ;
  assign n4200 = ( ~n72 & n3091 ) | ( ~n72 & n4199 ) | ( n3091 & n4199 ) ;
  assign n4201 = ~n3516 & n4200 ;
  assign n4202 = n53 | n68 ;
  assign n4203 = n506 & n4202 ;
  assign n4204 = n4201 | n4203 ;
  assign n4205 = ( n3609 & n4201 ) | ( n3609 & n4204 ) | ( n4201 & n4204 ) ;
  assign n4206 = x26 & ~n4205 ;
  assign n4207 = ( ~x26 & n4197 ) | ( ~x26 & n4205 ) | ( n4197 & n4205 ) ;
  assign n4208 = ( ~n4198 & n4206 ) | ( ~n4198 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = ( n4038 & n4049 ) | ( n4038 & ~n4051 ) | ( n4049 & ~n4051 ) ;
  assign n4210 = ( ~n4038 & n4052 ) | ( ~n4038 & n4209 ) | ( n4052 & n4209 ) ;
  assign n4211 = ( n4196 & n4208 ) | ( n4196 & n4210 ) | ( n4208 & n4210 ) ;
  assign n4212 = ( ~n4170 & n4180 ) | ( ~n4170 & n4182 ) | ( n4180 & n4182 ) ;
  assign n4213 = ( n4170 & ~n4183 ) | ( n4170 & n4212 ) | ( ~n4183 & n4212 ) ;
  assign n4214 = ~n3601 & n4200 ;
  assign n4215 = ~n506 & n4202 ;
  assign n4216 = ~n3533 & n4215 ;
  assign n4217 = n4214 | n4216 ;
  assign n4218 = n2083 & ~n3487 ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = n4203 | n4219 ;
  assign n4221 = ~n3602 & n3606 ;
  assign n4222 = ~n3603 & n3605 ;
  assign n4223 = ( n3533 & ~n4221 ) | ( n3533 & n4222 ) | ( ~n4221 & n4222 ) ;
  assign n4224 = ( n4219 & n4220 ) | ( n4219 & ~n4223 ) | ( n4220 & ~n4223 ) ;
  assign n4225 = x26 & ~n4224 ;
  assign n4226 = ~x26 & n4224 ;
  assign n4227 = n4225 | n4226 ;
  assign n4228 = n859 & n3536 ;
  assign n4229 = ~n721 & n3501 ;
  assign n4230 = n4228 | n4229 ;
  assign n4231 = n564 & n4039 ;
  assign n4232 = n4230 | n4231 ;
  assign n4233 = n3541 | n4232 ;
  assign n4234 = ( ~n3268 & n4232 ) | ( ~n3268 & n4233 ) | ( n4232 & n4233 ) ;
  assign n4235 = x29 & ~n4234 ;
  assign n4236 = ~x29 & n4234 ;
  assign n4237 = n4235 | n4236 ;
  assign n4238 = ( n4213 & n4227 ) | ( n4213 & n4237 ) | ( n4227 & n4237 ) ;
  assign n4239 = ( ~n4183 & n4185 ) | ( ~n4183 & n4195 ) | ( n4185 & n4195 ) ;
  assign n4240 = ( n4183 & ~n4196 ) | ( n4183 & n4239 ) | ( ~n4196 & n4239 ) ;
  assign n4241 = ~n3516 & n4215 ;
  assign n4242 = n2083 | n4241 ;
  assign n4243 = ( ~n3601 & n4241 ) | ( ~n3601 & n4242 ) | ( n4241 & n4242 ) ;
  assign n4244 = ~n3533 & n4200 ;
  assign n4245 = n4243 | n4244 ;
  assign n4246 = n4203 | n4245 ;
  assign n4247 = ( ~n4058 & n4245 ) | ( ~n4058 & n4246 ) | ( n4245 & n4246 ) ;
  assign n4248 = x26 & ~n4247 ;
  assign n4249 = ~x26 & n4247 ;
  assign n4250 = n4248 | n4249 ;
  assign n4251 = ( n4238 & n4240 ) | ( n4238 & n4250 ) | ( n4240 & n4250 ) ;
  assign n4252 = n1593 | n1793 ;
  assign n4253 = n440 | n989 ;
  assign n4254 = n1095 | n4253 ;
  assign n4255 = n4252 | n4254 ;
  assign n4256 = n70 | n976 ;
  assign n4257 = n1124 | n4256 ;
  assign n4258 = n4255 | n4257 ;
  assign n4259 = n3929 | n4258 ;
  assign n4260 = n3461 | n4259 ;
  assign n4261 = n1057 | n2655 ;
  assign n4262 = n396 | n1547 ;
  assign n4263 = n1277 | n2123 ;
  assign n4264 = n4262 | n4263 ;
  assign n4265 = n4261 | n4264 ;
  assign n4266 = n4260 | n4265 ;
  assign n4267 = n653 & ~n2942 ;
  assign n4268 = ~n4266 & n4267 ;
  assign n4269 = n1663 | n2211 ;
  assign n4270 = n104 | n455 ;
  assign n4271 = n308 | n440 ;
  assign n4272 = n4270 | n4271 ;
  assign n4273 = n4269 | n4272 ;
  assign n4274 = n606 | n4273 ;
  assign n4275 = n328 | n524 ;
  assign n4276 = n643 | n4275 ;
  assign n4277 = n1874 | n4276 ;
  assign n4278 = n4274 | n4277 ;
  assign n4279 = n150 | n989 ;
  assign n4280 = ( n217 & n1100 ) | ( n217 & ~n3761 ) | ( n1100 & ~n3761 ) ;
  assign n4281 = n4279 | n4280 ;
  assign n4282 = n1781 | n4281 ;
  assign n4283 = n4278 | n4282 ;
  assign n4284 = n160 | n1048 ;
  assign n4285 = n1745 | n4284 ;
  assign n4286 = n197 | n1074 ;
  assign n4287 = n4285 | n4286 ;
  assign n4288 = n640 | n850 ;
  assign n4289 = n1420 | n4288 ;
  assign n4290 = n683 | n2123 ;
  assign n4291 = n4289 | n4290 ;
  assign n4292 = n4287 | n4291 ;
  assign n4293 = n4283 | n4292 ;
  assign n4294 = n285 | n723 ;
  assign n4295 = n151 | n269 ;
  assign n4296 = n4294 | n4295 ;
  assign n4297 = n2172 | n4296 ;
  assign n4298 = n580 | n4297 ;
  assign n4299 = n379 | n1332 ;
  assign n4300 = n1199 | n4299 ;
  assign n4301 = n80 | n174 ;
  assign n4302 = n206 | n4301 ;
  assign n4303 = n4300 | n4302 ;
  assign n4304 = n1439 | n4303 ;
  assign n4305 = n4298 | n4304 ;
  assign n4306 = n173 | n321 ;
  assign n4307 = n3080 | n4306 ;
  assign n4308 = n3657 | n4307 ;
  assign n4309 = n1012 | n2030 ;
  assign n4310 = n1134 | n4309 ;
  assign n4311 = n4308 | n4310 ;
  assign n4312 = n4305 | n4311 ;
  assign n4313 = n4293 | n4312 ;
  assign n4314 = n911 | n4313 ;
  assign n4315 = ( x17 & n4268 ) | ( x17 & ~n4314 ) | ( n4268 & ~n4314 ) ;
  assign n4316 = ~n1529 & n3274 ;
  assign n4317 = n1600 & n3273 ;
  assign n4318 = n1398 & n3270 ;
  assign n4319 = n4317 | n4318 ;
  assign n4320 = n4316 | n4319 ;
  assign n4321 = n390 | n4320 ;
  assign n4322 = n3145 | n3257 ;
  assign n4323 = n3146 & ~n3256 ;
  assign n4324 = ( ~n1398 & n4322 ) | ( ~n1398 & n4323 ) | ( n4322 & n4323 ) ;
  assign n4325 = ( n4320 & n4321 ) | ( n4320 & ~n4324 ) | ( n4321 & ~n4324 ) ;
  assign n4326 = ( n3904 & n4315 ) | ( n3904 & ~n4325 ) | ( n4315 & ~n4325 ) ;
  assign n4327 = n3141 | n3252 ;
  assign n4328 = ~n1792 & n4327 ;
  assign n4329 = ( n1687 & n3141 ) | ( n1687 & n4328 ) | ( n3141 & n4328 ) ;
  assign n4330 = ( ~n1687 & n3141 ) | ( ~n1687 & n4328 ) | ( n3141 & n4328 ) ;
  assign n4331 = ( n1687 & ~n4329 ) | ( n1687 & n4330 ) | ( ~n4329 & n4330 ) ;
  assign n4332 = ~n1841 & n3273 ;
  assign n4333 = n1792 & n3274 ;
  assign n4334 = n4332 | n4333 ;
  assign n4335 = n1687 & n3270 ;
  assign n4336 = n4334 | n4335 ;
  assign n4337 = n390 | n4336 ;
  assign n4338 = ( n4331 & n4336 ) | ( n4331 & n4337 ) | ( n4336 & n4337 ) ;
  assign n4339 = n578 | n3080 ;
  assign n4340 = n3714 | n4339 ;
  assign n4341 = n232 | n446 ;
  assign n4342 = n372 | n1044 ;
  assign n4343 = n4341 | n4342 ;
  assign n4344 = n4340 | n4343 ;
  assign n4345 = n150 | n723 ;
  assign n4346 = n237 | n4345 ;
  assign n4347 = n3446 | n4346 ;
  assign n4348 = n303 | n331 ;
  assign n4349 = n683 | n4348 ;
  assign n4350 = n4347 | n4349 ;
  assign n4351 = n4344 | n4350 ;
  assign n4352 = n527 | n587 ;
  assign n4353 = n293 | n533 ;
  assign n4354 = n1682 | n4353 ;
  assign n4355 = n4352 | n4354 ;
  assign n4356 = n2805 | n4355 ;
  assign n4357 = n3875 | n4356 ;
  assign n4358 = n4351 | n4357 ;
  assign n4359 = n306 | n611 ;
  assign n4360 = n206 | n893 ;
  assign n4361 = n4359 | n4360 ;
  assign n4362 = n440 | n1041 ;
  assign n4363 = n925 | n4362 ;
  assign n4364 = n2164 | n4363 ;
  assign n4365 = n4361 | n4364 ;
  assign n4366 = n346 | n468 ;
  assign n4367 = n279 | n835 ;
  assign n4368 = n4366 | n4367 ;
  assign n4369 = n3475 | n4368 ;
  assign n4370 = n4365 | n4369 ;
  assign n4371 = n4358 | n4370 ;
  assign n4372 = n313 | n497 ;
  assign n4373 = n214 | n435 ;
  assign n4374 = n4372 | n4373 ;
  assign n4375 = n556 | n734 ;
  assign n4376 = n4270 | n4375 ;
  assign n4377 = n4374 | n4376 ;
  assign n4378 = n1056 | n1631 ;
  assign n4379 = n4377 | n4378 ;
  assign n4380 = n2981 | n4379 ;
  assign n4381 = n192 | n1176 ;
  assign n4382 = n402 | n4381 ;
  assign n4383 = n3617 | n4382 ;
  assign n4384 = n772 | n987 ;
  assign n4385 = n4383 | n4384 ;
  assign n4386 = n940 | n4385 ;
  assign n4387 = n4380 | n4386 ;
  assign n4388 = n4371 | n4387 ;
  assign n4389 = n1064 | n1489 ;
  assign n4390 = n1649 | n4389 ;
  assign n4391 = n165 | n210 ;
  assign n4392 = n808 | n4391 ;
  assign n4393 = n2923 | n4392 ;
  assign n4394 = n4390 | n4393 ;
  assign n4395 = n261 | n431 ;
  assign n4396 = n758 | n4395 ;
  assign n4397 = n144 | n524 ;
  assign n4398 = n1124 | n4397 ;
  assign n4399 = n4396 | n4398 ;
  assign n4400 = n3032 | n4399 ;
  assign n4401 = n705 | n1440 ;
  assign n4402 = n4400 | n4401 ;
  assign n4403 = n4394 | n4402 ;
  assign n4404 = n997 | n1637 ;
  assign n4405 = n125 | n174 ;
  assign n4406 = n82 | n4405 ;
  assign n4407 = n4404 | n4406 ;
  assign n4408 = n305 | n742 ;
  assign n4409 = n184 | n593 ;
  assign n4410 = n2592 | n4409 ;
  assign n4411 = n4408 | n4410 ;
  assign n4412 = n1308 | n2452 ;
  assign n4413 = n4411 | n4412 ;
  assign n4414 = n4407 | n4413 ;
  assign n4415 = n4403 | n4414 ;
  assign n4416 = n4388 | n4415 ;
  assign n4417 = n795 | n1590 ;
  assign n4418 = n2647 | n2744 ;
  assign n4419 = n4417 | n4418 ;
  assign n4420 = n4300 | n4419 ;
  assign n4421 = n368 | n493 ;
  assign n4422 = n294 | n4421 ;
  assign n4423 = n3355 | n4422 ;
  assign n4424 = n4420 | n4423 ;
  assign n4425 = n321 | n617 ;
  assign n4426 = n1860 | n4425 ;
  assign n4427 = n2051 | n4426 ;
  assign n4428 = n703 | n4427 ;
  assign n4429 = n4424 | n4428 ;
  assign n4430 = n305 | n441 ;
  assign n4431 = n2890 | n4430 ;
  assign n4432 = n480 | n977 ;
  assign n4433 = n4431 | n4432 ;
  assign n4434 = n174 | n350 ;
  assign n4435 = n860 | n4434 ;
  assign n4436 = n202 | n4435 ;
  assign n4437 = n4433 | n4436 ;
  assign n4438 = n4429 | n4437 ;
  assign n4439 = n711 | n969 ;
  assign n4440 = n440 | n1462 ;
  assign n4441 = n4439 | n4440 ;
  assign n4442 = n4120 | n4441 ;
  assign n4443 = n402 | n432 ;
  assign n4444 = n110 | n360 ;
  assign n4445 = n269 | n4444 ;
  assign n4446 = n4443 | n4445 ;
  assign n4447 = n1951 | n4446 ;
  assign n4448 = n133 | n442 ;
  assign n4449 = n257 | n623 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = n179 | n220 ;
  assign n4452 = n4450 | n4451 ;
  assign n4453 = n4447 | n4452 ;
  assign n4454 = n2803 | n4453 ;
  assign n4455 = n4442 | n4454 ;
  assign n4456 = n123 | n614 ;
  assign n4457 = n1345 | n4456 ;
  assign n4458 = n314 | n4457 ;
  assign n4459 = n2196 | n4458 ;
  assign n4460 = n285 | n297 ;
  assign n4461 = n1666 | n4460 ;
  assign n4462 = n3021 | n4461 ;
  assign n4463 = n1096 | n4462 ;
  assign n4464 = n4459 | n4463 ;
  assign n4465 = n164 | n392 ;
  assign n4466 = n618 & ~n4465 ;
  assign n4467 = ~n2775 & n4466 ;
  assign n4468 = ~n1752 & n4467 ;
  assign n4469 = n647 | n662 ;
  assign n4470 = n707 | n4469 ;
  assign n4471 = n323 | n912 ;
  assign n4472 = n1626 | n4471 ;
  assign n4473 = n4470 | n4472 ;
  assign n4474 = n4468 & ~n4473 ;
  assign n4475 = n358 | n404 ;
  assign n4476 = n747 | n1184 ;
  assign n4477 = n4475 | n4476 ;
  assign n4478 = n1437 | n1926 ;
  assign n4479 = n4477 | n4478 ;
  assign n4480 = n80 | n278 ;
  assign n4481 = n334 | n674 ;
  assign n4482 = n4480 | n4481 ;
  assign n4483 = n4479 | n4482 ;
  assign n4484 = n4474 & ~n4483 ;
  assign n4485 = ~n4464 & n4484 ;
  assign n4486 = ~n4455 & n4485 ;
  assign n4487 = ~n4438 & n4486 ;
  assign n4488 = ( x14 & ~n4416 ) | ( x14 & n4487 ) | ( ~n4416 & n4487 ) ;
  assign n4489 = n2795 | n3042 ;
  assign n4490 = n334 | n623 ;
  assign n4491 = n2307 | n4490 ;
  assign n4492 = n4489 | n4491 ;
  assign n4493 = n206 | n269 ;
  assign n4494 = n3754 | n4493 ;
  assign n4495 = n131 | n989 ;
  assign n4496 = n2863 | n4495 ;
  assign n4497 = n4494 | n4496 ;
  assign n4498 = n279 | n342 ;
  assign n4499 = n617 | n4498 ;
  assign n4500 = n1287 | n4499 ;
  assign n4501 = n4497 | n4500 ;
  assign n4502 = n2428 | n2979 ;
  assign n4503 = n316 | n4502 ;
  assign n4504 = n4501 | n4503 ;
  assign n4505 = n4492 | n4504 ;
  assign n4506 = n4394 | n4505 ;
  assign n4507 = n356 | n455 ;
  assign n4508 = n2781 | n4507 ;
  assign n4509 = n215 | n306 ;
  assign n4510 = n527 | n4509 ;
  assign n4511 = n4508 | n4510 ;
  assign n4512 = n87 | n4511 ;
  assign n4513 = n522 | n1066 ;
  assign n4514 = n330 | n4366 ;
  assign n4515 = n4513 | n4514 ;
  assign n4516 = n4512 | n4515 ;
  assign n4517 = n2513 | n4431 ;
  assign n4518 = n4516 | n4517 ;
  assign n4519 = n4506 | n4518 ;
  assign n4520 = n3629 | n4519 ;
  assign n4521 = ( n4338 & n4488 ) | ( n4338 & ~n4520 ) | ( n4488 & ~n4520 ) ;
  assign n4522 = ( n4268 & n4338 ) | ( n4268 & ~n4521 ) | ( n4338 & ~n4521 ) ;
  assign n4523 = ~n1529 & n3270 ;
  assign n4524 = n1687 & n3273 ;
  assign n4525 = n4523 | n4524 ;
  assign n4526 = n1600 & n3274 ;
  assign n4527 = n4525 | n4526 ;
  assign n4528 = n390 | n4527 ;
  assign n4529 = n3145 & n3255 ;
  assign n4530 = ~n3144 & n3256 ;
  assign n4531 = ( n1529 & ~n4529 ) | ( n1529 & n4530 ) | ( ~n4529 & n4530 ) ;
  assign n4532 = ( n4527 & n4528 ) | ( n4527 & ~n4531 ) | ( n4528 & ~n4531 ) ;
  assign n4533 = ( x17 & ~n4268 ) | ( x17 & n4314 ) | ( ~n4268 & n4314 ) ;
  assign n4534 = ( ~x17 & n4315 ) | ( ~x17 & n4533 ) | ( n4315 & n4533 ) ;
  assign n4535 = ( n4522 & n4532 ) | ( n4522 & n4534 ) | ( n4532 & n4534 ) ;
  assign n4536 = ~n1118 & n4039 ;
  assign n4537 = ~n1207 & n3501 ;
  assign n4538 = n4536 | n4537 ;
  assign n4539 = n1316 & n3536 ;
  assign n4540 = n4538 | n4539 ;
  assign n4541 = n3541 | n4540 ;
  assign n4542 = ( n3841 & n4540 ) | ( n3841 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4543 = x29 & ~n4542 ;
  assign n4544 = ~x29 & n4542 ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = ( n3904 & n4315 ) | ( n3904 & n4325 ) | ( n4315 & n4325 ) ;
  assign n4547 = ( n4325 & n4326 ) | ( n4325 & ~n4546 ) | ( n4326 & ~n4546 ) ;
  assign n4548 = ( n4535 & n4545 ) | ( n4535 & n4547 ) | ( n4545 & n4547 ) ;
  assign n4549 = ( n3904 & n4091 ) | ( n3904 & ~n4152 ) | ( n4091 & ~n4152 ) ;
  assign n4550 = ( ~n3904 & n4153 ) | ( ~n3904 & n4549 ) | ( n4153 & n4549 ) ;
  assign n4551 = ( ~n4326 & n4548 ) | ( ~n4326 & n4550 ) | ( n4548 & n4550 ) ;
  assign n4552 = ~n1118 & n3536 ;
  assign n4553 = n859 & n4039 ;
  assign n4554 = n4552 | n4553 ;
  assign n4555 = n995 & n3501 ;
  assign n4556 = n4554 | n4555 ;
  assign n4557 = n3541 | n4556 ;
  assign n4558 = ( ~n4034 & n4556 ) | ( ~n4034 & n4557 ) | ( n4556 & n4557 ) ;
  assign n4559 = x29 & ~n4558 ;
  assign n4560 = ~x29 & n4558 ;
  assign n4561 = n4559 | n4560 ;
  assign n4562 = ( n4153 & n4164 ) | ( n4153 & ~n4166 ) | ( n4164 & ~n4166 ) ;
  assign n4563 = ( ~n4153 & n4167 ) | ( ~n4153 & n4562 ) | ( n4167 & n4562 ) ;
  assign n4564 = ( n4551 & n4561 ) | ( n4551 & n4563 ) | ( n4561 & n4563 ) ;
  assign n4565 = ~n3487 & n4200 ;
  assign n4566 = ~n3601 & n4215 ;
  assign n4567 = ~n564 & n2083 ;
  assign n4568 = ( n2083 & n4566 ) | ( n2083 & ~n4567 ) | ( n4566 & ~n4567 ) ;
  assign n4569 = n4565 | n4568 ;
  assign n4570 = n4203 | n4569 ;
  assign n4571 = ( n3674 & n4569 ) | ( n3674 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = x26 & ~n4571 ;
  assign n4573 = ~x26 & n4571 ;
  assign n4574 = n4572 | n4573 ;
  assign n4575 = ( ~n4080 & n4167 ) | ( ~n4080 & n4169 ) | ( n4167 & n4169 ) ;
  assign n4576 = ( ~n4169 & n4170 ) | ( ~n4169 & n4575 ) | ( n4170 & n4575 ) ;
  assign n4577 = ( n4564 & n4574 ) | ( n4564 & ~n4576 ) | ( n4574 & ~n4576 ) ;
  assign n4578 = x20 | x22 ;
  assign n4579 = x21 | n4578 ;
  assign n4580 = x23 & ~n4579 ;
  assign n4581 = x21 & x22 ;
  assign n4582 = x20 & ~x23 ;
  assign n4583 = n4581 & n4582 ;
  assign n4584 = n4580 | n4583 ;
  assign n4585 = x22 & x23 ;
  assign n4586 = x22 | x23 ;
  assign n4587 = ~n4585 & n4586 ;
  assign n4588 = x20 & x21 ;
  assign n4589 = ~x20 & x21 ;
  assign n4590 = ( x20 & ~n4588 ) | ( x20 & n4589 ) | ( ~n4588 & n4589 ) ;
  assign n4591 = n4587 & n4590 ;
  assign n4592 = ( ~n3516 & n3608 ) | ( ~n3516 & n4591 ) | ( n3608 & n4591 ) ;
  assign n4593 = ( ~n3607 & n4584 ) | ( ~n3607 & n4592 ) | ( n4584 & n4592 ) ;
  assign n4594 = x23 & ~n4593 ;
  assign n4595 = ~x23 & n4593 ;
  assign n4596 = n4594 | n4595 ;
  assign n4597 = ( ~n4213 & n4227 ) | ( ~n4213 & n4237 ) | ( n4227 & n4237 ) ;
  assign n4598 = ( n4213 & ~n4238 ) | ( n4213 & n4597 ) | ( ~n4238 & n4597 ) ;
  assign n4599 = ( n4577 & n4596 ) | ( n4577 & n4598 ) | ( n4596 & n4598 ) ;
  assign n4600 = n564 & n4215 ;
  assign n4601 = ~n721 & n4200 ;
  assign n4602 = n4600 | n4601 ;
  assign n4603 = n859 & n2083 ;
  assign n4604 = n4602 | n4603 ;
  assign n4605 = n4203 | n4604 ;
  assign n4606 = ( ~n3268 & n4604 ) | ( ~n3268 & n4605 ) | ( n4604 & n4605 ) ;
  assign n4607 = x26 & ~n4606 ;
  assign n4608 = ~x26 & n4606 ;
  assign n4609 = n4607 | n4608 ;
  assign n4610 = n995 & n4039 ;
  assign n4611 = ~n1207 & n3536 ;
  assign n4612 = n4610 | n4611 ;
  assign n4613 = ~n1118 & n3501 ;
  assign n4614 = n4612 | n4613 ;
  assign n4615 = n3541 | n4614 ;
  assign n4616 = ( n4173 & n4614 ) | ( n4173 & n4615 ) | ( n4614 & n4615 ) ;
  assign n4617 = x29 & ~n4616 ;
  assign n4618 = ~x29 & n4616 ;
  assign n4619 = n4617 | n4618 ;
  assign n4620 = ( n4326 & n4548 ) | ( n4326 & n4550 ) | ( n4548 & n4550 ) ;
  assign n4621 = ( n4326 & n4551 ) | ( n4326 & ~n4620 ) | ( n4551 & ~n4620 ) ;
  assign n4622 = ( n4609 & n4619 ) | ( n4609 & ~n4621 ) | ( n4619 & ~n4621 ) ;
  assign n4623 = ( ~n4551 & n4561 ) | ( ~n4551 & n4563 ) | ( n4561 & n4563 ) ;
  assign n4624 = ( n4551 & ~n4564 ) | ( n4551 & n4623 ) | ( ~n4564 & n4623 ) ;
  assign n4625 = ~n3487 & n4215 ;
  assign n4626 = ~n721 & n2083 ;
  assign n4627 = n564 & n4200 ;
  assign n4628 = n4626 | n4627 ;
  assign n4629 = n4625 | n4628 ;
  assign n4630 = n4203 | n4629 ;
  assign n4631 = ( ~n3492 & n4629 ) | ( ~n3492 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4632 = x26 & ~n4631 ;
  assign n4633 = ~x26 & n4631 ;
  assign n4634 = n4632 | n4633 ;
  assign n4635 = ( n4622 & n4624 ) | ( n4622 & n4634 ) | ( n4624 & n4634 ) ;
  assign n4636 = n4578 & ~n4581 ;
  assign n4637 = ~n4590 & n4636 ;
  assign n4638 = ~n3516 & n4637 ;
  assign n4639 = x23 & n4638 ;
  assign n4640 = ~n3533 & n4584 ;
  assign n4641 = n4591 | n4640 ;
  assign n4642 = ( n3609 & n4640 ) | ( n3609 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4643 = x23 & ~n4642 ;
  assign n4644 = ( ~x23 & n4638 ) | ( ~x23 & n4642 ) | ( n4638 & n4642 ) ;
  assign n4645 = ( ~n4639 & n4643 ) | ( ~n4639 & n4644 ) | ( n4643 & n4644 ) ;
  assign n4646 = ( ~n4564 & n4574 ) | ( ~n4564 & n4576 ) | ( n4574 & n4576 ) ;
  assign n4647 = ( ~n4574 & n4577 ) | ( ~n4574 & n4646 ) | ( n4577 & n4646 ) ;
  assign n4648 = ( n4635 & n4645 ) | ( n4635 & ~n4647 ) | ( n4645 & ~n4647 ) ;
  assign n4649 = ~n4587 & n4590 ;
  assign n4650 = ~n3533 & n4649 ;
  assign n4651 = x23 & n4650 ;
  assign n4652 = ~n3601 & n4637 ;
  assign n4653 = ~n3487 & n4584 ;
  assign n4654 = n4652 | n4653 ;
  assign n4655 = n4591 | n4654 ;
  assign n4656 = ( ~n4223 & n4654 ) | ( ~n4223 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = x23 & ~n4656 ;
  assign n4658 = ( ~x23 & n4650 ) | ( ~x23 & n4656 ) | ( n4650 & n4656 ) ;
  assign n4659 = ( ~n4651 & n4657 ) | ( ~n4651 & n4658 ) | ( n4657 & n4658 ) ;
  assign n4660 = ~n1529 & n3536 ;
  assign n4661 = x29 & n4660 ;
  assign n4662 = n1316 & n4039 ;
  assign n4663 = n1398 & n3501 ;
  assign n4664 = n4662 | n4663 ;
  assign n4665 = n3541 | n4664 ;
  assign n4666 = ( n4084 & n4664 ) | ( n4084 & n4665 ) | ( n4664 & n4665 ) ;
  assign n4667 = x29 & ~n4666 ;
  assign n4668 = ( ~x29 & n4660 ) | ( ~x29 & n4666 ) | ( n4660 & n4666 ) ;
  assign n4669 = ( ~n4661 & n4667 ) | ( ~n4661 & n4668 ) | ( n4667 & n4668 ) ;
  assign n4670 = ( ~n4268 & n4338 ) | ( ~n4268 & n4521 ) | ( n4338 & n4521 ) ;
  assign n4671 = ( ~n4338 & n4522 ) | ( ~n4338 & n4670 ) | ( n4522 & n4670 ) ;
  assign n4672 = n1600 & n3254 ;
  assign n4673 = ( n1600 & n3143 ) | ( n1600 & ~n3254 ) | ( n3143 & ~n3254 ) ;
  assign n4674 = ( ~n3144 & n4672 ) | ( ~n3144 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4675 = n1687 & n3274 ;
  assign n4676 = n1792 & n3273 ;
  assign n4677 = n1600 & n3270 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = n4675 | n4678 ;
  assign n4680 = n390 | n4679 ;
  assign n4681 = ( n4674 & n4679 ) | ( n4674 & n4680 ) | ( n4679 & n4680 ) ;
  assign n4682 = ( n4669 & ~n4671 ) | ( n4669 & n4681 ) | ( ~n4671 & n4681 ) ;
  assign n4683 = ( ~n4522 & n4532 ) | ( ~n4522 & n4534 ) | ( n4532 & n4534 ) ;
  assign n4684 = ( n4522 & ~n4535 ) | ( n4522 & n4683 ) | ( ~n4535 & n4683 ) ;
  assign n4685 = n1316 & n3501 ;
  assign n4686 = ~n1207 & n4039 ;
  assign n4687 = n1398 & n3536 ;
  assign n4688 = n4686 | n4687 ;
  assign n4689 = n4685 | n4688 ;
  assign n4690 = n3541 | n4689 ;
  assign n4691 = ( ~n4157 & n4689 ) | ( ~n4157 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4692 = x29 & ~n4691 ;
  assign n4693 = ~x29 & n4691 ;
  assign n4694 = n4692 | n4693 ;
  assign n4695 = ( n4682 & n4684 ) | ( n4682 & n4694 ) | ( n4684 & n4694 ) ;
  assign n4696 = n859 & n4200 ;
  assign n4697 = ~n721 & n4215 ;
  assign n4698 = n4696 | n4697 ;
  assign n4699 = n995 & n2083 ;
  assign n4700 = n4698 | n4699 ;
  assign n4701 = n4203 | n4700 ;
  assign n4702 = ( ~n3829 & n4700 ) | ( ~n3829 & n4701 ) | ( n4700 & n4701 ) ;
  assign n4703 = x26 & ~n4702 ;
  assign n4704 = ~x26 & n4702 ;
  assign n4705 = n4703 | n4704 ;
  assign n4706 = ( ~n4535 & n4545 ) | ( ~n4535 & n4547 ) | ( n4545 & n4547 ) ;
  assign n4707 = ( n4535 & ~n4548 ) | ( n4535 & n4706 ) | ( ~n4548 & n4706 ) ;
  assign n4708 = ( n4695 & n4705 ) | ( n4695 & n4707 ) | ( n4705 & n4707 ) ;
  assign n4709 = ( n4609 & ~n4619 ) | ( n4609 & n4621 ) | ( ~n4619 & n4621 ) ;
  assign n4710 = ( ~n4609 & n4622 ) | ( ~n4609 & n4709 ) | ( n4622 & n4709 ) ;
  assign n4711 = ( n4659 & n4708 ) | ( n4659 & ~n4710 ) | ( n4708 & ~n4710 ) ;
  assign n4712 = ( n4622 & ~n4624 ) | ( n4622 & n4634 ) | ( ~n4624 & n4634 ) ;
  assign n4713 = ( n4624 & ~n4635 ) | ( n4624 & n4712 ) | ( ~n4635 & n4712 ) ;
  assign n4714 = ~n3533 & n4637 ;
  assign n4715 = x23 & n4714 ;
  assign n4716 = ~n3516 & n4649 ;
  assign n4717 = n4584 | n4716 ;
  assign n4718 = ( ~n3601 & n4716 ) | ( ~n3601 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4719 = n4591 | n4718 ;
  assign n4720 = ( ~n4058 & n4718 ) | ( ~n4058 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4721 = x23 & ~n4720 ;
  assign n4722 = ( ~x23 & n4714 ) | ( ~x23 & n4720 ) | ( n4714 & n4720 ) ;
  assign n4723 = ( ~n4715 & n4721 ) | ( ~n4715 & n4722 ) | ( n4721 & n4722 ) ;
  assign n4724 = ( n4711 & n4713 ) | ( n4711 & n4723 ) | ( n4713 & n4723 ) ;
  assign n4725 = n995 & n4215 ;
  assign n4726 = ~n1207 & n2083 ;
  assign n4727 = n4725 | n4726 ;
  assign n4728 = ~n1118 & n4200 ;
  assign n4729 = n4727 | n4728 ;
  assign n4730 = n4203 | n4729 ;
  assign n4731 = ( n4173 & n4729 ) | ( n4173 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4732 = x26 & ~n4731 ;
  assign n4733 = ~x26 & n4731 ;
  assign n4734 = n4732 | n4733 ;
  assign n4735 = ~n1529 & n3501 ;
  assign n4736 = n1600 & n3536 ;
  assign n4737 = n1398 & n4039 ;
  assign n4738 = n4736 | n4737 ;
  assign n4739 = n4735 | n4738 ;
  assign n4740 = x29 & n4739 ;
  assign n4741 = n3541 & ~n4324 ;
  assign n4742 = x29 & ~n4741 ;
  assign n4743 = ( ~x29 & n4739 ) | ( ~x29 & n4741 ) | ( n4739 & n4741 ) ;
  assign n4744 = ( ~n4740 & n4742 ) | ( ~n4740 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4745 = ~n1841 & n3270 ;
  assign n4746 = ~n2041 & n3273 ;
  assign n4747 = n4745 | n4746 ;
  assign n4748 = n1943 & n3274 ;
  assign n4749 = n4747 | n4748 ;
  assign n4750 = n390 | n4749 ;
  assign n4751 = n3141 & n3251 ;
  assign n4752 = ~n3140 & n3252 ;
  assign n4753 = ( n1841 & ~n4751 ) | ( n1841 & n4752 ) | ( ~n4751 & n4752 ) ;
  assign n4754 = ( n4749 & n4750 ) | ( n4749 & ~n4753 ) | ( n4750 & ~n4753 ) ;
  assign n4755 = n334 | n986 ;
  assign n4756 = n794 | n912 ;
  assign n4757 = n2276 | n4756 ;
  assign n4758 = n4755 | n4757 ;
  assign n4759 = n150 | n656 ;
  assign n4760 = n322 | n613 ;
  assign n4761 = n678 | n1020 ;
  assign n4762 = n4760 | n4761 ;
  assign n4763 = n4759 | n4762 ;
  assign n4764 = n4758 | n4763 ;
  assign n4765 = n2552 | n2870 ;
  assign n4766 = n661 | n4765 ;
  assign n4767 = n4764 | n4766 ;
  assign n4768 = n268 | n351 ;
  assign n4769 = n956 | n4768 ;
  assign n4770 = n816 | n4769 ;
  assign n4771 = n241 | n983 ;
  assign n4772 = n4770 | n4771 ;
  assign n4773 = n108 | n306 ;
  assign n4774 = n3994 | n4773 ;
  assign n4775 = n1429 | n4774 ;
  assign n4776 = n163 | n379 ;
  assign n4777 = n4775 | n4776 ;
  assign n4778 = n432 | n916 ;
  assign n4779 = n480 | n4778 ;
  assign n4780 = n2421 | n4779 ;
  assign n4781 = n148 | n441 ;
  assign n4782 = n1253 | n4781 ;
  assign n4783 = n2898 | n4782 ;
  assign n4784 = n4780 | n4783 ;
  assign n4785 = n4777 | n4784 ;
  assign n4786 = n4772 | n4785 ;
  assign n4787 = n4767 | n4786 ;
  assign n4788 = n303 | n535 ;
  assign n4789 = n3355 | n4788 ;
  assign n4790 = n1642 | n2719 ;
  assign n4791 = n4789 | n4790 ;
  assign n4792 = n3287 | n4791 ;
  assign n4793 = n1193 | n1586 ;
  assign n4794 = n298 | n1617 ;
  assign n4795 = n4793 | n4794 ;
  assign n4796 = n260 | n434 ;
  assign n4797 = n226 | n4796 ;
  assign n4798 = n4795 | n4797 ;
  assign n4799 = n3367 | n3395 ;
  assign n4800 = n3853 | n4799 ;
  assign n4801 = n4798 | n4800 ;
  assign n4802 = n4792 | n4801 ;
  assign n4803 = n4787 | n4802 ;
  assign n4804 = n210 | n999 ;
  assign n4805 = n1162 | n4804 ;
  assign n4806 = n269 | n704 ;
  assign n4807 = n4375 | n4806 ;
  assign n4808 = n1560 | n4253 ;
  assign n4809 = n4807 | n4808 ;
  assign n4810 = n4805 | n4809 ;
  assign n4811 = n291 | n2332 ;
  assign n4812 = n3686 | n4811 ;
  assign n4813 = n4810 | n4812 ;
  assign n4814 = n643 | n1150 ;
  assign n4815 = n4813 | n4814 ;
  assign n4816 = n368 | n922 ;
  assign n4817 = n508 | n1786 ;
  assign n4818 = n428 | n1332 ;
  assign n4819 = n4817 | n4818 ;
  assign n4820 = n4816 | n4819 ;
  assign n4821 = n4815 | n4820 ;
  assign n4822 = n4803 | n4821 ;
  assign n4823 = ( ~n4416 & n4754 ) | ( ~n4416 & n4822 ) | ( n4754 & n4822 ) ;
  assign n4824 = n1943 & n3273 ;
  assign n4825 = n1792 & n3270 ;
  assign n4826 = n4824 | n4825 ;
  assign n4827 = ~n1841 & n3274 ;
  assign n4828 = n4826 | n4827 ;
  assign n4829 = n390 | n4828 ;
  assign n4830 = n1792 & n3252 ;
  assign n4831 = ( n3142 & n4328 ) | ( n3142 & ~n4830 ) | ( n4328 & ~n4830 ) ;
  assign n4832 = ( n4828 & n4829 ) | ( n4828 & ~n4831 ) | ( n4829 & ~n4831 ) ;
  assign n4833 = ( x14 & n4416 ) | ( x14 & ~n4487 ) | ( n4416 & ~n4487 ) ;
  assign n4834 = ( ~x14 & n4488 ) | ( ~x14 & n4833 ) | ( n4488 & n4833 ) ;
  assign n4835 = ( n4823 & n4832 ) | ( n4823 & n4834 ) | ( n4832 & n4834 ) ;
  assign n4836 = ( n4338 & n4488 ) | ( n4338 & n4520 ) | ( n4488 & n4520 ) ;
  assign n4837 = ( n4520 & n4521 ) | ( n4520 & ~n4836 ) | ( n4521 & ~n4836 ) ;
  assign n4838 = ( n4744 & n4835 ) | ( n4744 & n4837 ) | ( n4835 & n4837 ) ;
  assign n4839 = ( n4669 & n4671 ) | ( n4669 & ~n4681 ) | ( n4671 & ~n4681 ) ;
  assign n4840 = ( ~n4669 & n4682 ) | ( ~n4669 & n4839 ) | ( n4682 & n4839 ) ;
  assign n4841 = ( n4734 & n4838 ) | ( n4734 & ~n4840 ) | ( n4838 & ~n4840 ) ;
  assign n4842 = n859 & n4215 ;
  assign n4843 = n995 & n4200 ;
  assign n4844 = n4842 | n4843 ;
  assign n4845 = ~n1118 & n2083 ;
  assign n4846 = n4844 | n4845 ;
  assign n4847 = n4203 | n4846 ;
  assign n4848 = ( ~n4034 & n4846 ) | ( ~n4034 & n4847 ) | ( n4846 & n4847 ) ;
  assign n4849 = x26 & ~n4848 ;
  assign n4850 = ~x26 & n4848 ;
  assign n4851 = n4849 | n4850 ;
  assign n4852 = ( ~n4682 & n4684 ) | ( ~n4682 & n4694 ) | ( n4684 & n4694 ) ;
  assign n4853 = ( n4682 & ~n4695 ) | ( n4682 & n4852 ) | ( ~n4695 & n4852 ) ;
  assign n4854 = ( n4841 & n4851 ) | ( n4841 & n4853 ) | ( n4851 & n4853 ) ;
  assign n4855 = ( ~n4695 & n4705 ) | ( ~n4695 & n4707 ) | ( n4705 & n4707 ) ;
  assign n4856 = ( n4695 & ~n4708 ) | ( n4695 & n4855 ) | ( ~n4708 & n4855 ) ;
  assign n4857 = ~n3487 & n4637 ;
  assign n4858 = ~n3601 & n4649 ;
  assign n4859 = ~n564 & n4584 ;
  assign n4860 = ( n4584 & n4858 ) | ( n4584 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  assign n4861 = n4857 | n4860 ;
  assign n4862 = n4591 | n4861 ;
  assign n4863 = ( n3674 & n4861 ) | ( n3674 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4864 = x23 & ~n4863 ;
  assign n4865 = ~x23 & n4863 ;
  assign n4866 = n4864 | n4865 ;
  assign n4867 = ( n4854 & n4856 ) | ( n4854 & n4866 ) | ( n4856 & n4866 ) ;
  assign n4868 = x17 & x18 ;
  assign n4869 = x19 & n4868 ;
  assign n4870 = ~x20 & n4869 ;
  assign n4871 = x17 | x18 ;
  assign n4872 = x19 | n4871 ;
  assign n4873 = x20 & ~n4872 ;
  assign n4874 = n4870 | n4873 ;
  assign n4875 = ~n4868 & n4871 ;
  assign n4876 = x19 & x20 ;
  assign n4877 = x19 | x20 ;
  assign n4878 = ( n4875 & n4876 ) | ( n4875 & ~n4877 ) | ( n4876 & ~n4877 ) ;
  assign n4879 = n4875 & ~n4878 ;
  assign n4880 = ( ~n3516 & n3608 ) | ( ~n3516 & n4879 ) | ( n3608 & n4879 ) ;
  assign n4881 = ( ~n3607 & n4874 ) | ( ~n3607 & n4880 ) | ( n4874 & n4880 ) ;
  assign n4882 = x20 & ~n4881 ;
  assign n4883 = ~x20 & n4881 ;
  assign n4884 = n4882 | n4883 ;
  assign n4885 = ( n4659 & ~n4708 ) | ( n4659 & n4710 ) | ( ~n4708 & n4710 ) ;
  assign n4886 = ( ~n4659 & n4711 ) | ( ~n4659 & n4885 ) | ( n4711 & n4885 ) ;
  assign n4887 = ( n4867 & n4884 ) | ( n4867 & ~n4886 ) | ( n4884 & ~n4886 ) ;
  assign n4888 = n192 | n942 ;
  assign n4889 = n1020 | n4888 ;
  assign n4890 = n1421 | n4889 ;
  assign n4891 = n256 | n567 ;
  assign n4892 = n405 | n4891 ;
  assign n4893 = n4890 | n4892 ;
  assign n4894 = n2866 | n3072 ;
  assign n4895 = n378 | n431 ;
  assign n4896 = n321 | n4895 ;
  assign n4897 = n48 | n3623 ;
  assign n4898 = n4896 | n4897 ;
  assign n4899 = n4894 | n4898 ;
  assign n4900 = n4893 | n4899 ;
  assign n4901 = n2160 | n4900 ;
  assign n4902 = n83 | n2964 ;
  assign n4903 = n3448 | n4469 ;
  assign n4904 = n290 | n347 ;
  assign n4905 = n4903 | n4904 ;
  assign n4906 = n4902 | n4905 ;
  assign n4907 = n674 | n1332 ;
  assign n4908 = n591 | n4907 ;
  assign n4909 = n4759 | n4908 ;
  assign n4910 = n844 | n3433 ;
  assign n4911 = n4909 | n4910 ;
  assign n4912 = n4906 | n4911 ;
  assign n4913 = n4344 | n4912 ;
  assign n4914 = n4901 | n4913 ;
  assign n4915 = n1117 | n4914 ;
  assign n4916 = n275 | n1048 ;
  assign n4917 = n742 | n4916 ;
  assign n4918 = n456 | n533 ;
  assign n4919 = n463 | n4918 ;
  assign n4920 = n613 | n1176 ;
  assign n4921 = n3791 | n4920 ;
  assign n4922 = n4919 | n4921 ;
  assign n4923 = n4917 | n4922 ;
  assign n4924 = n2317 | n3323 ;
  assign n4925 = n4359 | n4924 ;
  assign n4926 = n4923 | n4925 ;
  assign n4927 = n153 | n294 ;
  assign n4928 = n2479 | n4927 ;
  assign n4929 = n99 | n659 ;
  assign n4930 = n2222 | n4929 ;
  assign n4931 = n4928 | n4930 ;
  assign n4932 = n272 | n4931 ;
  assign n4933 = n4926 | n4932 ;
  assign n4934 = n4915 | n4933 ;
  assign n4935 = n3698 | n3890 ;
  assign n4936 = n4912 | n4935 ;
  assign n4937 = n449 | n628 ;
  assign n4938 = n2704 | n3995 ;
  assign n4939 = n4937 | n4938 ;
  assign n4940 = n850 | n1094 ;
  assign n4941 = n125 | n4940 ;
  assign n4942 = n358 | n2062 ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = n4939 | n4943 ;
  assign n4945 = n983 | n2611 ;
  assign n4946 = n1699 | n4945 ;
  assign n4947 = n4944 | n4946 ;
  assign n4948 = n2072 | n3446 ;
  assign n4949 = n454 | n922 ;
  assign n4950 = n4948 | n4949 ;
  assign n4951 = n279 | n659 ;
  assign n4952 = n97 | n4951 ;
  assign n4953 = n1048 | n4952 ;
  assign n4954 = n4950 | n4953 ;
  assign n4955 = n4947 | n4954 ;
  assign n4956 = n4936 | n4955 ;
  assign n4957 = n328 | n593 ;
  assign n4958 = n497 | n4957 ;
  assign n4959 = n70 | n238 ;
  assign n4960 = n3994 | n4959 ;
  assign n4961 = n4958 | n4960 ;
  assign n4962 = n133 | n197 ;
  assign n4963 = n700 | n942 ;
  assign n4964 = n4962 | n4963 ;
  assign n4965 = n4961 | n4964 ;
  assign n4966 = n2936 | n4965 ;
  assign n4967 = n218 | n360 ;
  assign n4968 = n368 | n4967 ;
  assign n4969 = n380 | n1872 ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = n3951 | n4460 ;
  assign n4972 = n2728 | n4971 ;
  assign n4973 = n2204 | n4972 ;
  assign n4974 = n4970 | n4973 ;
  assign n4975 = n1363 | n4974 ;
  assign n4976 = n4966 | n4975 ;
  assign n4977 = n413 | n3786 ;
  assign n4978 = n2189 | n4977 ;
  assign n4979 = n3657 | n4978 ;
  assign n4980 = n4976 | n4979 ;
  assign n4981 = n4956 | n4980 ;
  assign n4982 = ( ~x11 & n4934 ) | ( ~x11 & n4981 ) | ( n4934 & n4981 ) ;
  assign n4983 = n1943 & n3250 ;
  assign n4984 = ( ~n1943 & n3139 ) | ( ~n1943 & n3250 ) | ( n3139 & n3250 ) ;
  assign n4985 = ( n3140 & ~n4983 ) | ( n3140 & n4984 ) | ( ~n4983 & n4984 ) ;
  assign n4986 = n1943 & n3270 ;
  assign n4987 = ~n2041 & n3274 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = n2102 & n3273 ;
  assign n4990 = n4988 | n4989 ;
  assign n4991 = n390 | n4990 ;
  assign n4992 = ( ~n4985 & n4990 ) | ( ~n4985 & n4991 ) | ( n4990 & n4991 ) ;
  assign n4993 = ( ~n4416 & n4982 ) | ( ~n4416 & n4992 ) | ( n4982 & n4992 ) ;
  assign n4994 = n2041 | n3249 ;
  assign n4995 = ( n2041 & n3138 ) | ( n2041 & ~n3249 ) | ( n3138 & ~n3249 ) ;
  assign n4996 = n2041 | n3138 ;
  assign n4997 = ( n4994 & n4995 ) | ( n4994 & ~n4996 ) | ( n4995 & ~n4996 ) ;
  assign n4998 = n2102 & n3274 ;
  assign n4999 = ~n2041 & n3270 ;
  assign n5000 = n4998 | n4999 ;
  assign n5001 = n2187 & n3273 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = n390 | n5002 ;
  assign n5004 = ( ~n4997 & n5002 ) | ( ~n4997 & n5003 ) | ( n5002 & n5003 ) ;
  assign n5005 = ( x11 & n4934 ) | ( x11 & n4981 ) | ( n4934 & n4981 ) ;
  assign n5006 = ( x11 & n4982 ) | ( x11 & ~n5005 ) | ( n4982 & ~n5005 ) ;
  assign n5007 = n47 | n428 ;
  assign n5008 = n1323 | n3475 ;
  assign n5009 = n5007 | n5008 ;
  assign n5010 = n357 | n550 ;
  assign n5011 = n276 | n5010 ;
  assign n5012 = n1732 | n5011 ;
  assign n5013 = n5009 | n5012 ;
  assign n5014 = n1879 | n5013 ;
  assign n5015 = n662 | n863 ;
  assign n5016 = n4493 | n5015 ;
  assign n5017 = n2346 | n2717 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = n5014 | n5018 ;
  assign n5020 = n700 | n1074 ;
  assign n5021 = n351 | n5020 ;
  assign n5022 = n2553 & ~n2821 ;
  assign n5023 = ~n5021 & n5022 ;
  assign n5024 = n201 | n1126 ;
  assign n5025 = n5023 & ~n5024 ;
  assign n5026 = ~n3766 & n5025 ;
  assign n5027 = n177 | n2872 ;
  assign n5028 = n1612 | n5027 ;
  assign n5029 = n5026 & ~n5028 ;
  assign n5030 = ~n5019 & n5029 ;
  assign n5031 = n477 | n695 ;
  assign n5032 = n321 | n5031 ;
  assign n5033 = n3373 | n5032 ;
  assign n5034 = n378 | n600 ;
  assign n5035 = n4937 | n5034 ;
  assign n5036 = n5033 | n5035 ;
  assign n5037 = n1385 | n4977 ;
  assign n5038 = n5036 | n5037 ;
  assign n5039 = n465 | n2601 ;
  assign n5040 = n4471 | n5039 ;
  assign n5041 = n3073 | n5040 ;
  assign n5042 = n5038 | n5041 ;
  assign n5043 = n5030 & ~n5042 ;
  assign n5044 = n2918 | n3857 ;
  assign n5045 = n215 | n244 ;
  assign n5046 = n2059 | n5045 ;
  assign n5047 = n5044 | n5046 ;
  assign n5048 = n4459 | n5047 ;
  assign n5049 = n2348 | n3791 ;
  assign n5050 = n2659 | n5049 ;
  assign n5051 = n1737 | n2303 ;
  assign n5052 = n5050 | n5051 ;
  assign n5053 = n207 | n361 ;
  assign n5054 = n1678 | n5053 ;
  assign n5055 = n5052 | n5054 ;
  assign n5056 = n5048 | n5055 ;
  assign n5057 = n397 | n419 ;
  assign n5058 = n987 | n5057 ;
  assign n5059 = n2678 | n5058 ;
  assign n5060 = n1756 | n3114 ;
  assign n5061 = n4951 | n5060 ;
  assign n5062 = n5059 | n5061 ;
  assign n5063 = n528 | n4816 ;
  assign n5064 = n794 | n968 ;
  assign n5065 = n2834 | n5064 ;
  assign n5066 = n5063 | n5065 ;
  assign n5067 = n2314 | n5066 ;
  assign n5068 = n5062 | n5067 ;
  assign n5069 = n5056 | n5068 ;
  assign n5070 = n5043 & ~n5069 ;
  assign n5071 = n1094 | n1332 ;
  assign n5072 = n4443 | n5071 ;
  assign n5073 = n306 | n556 ;
  assign n5074 = n1862 | n5073 ;
  assign n5075 = n5072 | n5074 ;
  assign n5076 = n222 | n574 ;
  assign n5077 = n5075 | n5076 ;
  assign n5078 = n435 | n969 ;
  assign n5079 = n91 | n3192 ;
  assign n5080 = n5078 | n5079 ;
  assign n5081 = n5077 | n5080 ;
  assign n5082 = n293 | n455 ;
  assign n5083 = n218 | n591 ;
  assign n5084 = n5082 | n5083 ;
  assign n5085 = n1853 | n5084 ;
  assign n5086 = n416 | n623 ;
  assign n5087 = n1351 | n5086 ;
  assign n5088 = n498 | n2156 ;
  assign n5089 = n5087 | n5088 ;
  assign n5090 = n5085 | n5089 ;
  assign n5091 = n5081 | n5090 ;
  assign n5092 = n3384 | n4460 ;
  assign n5093 = n449 | n679 ;
  assign n5094 = n5092 | n5093 ;
  assign n5095 = n4108 | n5094 ;
  assign n5096 = n284 | n1193 ;
  assign n5097 = n913 | n3078 ;
  assign n5098 = n5096 | n5097 ;
  assign n5099 = n5095 | n5098 ;
  assign n5100 = n5091 | n5099 ;
  assign n5101 = n4138 | n5100 ;
  assign n5102 = n674 | n723 ;
  assign n5103 = n644 | n5102 ;
  assign n5104 = n1005 | n3365 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = n1272 | n1323 ;
  assign n5107 = n1589 | n5106 ;
  assign n5108 = n275 | n567 ;
  assign n5109 = n841 | n5108 ;
  assign n5110 = n2105 | n5109 ;
  assign n5111 = n5107 | n5110 ;
  assign n5112 = n5105 | n5111 ;
  assign n5113 = n1651 | n4469 ;
  assign n5114 = n1822 | n5113 ;
  assign n5115 = n3645 | n5114 ;
  assign n5116 = n4110 | n5115 ;
  assign n5117 = n148 | n210 ;
  assign n5118 = n4444 | n5117 ;
  assign n5119 = n356 | n2825 ;
  assign n5120 = n5118 | n5119 ;
  assign n5121 = n140 | n276 ;
  assign n5122 = n892 | n5121 ;
  assign n5123 = n4002 | n5122 ;
  assign n5124 = n5120 | n5123 ;
  assign n5125 = n5116 | n5124 ;
  assign n5126 = n5112 | n5125 ;
  assign n5127 = n5101 | n5126 ;
  assign n5128 = ( x8 & n5070 ) | ( x8 & ~n5127 ) | ( n5070 & ~n5127 ) ;
  assign n5129 = ~n2364 & n3273 ;
  assign n5130 = n2187 & n3270 ;
  assign n5131 = n5129 | n5130 ;
  assign n5132 = ~n2282 & n3274 ;
  assign n5133 = n5131 | n5132 ;
  assign n5134 = n390 | n5133 ;
  assign n5135 = n3137 & ~n3247 ;
  assign n5136 = n3136 & n3248 ;
  assign n5137 = ( n2187 & n5135 ) | ( n2187 & ~n5136 ) | ( n5135 & ~n5136 ) ;
  assign n5138 = ( n5133 & n5134 ) | ( n5133 & n5137 ) | ( n5134 & n5137 ) ;
  assign n5139 = ( n4934 & n5128 ) | ( n4934 & ~n5138 ) | ( n5128 & ~n5138 ) ;
  assign n5140 = n294 | n669 ;
  assign n5141 = n3360 | n5140 ;
  assign n5142 = n1048 | n2917 ;
  assign n5143 = n5141 | n5142 ;
  assign n5144 = n1578 | n2931 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = n3704 | n5145 ;
  assign n5147 = n2151 | n5146 ;
  assign n5148 = n2185 | n5147 ;
  assign n5149 = n1528 | n5148 ;
  assign n5150 = n556 | n623 ;
  assign n5151 = n356 | n554 ;
  assign n5152 = n5150 | n5151 ;
  assign n5153 = n1793 | n5152 ;
  assign n5154 = n261 | n308 ;
  assign n5155 = n280 | n5154 ;
  assign n5156 = n151 | n1006 ;
  assign n5157 = n271 | n5156 ;
  assign n5158 = n5155 | n5157 ;
  assign n5159 = n5153 | n5158 ;
  assign n5160 = n5149 | n5159 ;
  assign n5161 = ( n4934 & n5139 ) | ( n4934 & ~n5160 ) | ( n5139 & ~n5160 ) ;
  assign n5162 = ( ~n5004 & n5006 ) | ( ~n5004 & n5161 ) | ( n5006 & n5161 ) ;
  assign n5163 = ~n1841 & n3536 ;
  assign n5164 = n1687 & n4039 ;
  assign n5165 = n5163 | n5164 ;
  assign n5166 = n1792 & n3501 ;
  assign n5167 = n5165 | n5166 ;
  assign n5168 = x29 & n5167 ;
  assign n5169 = n3541 & n4331 ;
  assign n5170 = x29 & ~n5169 ;
  assign n5171 = ( ~x29 & n5167 ) | ( ~x29 & n5169 ) | ( n5167 & n5169 ) ;
  assign n5172 = ( ~n5168 & n5170 ) | ( ~n5168 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5173 = ( n4416 & n4982 ) | ( n4416 & n4992 ) | ( n4982 & n4992 ) ;
  assign n5174 = ( n4416 & n4993 ) | ( n4416 & ~n5173 ) | ( n4993 & ~n5173 ) ;
  assign n5175 = ( n5162 & ~n5172 ) | ( n5162 & n5174 ) | ( ~n5172 & n5174 ) ;
  assign n5176 = ( n4416 & n4754 ) | ( n4416 & n4822 ) | ( n4754 & n4822 ) ;
  assign n5177 = ( n4416 & n4823 ) | ( n4416 & ~n5176 ) | ( n4823 & ~n5176 ) ;
  assign n5178 = ( ~n4993 & n5175 ) | ( ~n4993 & n5177 ) | ( n5175 & n5177 ) ;
  assign n5179 = ~n1529 & n4039 ;
  assign n5180 = n1687 & n3536 ;
  assign n5181 = n5179 | n5180 ;
  assign n5182 = n1600 & n3501 ;
  assign n5183 = n5181 | n5182 ;
  assign n5184 = x29 & n5183 ;
  assign n5185 = n3541 & ~n4531 ;
  assign n5186 = x29 & ~n5185 ;
  assign n5187 = ( ~x29 & n5183 ) | ( ~x29 & n5185 ) | ( n5183 & n5185 ) ;
  assign n5188 = ( ~n5184 & n5186 ) | ( ~n5184 & n5187 ) | ( n5186 & n5187 ) ;
  assign n5189 = ( ~n4823 & n4832 ) | ( ~n4823 & n4834 ) | ( n4832 & n4834 ) ;
  assign n5190 = ( n4823 & ~n4835 ) | ( n4823 & n5189 ) | ( ~n4835 & n5189 ) ;
  assign n5191 = ( ~n5178 & n5188 ) | ( ~n5178 & n5190 ) | ( n5188 & n5190 ) ;
  assign n5192 = n1316 & n2083 ;
  assign n5193 = x26 & n5192 ;
  assign n5194 = ~n1118 & n4215 ;
  assign n5195 = ~n1207 & n4200 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = n4203 | n5196 ;
  assign n5198 = ( n3841 & n5196 ) | ( n3841 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5199 = x26 & ~n5198 ;
  assign n5200 = ( ~x26 & n5192 ) | ( ~x26 & n5198 ) | ( n5192 & n5198 ) ;
  assign n5201 = ( ~n5193 & n5199 ) | ( ~n5193 & n5200 ) | ( n5199 & n5200 ) ;
  assign n5202 = ( ~n4744 & n4835 ) | ( ~n4744 & n4837 ) | ( n4835 & n4837 ) ;
  assign n5203 = ( n4744 & ~n4838 ) | ( n4744 & n5202 ) | ( ~n4838 & n5202 ) ;
  assign n5204 = ( n5191 & n5201 ) | ( n5191 & n5203 ) | ( n5201 & n5203 ) ;
  assign n5205 = n564 & n4649 ;
  assign n5206 = n4591 | n5205 ;
  assign n5207 = ( ~n3268 & n5205 ) | ( ~n3268 & n5206 ) | ( n5205 & n5206 ) ;
  assign n5208 = n859 & n4584 ;
  assign n5209 = ( ~x23 & n5207 ) | ( ~x23 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5210 = ~n721 & n4637 ;
  assign n5211 = x23 & ~n5208 ;
  assign n5212 = n5210 | n5211 ;
  assign n5213 = ( n5207 & n5210 ) | ( n5207 & n5211 ) | ( n5210 & n5211 ) ;
  assign n5214 = ( n5209 & n5212 ) | ( n5209 & ~n5213 ) | ( n5212 & ~n5213 ) ;
  assign n5215 = ( n4734 & ~n4838 ) | ( n4734 & n4840 ) | ( ~n4838 & n4840 ) ;
  assign n5216 = ( ~n4734 & n4841 ) | ( ~n4734 & n5215 ) | ( n4841 & n5215 ) ;
  assign n5217 = ( n5204 & n5214 ) | ( n5204 & ~n5216 ) | ( n5214 & ~n5216 ) ;
  assign n5218 = ~n3487 & n4649 ;
  assign n5219 = ~n721 & n4584 ;
  assign n5220 = n564 & n4637 ;
  assign n5221 = n5219 | n5220 ;
  assign n5222 = n5218 | n5221 ;
  assign n5223 = n4591 | n5222 ;
  assign n5224 = ( ~n3492 & n5222 ) | ( ~n3492 & n5223 ) | ( n5222 & n5223 ) ;
  assign n5225 = x23 & ~n5224 ;
  assign n5226 = ~x23 & n5224 ;
  assign n5227 = n5225 | n5226 ;
  assign n5228 = ( ~n4841 & n4851 ) | ( ~n4841 & n4853 ) | ( n4851 & n4853 ) ;
  assign n5229 = ( n4841 & ~n4854 ) | ( n4841 & n5228 ) | ( ~n4854 & n5228 ) ;
  assign n5230 = ( n5217 & n5227 ) | ( n5217 & n5229 ) | ( n5227 & n5229 ) ;
  assign n5231 = n4872 & ~n4875 ;
  assign n5232 = ~n4869 & n5231 ;
  assign n5233 = ~n3516 & n5232 ;
  assign n5234 = x20 & n5233 ;
  assign n5235 = ~n3533 & n4874 ;
  assign n5236 = n4879 | n5235 ;
  assign n5237 = ( n3609 & n5235 ) | ( n3609 & n5236 ) | ( n5235 & n5236 ) ;
  assign n5238 = x20 & ~n5237 ;
  assign n5239 = ( ~x20 & n5233 ) | ( ~x20 & n5237 ) | ( n5233 & n5237 ) ;
  assign n5240 = ( ~n5234 & n5238 ) | ( ~n5234 & n5239 ) | ( n5238 & n5239 ) ;
  assign n5241 = ( ~n4854 & n4856 ) | ( ~n4854 & n4866 ) | ( n4856 & n4866 ) ;
  assign n5242 = ( n4854 & ~n4867 ) | ( n4854 & n5241 ) | ( ~n4867 & n5241 ) ;
  assign n5243 = ( n5230 & n5240 ) | ( n5230 & n5242 ) | ( n5240 & n5242 ) ;
  assign n5244 = ( ~n5217 & n5227 ) | ( ~n5217 & n5229 ) | ( n5227 & n5229 ) ;
  assign n5245 = ( n5217 & ~n5230 ) | ( n5217 & n5244 ) | ( ~n5230 & n5244 ) ;
  assign n5246 = ( ~n5191 & n5201 ) | ( ~n5191 & n5203 ) | ( n5201 & n5203 ) ;
  assign n5247 = ( n5191 & ~n5204 ) | ( n5191 & n5246 ) | ( ~n5204 & n5246 ) ;
  assign n5248 = n1316 & n4215 ;
  assign n5249 = n1398 & n4200 ;
  assign n5250 = n5248 | n5249 ;
  assign n5251 = ~n1529 & n2083 ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = x26 & n5252 ;
  assign n5254 = n4084 & n4203 ;
  assign n5255 = ( ~x26 & n5252 ) | ( ~x26 & n5254 ) | ( n5252 & n5254 ) ;
  assign n5256 = x26 & ~n5254 ;
  assign n5257 = ( ~n5253 & n5255 ) | ( ~n5253 & n5256 ) | ( n5255 & n5256 ) ;
  assign n5258 = n1687 & n3501 ;
  assign n5259 = n1600 & n4039 ;
  assign n5260 = n1792 & n3536 ;
  assign n5261 = n5259 | n5260 ;
  assign n5262 = n5258 | n5261 ;
  assign n5263 = n3541 | n5262 ;
  assign n5264 = ( n4674 & n5262 ) | ( n4674 & n5263 ) | ( n5262 & n5263 ) ;
  assign n5265 = x29 & ~n5264 ;
  assign n5266 = ~x29 & n5264 ;
  assign n5267 = n5265 | n5266 ;
  assign n5268 = ( n4993 & n5175 ) | ( n4993 & ~n5177 ) | ( n5175 & ~n5177 ) ;
  assign n5269 = ( ~n5175 & n5178 ) | ( ~n5175 & n5268 ) | ( n5178 & n5268 ) ;
  assign n5270 = ( n5257 & n5267 ) | ( n5257 & n5269 ) | ( n5267 & n5269 ) ;
  assign n5271 = n1398 & n2083 ;
  assign n5272 = x26 & n5271 ;
  assign n5273 = n1316 & n4200 ;
  assign n5274 = ~n1207 & n4215 ;
  assign n5275 = n5273 | n5274 ;
  assign n5276 = n4203 | n5275 ;
  assign n5277 = ( ~n4157 & n5275 ) | ( ~n4157 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5278 = x26 & ~n5277 ;
  assign n5279 = ( ~x26 & n5271 ) | ( ~x26 & n5277 ) | ( n5271 & n5277 ) ;
  assign n5280 = ( ~n5272 & n5278 ) | ( ~n5272 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = ( n5178 & n5188 ) | ( n5178 & n5190 ) | ( n5188 & n5190 ) ;
  assign n5282 = ( n5178 & n5191 ) | ( n5178 & ~n5281 ) | ( n5191 & ~n5281 ) ;
  assign n5283 = ( n5270 & n5280 ) | ( n5270 & ~n5282 ) | ( n5280 & ~n5282 ) ;
  assign n5284 = n859 & n4637 ;
  assign n5285 = ~n721 & n4649 ;
  assign n5286 = n5284 | n5285 ;
  assign n5287 = n995 & n4584 ;
  assign n5288 = n5286 | n5287 ;
  assign n5289 = n4591 | n5288 ;
  assign n5290 = ( ~n3829 & n5288 ) | ( ~n3829 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5291 = x23 & ~n5290 ;
  assign n5292 = ~x23 & n5290 ;
  assign n5293 = n5291 | n5292 ;
  assign n5294 = ( n5247 & n5283 ) | ( n5247 & n5293 ) | ( n5283 & n5293 ) ;
  assign n5295 = ~n3601 & n5232 ;
  assign n5296 = ~n3533 & n4878 ;
  assign n5297 = n5295 | n5296 ;
  assign n5298 = ~n3487 & n4874 ;
  assign n5299 = n5297 | n5298 ;
  assign n5300 = n4879 | n5299 ;
  assign n5301 = ( ~n4223 & n5299 ) | ( ~n4223 & n5300 ) | ( n5299 & n5300 ) ;
  assign n5302 = x20 & ~n5301 ;
  assign n5303 = ~x20 & n5301 ;
  assign n5304 = n5302 | n5303 ;
  assign n5305 = ( ~n5204 & n5214 ) | ( ~n5204 & n5216 ) | ( n5214 & n5216 ) ;
  assign n5306 = ( ~n5214 & n5217 ) | ( ~n5214 & n5305 ) | ( n5217 & n5305 ) ;
  assign n5307 = ( n5294 & n5304 ) | ( n5294 & ~n5306 ) | ( n5304 & ~n5306 ) ;
  assign n5308 = ~n3533 & n5232 ;
  assign n5309 = x20 & n5308 ;
  assign n5310 = ~n3516 & n4878 ;
  assign n5311 = n4874 | n5310 ;
  assign n5312 = ( ~n3601 & n5310 ) | ( ~n3601 & n5311 ) | ( n5310 & n5311 ) ;
  assign n5313 = n4879 | n5312 ;
  assign n5314 = ( ~n4058 & n5312 ) | ( ~n4058 & n5313 ) | ( n5312 & n5313 ) ;
  assign n5315 = x20 & ~n5314 ;
  assign n5316 = ( ~x20 & n5308 ) | ( ~x20 & n5314 ) | ( n5308 & n5314 ) ;
  assign n5317 = ( ~n5309 & n5315 ) | ( ~n5309 & n5316 ) | ( n5315 & n5316 ) ;
  assign n5318 = ( n5245 & n5307 ) | ( n5245 & n5317 ) | ( n5307 & n5317 ) ;
  assign n5319 = ~n2041 & n3536 ;
  assign n5320 = n1943 & n3501 ;
  assign n5321 = n5319 | n5320 ;
  assign n5322 = ~n1841 & n4039 ;
  assign n5323 = n5321 | n5322 ;
  assign n5324 = x29 & n5323 ;
  assign n5325 = n3541 & ~n4753 ;
  assign n5326 = x29 & ~n5325 ;
  assign n5327 = ( ~x29 & n5323 ) | ( ~x29 & n5325 ) | ( n5323 & n5325 ) ;
  assign n5328 = ( ~n5324 & n5326 ) | ( ~n5324 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5329 = n2102 & n3248 ;
  assign n5330 = ( ~n2102 & n3137 ) | ( ~n2102 & n3248 ) | ( n3137 & n3248 ) ;
  assign n5331 = ( n3138 & ~n5329 ) | ( n3138 & n5330 ) | ( ~n5329 & n5330 ) ;
  assign n5332 = n2102 & n3270 ;
  assign n5333 = n2187 & n3274 ;
  assign n5334 = n5332 | n5333 ;
  assign n5335 = ~n2282 & n3273 ;
  assign n5336 = n5334 | n5335 ;
  assign n5337 = n390 | n5336 ;
  assign n5338 = ( ~n5331 & n5336 ) | ( ~n5331 & n5337 ) | ( n5336 & n5337 ) ;
  assign n5339 = ( n4934 & ~n5139 ) | ( n4934 & n5160 ) | ( ~n5139 & n5160 ) ;
  assign n5340 = ( ~n4934 & n5161 ) | ( ~n4934 & n5339 ) | ( n5161 & n5339 ) ;
  assign n5341 = ( n5328 & n5338 ) | ( n5328 & n5340 ) | ( n5338 & n5340 ) ;
  assign n5342 = n1943 & n3536 ;
  assign n5343 = x29 & n5342 ;
  assign n5344 = n1792 & n4039 ;
  assign n5345 = ~n1841 & n3501 ;
  assign n5346 = n5344 | n5345 ;
  assign n5347 = n3541 | n5346 ;
  assign n5348 = ( ~n4831 & n5346 ) | ( ~n4831 & n5347 ) | ( n5346 & n5347 ) ;
  assign n5349 = x29 & ~n5348 ;
  assign n5350 = ( ~x29 & n5342 ) | ( ~x29 & n5348 ) | ( n5342 & n5348 ) ;
  assign n5351 = ( ~n5343 & n5349 ) | ( ~n5343 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5352 = ( n5004 & n5006 ) | ( n5004 & n5161 ) | ( n5006 & n5161 ) ;
  assign n5353 = ( n5004 & n5162 ) | ( n5004 & ~n5352 ) | ( n5162 & ~n5352 ) ;
  assign n5354 = ( n5341 & n5351 ) | ( n5341 & n5353 ) | ( n5351 & n5353 ) ;
  assign n5355 = ~n1529 & n4200 ;
  assign n5356 = n1600 & n2083 ;
  assign n5357 = n1398 & n4215 ;
  assign n5358 = n5356 | n5357 ;
  assign n5359 = n5355 | n5358 ;
  assign n5360 = x26 & n5359 ;
  assign n5361 = n4203 & ~n4324 ;
  assign n5362 = ( ~x26 & n5359 ) | ( ~x26 & n5361 ) | ( n5359 & n5361 ) ;
  assign n5363 = x26 & ~n5361 ;
  assign n5364 = ( ~n5360 & n5362 ) | ( ~n5360 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5365 = ( n5162 & n5172 ) | ( n5162 & n5174 ) | ( n5172 & n5174 ) ;
  assign n5366 = ( n5172 & n5175 ) | ( n5172 & ~n5365 ) | ( n5175 & ~n5365 ) ;
  assign n5367 = ( n5354 & n5364 ) | ( n5354 & n5366 ) | ( n5364 & n5366 ) ;
  assign n5368 = n995 & n4649 ;
  assign n5369 = ~n1207 & n4584 ;
  assign n5370 = n5368 | n5369 ;
  assign n5371 = ~n1118 & n4637 ;
  assign n5372 = n5370 | n5371 ;
  assign n5373 = n4591 | n5372 ;
  assign n5374 = ( n4173 & n5372 ) | ( n4173 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5375 = x23 & ~n5374 ;
  assign n5376 = ~x23 & n5374 ;
  assign n5377 = n5375 | n5376 ;
  assign n5378 = ( ~n5257 & n5267 ) | ( ~n5257 & n5269 ) | ( n5267 & n5269 ) ;
  assign n5379 = ( n5257 & ~n5270 ) | ( n5257 & n5378 ) | ( ~n5270 & n5378 ) ;
  assign n5380 = ( n5367 & n5377 ) | ( n5367 & n5379 ) | ( n5377 & n5379 ) ;
  assign n5381 = n859 & n4649 ;
  assign n5382 = n995 & n4637 ;
  assign n5383 = n5381 | n5382 ;
  assign n5384 = ~n1118 & n4584 ;
  assign n5385 = n5383 | n5384 ;
  assign n5386 = n4591 | n5385 ;
  assign n5387 = ( ~n4034 & n5385 ) | ( ~n4034 & n5386 ) | ( n5385 & n5386 ) ;
  assign n5388 = x23 & ~n5387 ;
  assign n5389 = ~x23 & n5387 ;
  assign n5390 = n5388 | n5389 ;
  assign n5391 = ( n5270 & ~n5280 ) | ( n5270 & n5282 ) | ( ~n5280 & n5282 ) ;
  assign n5392 = ( ~n5270 & n5283 ) | ( ~n5270 & n5391 ) | ( n5283 & n5391 ) ;
  assign n5393 = ( n5380 & n5390 ) | ( n5380 & ~n5392 ) | ( n5390 & ~n5392 ) ;
  assign n5394 = ( ~n5247 & n5283 ) | ( ~n5247 & n5293 ) | ( n5283 & n5293 ) ;
  assign n5395 = ( n5247 & ~n5294 ) | ( n5247 & n5394 ) | ( ~n5294 & n5394 ) ;
  assign n5396 = ~n3487 & n5232 ;
  assign n5397 = ~n3601 & n4878 ;
  assign n5398 = n564 & n4874 ;
  assign n5399 = n5397 | n5398 ;
  assign n5400 = n5396 | n5399 ;
  assign n5401 = n4879 | n5400 ;
  assign n5402 = ( n3674 & n5400 ) | ( n3674 & n5401 ) | ( n5400 & n5401 ) ;
  assign n5403 = x20 & ~n5402 ;
  assign n5404 = ~x20 & n5402 ;
  assign n5405 = n5403 | n5404 ;
  assign n5406 = ( n5393 & n5395 ) | ( n5393 & n5405 ) | ( n5395 & n5405 ) ;
  assign n5407 = x14 | x15 ;
  assign n5408 = x16 | n5407 ;
  assign n5409 = x17 & ~n5408 ;
  assign n5410 = x14 & x15 ;
  assign n5411 = x16 & n5410 ;
  assign n5412 = ~x17 & n5411 ;
  assign n5413 = n5409 | n5412 ;
  assign n5414 = n5407 & ~n5410 ;
  assign n5415 = x16 & x17 ;
  assign n5416 = x16 | x17 ;
  assign n5417 = ( n5414 & n5415 ) | ( n5414 & ~n5416 ) | ( n5415 & ~n5416 ) ;
  assign n5418 = n5414 & ~n5417 ;
  assign n5419 = ( ~n3516 & n3608 ) | ( ~n3516 & n5418 ) | ( n3608 & n5418 ) ;
  assign n5420 = ( ~n3607 & n5413 ) | ( ~n3607 & n5419 ) | ( n5413 & n5419 ) ;
  assign n5421 = x17 & ~n5420 ;
  assign n5422 = ~x17 & n5420 ;
  assign n5423 = n5421 | n5422 ;
  assign n5424 = ( ~n5294 & n5304 ) | ( ~n5294 & n5306 ) | ( n5304 & n5306 ) ;
  assign n5425 = ( ~n5304 & n5307 ) | ( ~n5304 & n5424 ) | ( n5307 & n5424 ) ;
  assign n5426 = ( n5406 & n5423 ) | ( n5406 & ~n5425 ) | ( n5423 & ~n5425 ) ;
  assign n5427 = n225 | n456 ;
  assign n5428 = n3312 | n5427 ;
  assign n5429 = n428 | n589 ;
  assign n5430 = n678 | n5429 ;
  assign n5431 = n5428 | n5430 ;
  assign n5432 = n917 | n1302 ;
  assign n5433 = n1111 | n5432 ;
  assign n5434 = n1338 | n5433 ;
  assign n5435 = n5431 | n5434 ;
  assign n5436 = n899 | n1010 ;
  assign n5437 = n5435 | n5436 ;
  assign n5438 = n497 | n554 ;
  assign n5439 = n1081 | n5438 ;
  assign n5440 = n923 | n2081 ;
  assign n5441 = n5439 | n5440 ;
  assign n5442 = n669 | n780 ;
  assign n5443 = n5441 | n5442 ;
  assign n5444 = n5437 | n5443 ;
  assign n5445 = n4438 | n5444 ;
  assign n5446 = n170 | n1078 ;
  assign n5447 = n5445 | n5446 ;
  assign n5448 = ( x2 & x5 ) | ( x2 & ~n5447 ) | ( x5 & ~n5447 ) ;
  assign n5449 = ~n3133 & n3244 ;
  assign n5450 = n2398 | n5449 ;
  assign n5451 = n3134 & n3244 ;
  assign n5452 = n5450 & ~n5451 ;
  assign n5453 = ~n2467 & n3274 ;
  assign n5454 = n2398 & n3270 ;
  assign n5455 = ~n2521 & n3273 ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = n5453 | n5456 ;
  assign n5458 = n390 | n5457 ;
  assign n5459 = ( n5452 & n5457 ) | ( n5452 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5460 = ( n5070 & ~n5448 ) | ( n5070 & n5459 ) | ( ~n5448 & n5459 ) ;
  assign n5461 = n221 | n942 ;
  assign n5462 = n359 | n5461 ;
  assign n5463 = n1151 | n5462 ;
  assign n5464 = n752 | n5463 ;
  assign n5465 = n161 | n614 ;
  assign n5466 = n140 | n5465 ;
  assign n5467 = n4507 | n5466 ;
  assign n5468 = n5464 | n5467 ;
  assign n5469 = n5105 | n5468 ;
  assign n5470 = n1357 | n2201 ;
  assign n5471 = n4755 | n5470 ;
  assign n5472 = n5041 | n5471 ;
  assign n5473 = n1432 | n5472 ;
  assign n5474 = n5469 | n5473 ;
  assign n5475 = n3950 | n5474 ;
  assign n5476 = n1110 | n1193 ;
  assign n5477 = n946 | n5476 ;
  assign n5478 = n775 | n5477 ;
  assign n5479 = n2019 | n2105 ;
  assign n5480 = n5478 | n5479 ;
  assign n5481 = n1971 | n3905 ;
  assign n5482 = n3724 | n5481 ;
  assign n5483 = n285 | n669 ;
  assign n5484 = n5117 | n5483 ;
  assign n5485 = n260 | n1074 ;
  assign n5486 = n1649 | n5485 ;
  assign n5487 = n5484 | n5486 ;
  assign n5488 = n5482 | n5487 ;
  assign n5489 = n5480 | n5488 ;
  assign n5490 = n5475 | n5489 ;
  assign n5491 = ( n5070 & n5460 ) | ( n5070 & n5490 ) | ( n5460 & n5490 ) ;
  assign n5492 = n2282 | n3246 ;
  assign n5493 = ( n2282 & n3135 ) | ( n2282 & ~n3246 ) | ( n3135 & ~n3246 ) ;
  assign n5494 = ( ~n3136 & n5492 ) | ( ~n3136 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5495 = ~n2364 & n3274 ;
  assign n5496 = ~n2282 & n3270 ;
  assign n5497 = n5495 | n5496 ;
  assign n5498 = n2398 & n3273 ;
  assign n5499 = n5497 | n5498 ;
  assign n5500 = n390 | n5499 ;
  assign n5501 = ( ~n5494 & n5499 ) | ( ~n5494 & n5500 ) | ( n5499 & n5500 ) ;
  assign n5502 = ( x8 & ~n5070 ) | ( x8 & n5127 ) | ( ~n5070 & n5127 ) ;
  assign n5503 = ( ~x8 & n5128 ) | ( ~x8 & n5502 ) | ( n5128 & n5502 ) ;
  assign n5504 = ( n5491 & n5501 ) | ( n5491 & n5503 ) | ( n5501 & n5503 ) ;
  assign n5505 = n2102 & n3536 ;
  assign n5506 = n1943 & n4039 ;
  assign n5507 = n5505 | n5506 ;
  assign n5508 = ~n2041 & n3501 ;
  assign n5509 = n5507 | n5508 ;
  assign n5510 = x29 & n5509 ;
  assign n5511 = n3541 & ~n4985 ;
  assign n5512 = x29 & ~n5511 ;
  assign n5513 = ( ~x29 & n5509 ) | ( ~x29 & n5511 ) | ( n5509 & n5511 ) ;
  assign n5514 = ( ~n5510 & n5512 ) | ( ~n5510 & n5513 ) | ( n5512 & n5513 ) ;
  assign n5515 = ( n4934 & ~n5128 ) | ( n4934 & n5138 ) | ( ~n5128 & n5138 ) ;
  assign n5516 = ( ~n4934 & n5139 ) | ( ~n4934 & n5515 ) | ( n5139 & n5515 ) ;
  assign n5517 = ( n5504 & n5514 ) | ( n5504 & n5516 ) | ( n5514 & n5516 ) ;
  assign n5518 = ( ~n5328 & n5338 ) | ( ~n5328 & n5340 ) | ( n5338 & n5340 ) ;
  assign n5519 = ( n5328 & ~n5341 ) | ( n5328 & n5518 ) | ( ~n5341 & n5518 ) ;
  assign n5520 = n1687 & n4200 ;
  assign n5521 = n1792 & n2083 ;
  assign n5522 = n1600 & n4215 ;
  assign n5523 = n5521 | n5522 ;
  assign n5524 = n5520 | n5523 ;
  assign n5525 = x26 & n5524 ;
  assign n5526 = n4203 & n4674 ;
  assign n5527 = x26 & ~n5526 ;
  assign n5528 = ( ~x26 & n5524 ) | ( ~x26 & n5526 ) | ( n5524 & n5526 ) ;
  assign n5529 = ( ~n5525 & n5527 ) | ( ~n5525 & n5528 ) | ( n5527 & n5528 ) ;
  assign n5530 = ( n5517 & n5519 ) | ( n5517 & n5529 ) | ( n5519 & n5529 ) ;
  assign n5531 = ~n1529 & n4215 ;
  assign n5532 = n1687 & n2083 ;
  assign n5533 = n5531 | n5532 ;
  assign n5534 = n1600 & n4200 ;
  assign n5535 = n5533 | n5534 ;
  assign n5536 = x26 & n5535 ;
  assign n5537 = n4203 & ~n4531 ;
  assign n5538 = x26 & ~n5537 ;
  assign n5539 = ( ~x26 & n5535 ) | ( ~x26 & n5537 ) | ( n5535 & n5537 ) ;
  assign n5540 = ( ~n5536 & n5538 ) | ( ~n5536 & n5539 ) | ( n5538 & n5539 ) ;
  assign n5541 = ( n5341 & ~n5351 ) | ( n5341 & n5353 ) | ( ~n5351 & n5353 ) ;
  assign n5542 = ( n5351 & ~n5354 ) | ( n5351 & n5541 ) | ( ~n5354 & n5541 ) ;
  assign n5543 = ( n5530 & n5540 ) | ( n5530 & n5542 ) | ( n5540 & n5542 ) ;
  assign n5544 = n1316 & n4584 ;
  assign n5545 = ~n1207 & n4637 ;
  assign n5546 = n5544 | n5545 ;
  assign n5547 = ~n1118 & n4649 ;
  assign n5548 = n5546 | n5547 ;
  assign n5549 = n4591 | n5548 ;
  assign n5550 = ( n3841 & n5548 ) | ( n3841 & n5549 ) | ( n5548 & n5549 ) ;
  assign n5551 = x23 & ~n5550 ;
  assign n5552 = ~x23 & n5550 ;
  assign n5553 = n5551 | n5552 ;
  assign n5554 = ( ~n5354 & n5364 ) | ( ~n5354 & n5366 ) | ( n5364 & n5366 ) ;
  assign n5555 = ( n5354 & ~n5367 ) | ( n5354 & n5554 ) | ( ~n5367 & n5554 ) ;
  assign n5556 = ( n5543 & n5553 ) | ( n5543 & n5555 ) | ( n5553 & n5555 ) ;
  assign n5557 = n859 & n4874 ;
  assign n5558 = ~n721 & n5232 ;
  assign n5559 = n5557 | n5558 ;
  assign n5560 = n564 & n4878 ;
  assign n5561 = n5559 | n5560 ;
  assign n5562 = n4879 | n5561 ;
  assign n5563 = ( ~n3268 & n5561 ) | ( ~n3268 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = x20 & ~n5563 ;
  assign n5565 = ~x20 & n5563 ;
  assign n5566 = n5564 | n5565 ;
  assign n5567 = ( ~n5367 & n5377 ) | ( ~n5367 & n5379 ) | ( n5377 & n5379 ) ;
  assign n5568 = ( n5367 & ~n5380 ) | ( n5367 & n5567 ) | ( ~n5380 & n5567 ) ;
  assign n5569 = ( n5556 & n5566 ) | ( n5556 & n5568 ) | ( n5566 & n5568 ) ;
  assign n5570 = ~n3487 & n4878 ;
  assign n5571 = ~n721 & n4874 ;
  assign n5572 = n564 & n5232 ;
  assign n5573 = n5571 | n5572 ;
  assign n5574 = n5570 | n5573 ;
  assign n5575 = n4879 | n5574 ;
  assign n5576 = ( ~n3492 & n5574 ) | ( ~n3492 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5577 = x20 & ~n5576 ;
  assign n5578 = ~x20 & n5576 ;
  assign n5579 = n5577 | n5578 ;
  assign n5580 = ( n5380 & ~n5390 ) | ( n5380 & n5392 ) | ( ~n5390 & n5392 ) ;
  assign n5581 = ( ~n5380 & n5393 ) | ( ~n5380 & n5580 ) | ( n5393 & n5580 ) ;
  assign n5582 = ( n5569 & n5579 ) | ( n5569 & ~n5581 ) | ( n5579 & ~n5581 ) ;
  assign n5583 = n5411 | n5414 ;
  assign n5584 = n5408 & ~n5583 ;
  assign n5585 = ~n3516 & n5584 ;
  assign n5586 = x17 & n5585 ;
  assign n5587 = ~n3533 & n5413 ;
  assign n5588 = n5418 | n5587 ;
  assign n5589 = ( n3609 & n5587 ) | ( n3609 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = x17 & ~n5589 ;
  assign n5591 = ( ~x17 & n5585 ) | ( ~x17 & n5589 ) | ( n5585 & n5589 ) ;
  assign n5592 = ( ~n5586 & n5590 ) | ( ~n5586 & n5591 ) | ( n5590 & n5591 ) ;
  assign n5593 = ( ~n5393 & n5395 ) | ( ~n5393 & n5405 ) | ( n5395 & n5405 ) ;
  assign n5594 = ( n5393 & ~n5406 ) | ( n5393 & n5593 ) | ( ~n5406 & n5593 ) ;
  assign n5595 = ( n5582 & n5592 ) | ( n5582 & n5594 ) | ( n5592 & n5594 ) ;
  assign n5596 = n2642 & n3240 ;
  assign n5597 = ( n2642 & n3129 ) | ( n2642 & ~n3240 ) | ( n3129 & ~n3240 ) ;
  assign n5598 = ( ~n3130 & n5596 ) | ( ~n3130 & n5597 ) | ( n5596 & n5597 ) ;
  assign n5599 = n2735 & n3274 ;
  assign n5600 = n2642 & n3270 ;
  assign n5601 = n5599 | n5600 ;
  assign n5602 = n2820 & n3273 ;
  assign n5603 = n5601 | n5602 ;
  assign n5604 = n390 | n5603 ;
  assign n5605 = ( n5598 & n5603 ) | ( n5598 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5606 = n269 | n616 ;
  assign n5607 = n178 | n542 ;
  assign n5608 = n5606 | n5607 ;
  assign n5609 = n5150 | n5608 ;
  assign n5610 = n3356 | n5609 ;
  assign n5611 = n342 | n485 ;
  assign n5612 = n533 | n550 ;
  assign n5613 = n5611 | n5612 ;
  assign n5614 = n257 | n1069 ;
  assign n5615 = n5613 | n5614 ;
  assign n5616 = n5610 | n5615 ;
  assign n5617 = n298 | n321 ;
  assign n5618 = n758 | n3167 ;
  assign n5619 = n5617 | n5618 ;
  assign n5620 = n3394 | n5619 ;
  assign n5621 = n5616 | n5620 ;
  assign n5622 = n3212 | n5621 ;
  assign n5623 = n1883 | n5622 ;
  assign n5624 = n928 | n1691 ;
  assign n5625 = n1660 | n5624 ;
  assign n5626 = n5155 | n5625 ;
  assign n5627 = n2918 | n4006 ;
  assign n5628 = n82 | n2440 ;
  assign n5629 = n5627 | n5628 ;
  assign n5630 = n1275 | n5629 ;
  assign n5631 = n5626 | n5630 ;
  assign n5632 = n1955 | n5066 ;
  assign n5633 = n5631 | n5632 ;
  assign n5634 = n5623 | n5633 ;
  assign n5635 = n3686 | n3852 ;
  assign n5636 = n210 | n278 ;
  assign n5637 = n2024 | n5636 ;
  assign n5638 = n269 | n835 ;
  assign n5639 = n5637 | n5638 ;
  assign n5640 = n5635 | n5639 ;
  assign n5641 = n4399 | n5640 ;
  assign n5642 = n355 | n5641 ;
  assign n5643 = n1012 | n1518 ;
  assign n5644 = n96 | n185 ;
  assign n5645 = n678 | n5644 ;
  assign n5646 = n5643 | n5645 ;
  assign n5647 = n757 | n4782 ;
  assign n5648 = n5646 | n5647 ;
  assign n5649 = n1105 | n5648 ;
  assign n5650 = n5642 | n5649 ;
  assign n5651 = n1205 | n5650 ;
  assign n5652 = n3122 | n5651 ;
  assign n5653 = n5634 | n5652 ;
  assign n5654 = x2 & n5653 ;
  assign n5655 = ( x2 & n5605 ) | ( x2 & n5654 ) | ( n5605 & n5654 ) ;
  assign n5656 = x2 | n5652 ;
  assign n5657 = ( x2 & n5634 ) | ( x2 & n5656 ) | ( n5634 & n5656 ) ;
  assign n5658 = ( x2 & n5605 ) | ( x2 & n5657 ) | ( n5605 & n5657 ) ;
  assign n5659 = n614 | n3761 ;
  assign n5660 = n2576 | n5659 ;
  assign n5661 = n48 | n667 ;
  assign n5662 = n5660 | n5661 ;
  assign n5663 = n1768 | n5662 ;
  assign n5664 = n298 | n1392 ;
  assign n5665 = n4348 | n5664 ;
  assign n5666 = n4964 | n5665 ;
  assign n5667 = n5663 | n5666 ;
  assign n5668 = n3971 | n5667 ;
  assign n5669 = n89 | n392 ;
  assign n5670 = n987 | n5669 ;
  assign n5671 = n308 | n329 ;
  assign n5672 = n5670 | n5671 ;
  assign n5673 = n765 | n5672 ;
  assign n5674 = n2995 | n5673 ;
  assign n5675 = n351 | n928 ;
  assign n5676 = n225 | n5157 ;
  assign n5677 = n5675 | n5676 ;
  assign n5678 = n5674 | n5677 ;
  assign n5679 = n813 | n5678 ;
  assign n5680 = n5668 | n5679 ;
  assign n5681 = n2543 | n5680 ;
  assign n5682 = n2847 & ~n5681 ;
  assign n5683 = n5658 & ~n5682 ;
  assign n5684 = n5655 | n5683 ;
  assign n5685 = ~n2467 & n3270 ;
  assign n5686 = ~n2521 & n3274 ;
  assign n5687 = ~n2608 & n3273 ;
  assign n5688 = n5686 | n5687 ;
  assign n5689 = n5685 | n5688 ;
  assign n5690 = n390 | n5689 ;
  assign n5691 = n3133 & ~n3243 ;
  assign n5692 = n3132 & ~n3244 ;
  assign n5693 = ( n2467 & ~n5691 ) | ( n2467 & n5692 ) | ( ~n5691 & n5692 ) ;
  assign n5694 = ( n5689 & n5690 ) | ( n5689 & ~n5693 ) | ( n5690 & ~n5693 ) ;
  assign n5695 = ( x2 & ~x5 ) | ( x2 & n5447 ) | ( ~x5 & n5447 ) ;
  assign n5696 = ( ~x2 & n5448 ) | ( ~x2 & n5695 ) | ( n5448 & n5695 ) ;
  assign n5697 = ( n5684 & n5694 ) | ( n5684 & n5696 ) | ( n5694 & n5696 ) ;
  assign n5698 = ~n2364 & n3536 ;
  assign n5699 = n2187 & n4039 ;
  assign n5700 = n5698 | n5699 ;
  assign n5701 = ~n2282 & n3501 ;
  assign n5702 = n5700 | n5701 ;
  assign n5703 = x29 & n5702 ;
  assign n5704 = n3541 & n5137 ;
  assign n5705 = x29 & ~n5704 ;
  assign n5706 = ( ~x29 & n5702 ) | ( ~x29 & n5704 ) | ( n5702 & n5704 ) ;
  assign n5707 = ( ~n5703 & n5705 ) | ( ~n5703 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = ( n5070 & n5448 ) | ( n5070 & ~n5459 ) | ( n5448 & ~n5459 ) ;
  assign n5709 = ( ~n5070 & n5460 ) | ( ~n5070 & n5708 ) | ( n5460 & n5708 ) ;
  assign n5710 = ( n5697 & n5707 ) | ( n5697 & ~n5709 ) | ( n5707 & ~n5709 ) ;
  assign n5711 = ( n2364 & ~n3133 ) | ( n2364 & n5450 ) | ( ~n3133 & n5450 ) ;
  assign n5712 = ( n2364 & n3133 ) | ( n2364 & ~n5450 ) | ( n3133 & ~n5450 ) ;
  assign n5713 = ( ~n2364 & n5711 ) | ( ~n2364 & n5712 ) | ( n5711 & n5712 ) ;
  assign n5714 = ~n2467 & n3273 ;
  assign n5715 = ~n2364 & n3270 ;
  assign n5716 = n5714 | n5715 ;
  assign n5717 = n2398 & n3274 ;
  assign n5718 = n5716 | n5717 ;
  assign n5719 = n390 | n5718 ;
  assign n5720 = ( n5713 & n5718 ) | ( n5713 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5721 = ( ~n5070 & n5460 ) | ( ~n5070 & n5490 ) | ( n5460 & n5490 ) ;
  assign n5722 = ( n5070 & ~n5491 ) | ( n5070 & n5721 ) | ( ~n5491 & n5721 ) ;
  assign n5723 = ( n5710 & n5720 ) | ( n5710 & n5722 ) | ( n5720 & n5722 ) ;
  assign n5724 = n2102 & n3501 ;
  assign n5725 = ~n2041 & n4039 ;
  assign n5726 = n5724 | n5725 ;
  assign n5727 = n2187 & n3536 ;
  assign n5728 = n5726 | n5727 ;
  assign n5729 = n3541 | n5728 ;
  assign n5730 = ( ~n4997 & n5728 ) | ( ~n4997 & n5729 ) | ( n5728 & n5729 ) ;
  assign n5731 = x29 & ~n5730 ;
  assign n5732 = ~x29 & n5730 ;
  assign n5733 = n5731 | n5732 ;
  assign n5734 = ( ~n5491 & n5501 ) | ( ~n5491 & n5503 ) | ( n5501 & n5503 ) ;
  assign n5735 = ( n5491 & ~n5504 ) | ( n5491 & n5734 ) | ( ~n5504 & n5734 ) ;
  assign n5736 = ( n5723 & n5733 ) | ( n5723 & n5735 ) | ( n5733 & n5735 ) ;
  assign n5737 = n1687 & n4215 ;
  assign n5738 = n1792 & n4200 ;
  assign n5739 = n5737 | n5738 ;
  assign n5740 = ~n1841 & n2083 ;
  assign n5741 = n5739 | n5740 ;
  assign n5742 = x26 & n5741 ;
  assign n5743 = n4203 & n4331 ;
  assign n5744 = ( ~x26 & n5741 ) | ( ~x26 & n5743 ) | ( n5741 & n5743 ) ;
  assign n5745 = x26 & ~n5743 ;
  assign n5746 = ( ~n5742 & n5744 ) | ( ~n5742 & n5745 ) | ( n5744 & n5745 ) ;
  assign n5747 = ( ~n5504 & n5514 ) | ( ~n5504 & n5516 ) | ( n5514 & n5516 ) ;
  assign n5748 = ( n5504 & ~n5517 ) | ( n5504 & n5747 ) | ( ~n5517 & n5747 ) ;
  assign n5749 = ( n5736 & n5746 ) | ( n5736 & n5748 ) | ( n5746 & n5748 ) ;
  assign n5750 = ~n1529 & n4584 ;
  assign n5751 = n1316 & n4649 ;
  assign n5752 = n5750 | n5751 ;
  assign n5753 = n1398 & n4637 ;
  assign n5754 = n5752 | n5753 ;
  assign n5755 = n4591 | n5754 ;
  assign n5756 = ( n4084 & n5754 ) | ( n4084 & n5755 ) | ( n5754 & n5755 ) ;
  assign n5757 = x23 & ~n5756 ;
  assign n5758 = ~x23 & n5756 ;
  assign n5759 = n5757 | n5758 ;
  assign n5760 = ( n5517 & ~n5519 ) | ( n5517 & n5529 ) | ( ~n5519 & n5529 ) ;
  assign n5761 = ( n5519 & ~n5530 ) | ( n5519 & n5760 ) | ( ~n5530 & n5760 ) ;
  assign n5762 = ( n5749 & n5759 ) | ( n5749 & n5761 ) | ( n5759 & n5761 ) ;
  assign n5763 = ( ~n5530 & n5540 ) | ( ~n5530 & n5542 ) | ( n5540 & n5542 ) ;
  assign n5764 = ( n5530 & ~n5543 ) | ( n5530 & n5763 ) | ( ~n5543 & n5763 ) ;
  assign n5765 = n1316 & n4637 ;
  assign n5766 = ~n1207 & n4649 ;
  assign n5767 = n1398 & n4584 ;
  assign n5768 = n5766 | n5767 ;
  assign n5769 = n5765 | n5768 ;
  assign n5770 = n4591 | n5769 ;
  assign n5771 = ( ~n4157 & n5769 ) | ( ~n4157 & n5770 ) | ( n5769 & n5770 ) ;
  assign n5772 = x23 & ~n5771 ;
  assign n5773 = ~x23 & n5771 ;
  assign n5774 = n5772 | n5773 ;
  assign n5775 = ( n5762 & n5764 ) | ( n5762 & n5774 ) | ( n5764 & n5774 ) ;
  assign n5776 = n859 & n5232 ;
  assign n5777 = ~n721 & n4878 ;
  assign n5778 = n5776 | n5777 ;
  assign n5779 = n995 & n4874 ;
  assign n5780 = n5778 | n5779 ;
  assign n5781 = n4879 | n5780 ;
  assign n5782 = ( ~n3829 & n5780 ) | ( ~n3829 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5783 = x20 & ~n5782 ;
  assign n5784 = ~x20 & n5782 ;
  assign n5785 = n5783 | n5784 ;
  assign n5786 = ( ~n5543 & n5553 ) | ( ~n5543 & n5555 ) | ( n5553 & n5555 ) ;
  assign n5787 = ( n5543 & ~n5556 ) | ( n5543 & n5786 ) | ( ~n5556 & n5786 ) ;
  assign n5788 = ( n5775 & n5785 ) | ( n5775 & n5787 ) | ( n5785 & n5787 ) ;
  assign n5789 = ~n3487 & n5413 ;
  assign n5790 = ~n3601 & n5584 ;
  assign n5791 = n3533 & n5417 ;
  assign n5792 = ( n5417 & n5790 ) | ( n5417 & ~n5791 ) | ( n5790 & ~n5791 ) ;
  assign n5793 = n5789 | n5792 ;
  assign n5794 = n5418 | n5793 ;
  assign n5795 = ( ~n4223 & n5793 ) | ( ~n4223 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5796 = x17 & ~n5795 ;
  assign n5797 = ~x17 & n5795 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = ( n5556 & ~n5566 ) | ( n5556 & n5568 ) | ( ~n5566 & n5568 ) ;
  assign n5800 = ( n5566 & ~n5569 ) | ( n5566 & n5799 ) | ( ~n5569 & n5799 ) ;
  assign n5801 = ( n5788 & n5798 ) | ( n5788 & n5800 ) | ( n5798 & n5800 ) ;
  assign n5802 = ~n3533 & n5584 ;
  assign n5803 = x17 & n5802 ;
  assign n5804 = ~n3516 & n5417 ;
  assign n5805 = n5413 | n5804 ;
  assign n5806 = ( ~n3601 & n5804 ) | ( ~n3601 & n5805 ) | ( n5804 & n5805 ) ;
  assign n5807 = n5418 | n5806 ;
  assign n5808 = ( ~n4058 & n5806 ) | ( ~n4058 & n5807 ) | ( n5806 & n5807 ) ;
  assign n5809 = x17 & ~n5808 ;
  assign n5810 = ( ~x17 & n5802 ) | ( ~x17 & n5808 ) | ( n5802 & n5808 ) ;
  assign n5811 = ( ~n5803 & n5809 ) | ( ~n5803 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5812 = ( n5569 & ~n5579 ) | ( n5569 & n5581 ) | ( ~n5579 & n5581 ) ;
  assign n5813 = ( ~n5569 & n5582 ) | ( ~n5569 & n5812 ) | ( n5582 & n5812 ) ;
  assign n5814 = ( n5801 & n5811 ) | ( n5801 & ~n5813 ) | ( n5811 & ~n5813 ) ;
  assign n5815 = ( ~n5723 & n5733 ) | ( ~n5723 & n5735 ) | ( n5733 & n5735 ) ;
  assign n5816 = ( n5723 & ~n5736 ) | ( n5723 & n5815 ) | ( ~n5736 & n5815 ) ;
  assign n5817 = n1943 & n2083 ;
  assign n5818 = n1792 & n4215 ;
  assign n5819 = n5817 | n5818 ;
  assign n5820 = ~n1841 & n4200 ;
  assign n5821 = n5819 | n5820 ;
  assign n5822 = x26 & n5821 ;
  assign n5823 = n4203 & ~n4831 ;
  assign n5824 = x26 & ~n5823 ;
  assign n5825 = ( ~x26 & n5821 ) | ( ~x26 & n5823 ) | ( n5821 & n5823 ) ;
  assign n5826 = ( ~n5822 & n5824 ) | ( ~n5822 & n5825 ) | ( n5824 & n5825 ) ;
  assign n5827 = ( ~n5710 & n5720 ) | ( ~n5710 & n5722 ) | ( n5720 & n5722 ) ;
  assign n5828 = ( n5710 & ~n5723 ) | ( n5710 & n5827 ) | ( ~n5723 & n5827 ) ;
  assign n5829 = ~n1841 & n4215 ;
  assign n5830 = ~n2041 & n2083 ;
  assign n5831 = n5829 | n5830 ;
  assign n5832 = n1943 & n4200 ;
  assign n5833 = n5831 | n5832 ;
  assign n5834 = n4203 | n5833 ;
  assign n5835 = ( ~n4753 & n5833 ) | ( ~n4753 & n5834 ) | ( n5833 & n5834 ) ;
  assign n5836 = x26 & ~n5835 ;
  assign n5837 = ~x26 & n5835 ;
  assign n5838 = n5836 | n5837 ;
  assign n5839 = n2102 & n4039 ;
  assign n5840 = n2187 & n3501 ;
  assign n5841 = n5839 | n5840 ;
  assign n5842 = ~n2282 & n3536 ;
  assign n5843 = n5841 | n5842 ;
  assign n5844 = n3541 | n5843 ;
  assign n5845 = ( ~n5331 & n5843 ) | ( ~n5331 & n5844 ) | ( n5843 & n5844 ) ;
  assign n5846 = x29 & ~n5845 ;
  assign n5847 = ~x29 & n5845 ;
  assign n5848 = n5846 | n5847 ;
  assign n5849 = ( n5828 & n5838 ) | ( n5828 & n5848 ) | ( n5838 & n5848 ) ;
  assign n5850 = ( n5816 & n5826 ) | ( n5816 & n5849 ) | ( n5826 & n5849 ) ;
  assign n5851 = ( ~n5736 & n5746 ) | ( ~n5736 & n5748 ) | ( n5746 & n5748 ) ;
  assign n5852 = ( n5736 & ~n5749 ) | ( n5736 & n5851 ) | ( ~n5749 & n5851 ) ;
  assign n5853 = n1600 & n4584 ;
  assign n5854 = x23 & n5853 ;
  assign n5855 = n1398 & n4649 ;
  assign n5856 = n4637 | n5855 ;
  assign n5857 = ( ~n1529 & n5855 ) | ( ~n1529 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5858 = n4591 | n5857 ;
  assign n5859 = ( ~n4324 & n5857 ) | ( ~n4324 & n5858 ) | ( n5857 & n5858 ) ;
  assign n5860 = x23 & ~n5859 ;
  assign n5861 = ( ~x23 & n5853 ) | ( ~x23 & n5859 ) | ( n5853 & n5859 ) ;
  assign n5862 = ( ~n5854 & n5860 ) | ( ~n5854 & n5861 ) | ( n5860 & n5861 ) ;
  assign n5863 = ( n5850 & n5852 ) | ( n5850 & n5862 ) | ( n5852 & n5862 ) ;
  assign n5864 = ( ~n5749 & n5759 ) | ( ~n5749 & n5761 ) | ( n5759 & n5761 ) ;
  assign n5865 = ( n5749 & ~n5762 ) | ( n5749 & n5864 ) | ( ~n5762 & n5864 ) ;
  assign n5866 = n995 & n4878 ;
  assign n5867 = ~n1207 & n4874 ;
  assign n5868 = n5866 | n5867 ;
  assign n5869 = ~n1118 & n5232 ;
  assign n5870 = n5868 | n5869 ;
  assign n5871 = n4879 | n5870 ;
  assign n5872 = ( n4173 & n5870 ) | ( n4173 & n5871 ) | ( n5870 & n5871 ) ;
  assign n5873 = x20 & ~n5872 ;
  assign n5874 = ~x20 & n5872 ;
  assign n5875 = n5873 | n5874 ;
  assign n5876 = ( n5863 & n5865 ) | ( n5863 & n5875 ) | ( n5865 & n5875 ) ;
  assign n5877 = ( ~n5762 & n5764 ) | ( ~n5762 & n5774 ) | ( n5764 & n5774 ) ;
  assign n5878 = ( n5762 & ~n5775 ) | ( n5762 & n5877 ) | ( ~n5775 & n5877 ) ;
  assign n5879 = n859 & n4878 ;
  assign n5880 = n995 & n5232 ;
  assign n5881 = n5879 | n5880 ;
  assign n5882 = ~n1118 & n4874 ;
  assign n5883 = n5881 | n5882 ;
  assign n5884 = n4879 | n5883 ;
  assign n5885 = ( ~n4034 & n5883 ) | ( ~n4034 & n5884 ) | ( n5883 & n5884 ) ;
  assign n5886 = x20 & ~n5885 ;
  assign n5887 = ~x20 & n5885 ;
  assign n5888 = n5886 | n5887 ;
  assign n5889 = ( n5876 & n5878 ) | ( n5876 & n5888 ) | ( n5878 & n5888 ) ;
  assign n5890 = ~n3487 & n5584 ;
  assign n5891 = ~n3601 & n5417 ;
  assign n5892 = ~n564 & n5413 ;
  assign n5893 = ( n5413 & n5891 ) | ( n5413 & ~n5892 ) | ( n5891 & ~n5892 ) ;
  assign n5894 = n5890 | n5893 ;
  assign n5895 = n5418 | n5894 ;
  assign n5896 = ( n3674 & n5894 ) | ( n3674 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5897 = x17 & ~n5896 ;
  assign n5898 = ~x17 & n5896 ;
  assign n5899 = n5897 | n5898 ;
  assign n5900 = ( ~n5775 & n5785 ) | ( ~n5775 & n5787 ) | ( n5785 & n5787 ) ;
  assign n5901 = ( n5775 & ~n5788 ) | ( n5775 & n5900 ) | ( ~n5788 & n5900 ) ;
  assign n5902 = ( n5889 & n5899 ) | ( n5889 & n5901 ) | ( n5899 & n5901 ) ;
  assign n5903 = x11 | x12 ;
  assign n5904 = x13 | n5903 ;
  assign n5905 = x14 & ~n5904 ;
  assign n5906 = x11 & x13 ;
  assign n5907 = x12 & ~x14 ;
  assign n5908 = n5906 & n5907 ;
  assign n5909 = n5905 | n5908 ;
  assign n5910 = x11 & ~x12 ;
  assign n5911 = ( ~x11 & n5903 ) | ( ~x11 & n5910 ) | ( n5903 & n5910 ) ;
  assign n5912 = x13 & x14 ;
  assign n5913 = x13 | x14 ;
  assign n5914 = ( n5911 & n5912 ) | ( n5911 & ~n5913 ) | ( n5912 & ~n5913 ) ;
  assign n5915 = n5911 & ~n5914 ;
  assign n5916 = ( ~n3516 & n3608 ) | ( ~n3516 & n5915 ) | ( n3608 & n5915 ) ;
  assign n5917 = ( ~n3607 & n5909 ) | ( ~n3607 & n5916 ) | ( n5909 & n5916 ) ;
  assign n5918 = x14 & ~n5917 ;
  assign n5919 = ~x14 & n5917 ;
  assign n5920 = n5918 | n5919 ;
  assign n5921 = ( ~n5788 & n5798 ) | ( ~n5788 & n5800 ) | ( n5798 & n5800 ) ;
  assign n5922 = ( n5788 & ~n5801 ) | ( n5788 & n5921 ) | ( ~n5801 & n5921 ) ;
  assign n5923 = ( n5902 & n5920 ) | ( n5902 & n5922 ) | ( n5920 & n5922 ) ;
  assign n5924 = n2944 | n3236 ;
  assign n5925 = ( n2944 & n3125 ) | ( n2944 & ~n3236 ) | ( n3125 & ~n3236 ) ;
  assign n5926 = ( ~n3126 & n5924 ) | ( ~n3126 & n5925 ) | ( n5924 & n5925 ) ;
  assign n5927 = ~n2944 & n3270 ;
  assign n5928 = ~n2977 & n3274 ;
  assign n5929 = n5927 | n5928 ;
  assign n5930 = n3123 & n3273 ;
  assign n5931 = n5929 | n5930 ;
  assign n5932 = n390 | n5931 ;
  assign n5933 = ( ~n5926 & n5931 ) | ( ~n5926 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5934 = n570 | n4397 ;
  assign n5935 = n4142 | n5934 ;
  assign n5936 = n557 | n586 ;
  assign n5937 = n5935 | n5936 ;
  assign n5938 = n281 | n617 ;
  assign n5939 = n163 | n455 ;
  assign n5940 = n63 | n5939 ;
  assign n5941 = n5938 | n5940 ;
  assign n5942 = n5937 | n5941 ;
  assign n5943 = n96 | n616 ;
  assign n5944 = n413 | n5943 ;
  assign n5945 = n3756 | n5944 ;
  assign n5946 = n2999 | n3934 ;
  assign n5947 = n5945 | n5946 ;
  assign n5948 = n191 | n1414 ;
  assign n5949 = n1906 | n3454 ;
  assign n5950 = n5948 | n5949 ;
  assign n5951 = n208 | n215 ;
  assign n5952 = n1720 | n5951 ;
  assign n5953 = n5950 | n5952 ;
  assign n5954 = n264 | n401 ;
  assign n5955 = n205 | n5954 ;
  assign n5956 = n3052 | n3229 ;
  assign n5957 = n5955 | n5956 ;
  assign n5958 = n758 | n2145 ;
  assign n5959 = n5957 | n5958 ;
  assign n5960 = n5953 | n5959 ;
  assign n5961 = n5947 | n5960 ;
  assign n5962 = n5942 | n5961 ;
  assign n5963 = n2722 | n5962 ;
  assign n5964 = n3123 & ~n3233 ;
  assign n5965 = n3234 | n5964 ;
  assign n5966 = n390 & n5965 ;
  assign n5967 = n3123 & n3270 ;
  assign n5968 = ~n3049 & n3274 ;
  assign n5969 = n5967 | n5968 ;
  assign n5970 = ~n3232 & n3273 ;
  assign n5971 = n5969 | n5970 ;
  assign n5972 = n5966 | n5971 ;
  assign n5973 = n3648 | n3714 ;
  assign n5974 = n614 | n678 ;
  assign n5975 = n5973 | n5974 ;
  assign n5976 = n164 | n780 ;
  assign n5977 = n809 | n5976 ;
  assign n5978 = n709 | n5977 ;
  assign n5979 = n5975 | n5978 ;
  assign n5980 = n1108 | n1131 ;
  assign n5981 = n5979 | n5980 ;
  assign n5982 = n200 | n1176 ;
  assign n5983 = n542 | n647 ;
  assign n5984 = n5982 | n5983 ;
  assign n5985 = n3000 | n5984 ;
  assign n5986 = n2940 | n5985 ;
  assign n5987 = n232 | n1041 ;
  assign n5988 = n657 | n5987 ;
  assign n5989 = n941 | n1294 ;
  assign n5990 = n5988 | n5989 ;
  assign n5991 = n5986 | n5990 ;
  assign n5992 = n5981 | n5991 ;
  assign n5993 = n2557 & ~n5992 ;
  assign n5994 = ~n3769 & n5993 ;
  assign n5995 = ~n4293 & n5994 ;
  assign n5996 = n5972 & ~n5995 ;
  assign n5997 = ~n2977 & n3235 ;
  assign n5998 = ( n2977 & n3124 ) | ( n2977 & n3235 ) | ( n3124 & n3235 ) ;
  assign n5999 = n2977 | n3124 ;
  assign n6000 = ( n5997 & ~n5998 ) | ( n5997 & n5999 ) | ( ~n5998 & n5999 ) ;
  assign n6001 = ~n2977 & n3270 ;
  assign n6002 = ~n3049 & n3273 ;
  assign n6003 = n6001 | n6002 ;
  assign n6004 = n3123 & n3274 ;
  assign n6005 = n6003 | n6004 ;
  assign n6006 = n390 | n6005 ;
  assign n6007 = ( n6000 & n6005 ) | ( n6000 & n6006 ) | ( n6005 & n6006 ) ;
  assign n6008 = n206 | n635 ;
  assign n6009 = n3622 | n6008 ;
  assign n6010 = n161 | n572 ;
  assign n6011 = n6009 | n6010 ;
  assign n6012 = n2173 | n6011 ;
  assign n6013 = n70 | n1542 ;
  assign n6014 = n331 | n6013 ;
  assign n6015 = n6012 | n6014 ;
  assign n6016 = n541 & n4202 ;
  assign n6017 = n124 | n589 ;
  assign n6018 = n6016 | n6017 ;
  assign n6019 = n892 | n6018 ;
  assign n6020 = n1824 | n4286 ;
  assign n6021 = n6019 | n6020 ;
  assign n6022 = n3638 | n6021 ;
  assign n6023 = n3085 | n6022 ;
  assign n6024 = n6015 | n6023 ;
  assign n6025 = n1974 | n6024 ;
  assign n6026 = n232 | n303 ;
  assign n6027 = n209 | n6026 ;
  assign n6028 = n3449 | n6027 ;
  assign n6029 = n1153 & ~n2162 ;
  assign n6030 = ~n6028 & n6029 ;
  assign n6031 = n1413 | n1537 ;
  assign n6032 = n2834 | n6031 ;
  assign n6033 = n321 | n545 ;
  assign n6034 = n774 | n6033 ;
  assign n6035 = n6032 | n6034 ;
  assign n6036 = n6030 & ~n6035 ;
  assign n6037 = n287 | n1086 ;
  assign n6038 = n550 | n6037 ;
  assign n6039 = n2263 | n6038 ;
  assign n6040 = n2787 | n3335 ;
  assign n6041 = n264 | n942 ;
  assign n6042 = n6040 | n6041 ;
  assign n6043 = n6039 | n6042 ;
  assign n6044 = n140 | n434 ;
  assign n6045 = n262 | n6044 ;
  assign n6046 = n2057 | n6045 ;
  assign n6047 = n6043 | n6046 ;
  assign n6048 = n6036 & ~n6047 ;
  assign n6049 = ~n6025 & n6048 ;
  assign n6050 = ( n5996 & n6007 ) | ( n5996 & ~n6049 ) | ( n6007 & ~n6049 ) ;
  assign n6051 = ( n5933 & n5963 ) | ( n5933 & n6050 ) | ( n5963 & n6050 ) ;
  assign n6052 = ~n2888 & n3237 ;
  assign n6053 = ( n2888 & ~n3126 ) | ( n2888 & n3237 ) | ( ~n3126 & n3237 ) ;
  assign n6054 = ~n2888 & n3126 ;
  assign n6055 = ( ~n6052 & n6053 ) | ( ~n6052 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6056 = ~n2888 & n3270 ;
  assign n6057 = ~n2977 & n3273 ;
  assign n6058 = ~n2944 & n3274 ;
  assign n6059 = n6057 | n6058 ;
  assign n6060 = n6056 | n6059 ;
  assign n6061 = n390 | n6060 ;
  assign n6062 = ( ~n6055 & n6060 ) | ( ~n6055 & n6061 ) | ( n6060 & n6061 ) ;
  assign n6063 = n192 | n435 ;
  assign n6064 = n968 | n6063 ;
  assign n6065 = n2805 | n6064 ;
  assign n6066 = n2756 | n6065 ;
  assign n6067 = n226 | n2081 ;
  assign n6068 = n74 | n1048 ;
  assign n6069 = n6067 | n6068 ;
  assign n6070 = n208 | n296 ;
  assign n6071 = n526 | n6070 ;
  assign n6072 = n3445 | n6071 ;
  assign n6073 = n6069 | n6072 ;
  assign n6074 = n511 | n6073 ;
  assign n6075 = n6066 | n6074 ;
  assign n6076 = n1199 | n2670 ;
  assign n6077 = n5974 | n6076 ;
  assign n6078 = n1572 | n6077 ;
  assign n6079 = n329 | n661 ;
  assign n6080 = n380 | n6079 ;
  assign n6081 = n91 | n6080 ;
  assign n6082 = n6078 | n6081 ;
  assign n6083 = n6075 | n6082 ;
  assign n6084 = n178 | n2971 ;
  assign n6085 = n2357 | n6084 ;
  assign n6086 = n3194 | n6085 ;
  assign n6087 = n5153 | n6086 ;
  assign n6088 = n284 | n328 ;
  assign n6089 = n688 | n6088 ;
  assign n6090 = n207 | n468 ;
  assign n6091 = n656 | n6090 ;
  assign n6092 = n6089 | n6091 ;
  assign n6093 = n110 | n125 ;
  assign n6094 = n1579 | n6093 ;
  assign n6095 = n6092 | n6094 ;
  assign n6096 = n2134 | n2789 ;
  assign n6097 = n6095 | n6096 ;
  assign n6098 = n1971 | n2373 ;
  assign n6099 = n6097 | n6098 ;
  assign n6100 = n6087 | n6099 ;
  assign n6101 = n6083 | n6100 ;
  assign n6102 = n5030 & ~n6101 ;
  assign n6103 = ( n6051 & n6062 ) | ( n6051 & ~n6102 ) | ( n6062 & ~n6102 ) ;
  assign n6104 = n2820 & ~n3238 ;
  assign n6105 = ( n2820 & ~n3127 ) | ( n2820 & n3238 ) | ( ~n3127 & n3238 ) ;
  assign n6106 = ( ~n3128 & n6104 ) | ( ~n3128 & n6105 ) | ( n6104 & n6105 ) ;
  assign n6107 = ~n2944 & n3273 ;
  assign n6108 = n2820 & n3270 ;
  assign n6109 = n6107 | n6108 ;
  assign n6110 = ~n2888 & n3274 ;
  assign n6111 = n6109 | n6110 ;
  assign n6112 = n390 | n6111 ;
  assign n6113 = ( n6106 & n6111 ) | ( n6106 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6114 = n1783 | n3450 ;
  assign n6115 = n941 | n3614 ;
  assign n6116 = n6114 | n6115 ;
  assign n6117 = n207 | n287 ;
  assign n6118 = n1094 | n6117 ;
  assign n6119 = n3037 | n6118 ;
  assign n6120 = n4917 | n6119 ;
  assign n6121 = n6116 | n6120 ;
  assign n6122 = n285 | n556 ;
  assign n6123 = n91 | n6122 ;
  assign n6124 = n225 | n6123 ;
  assign n6125 = n4282 | n6124 ;
  assign n6126 = n6121 | n6125 ;
  assign n6127 = n1142 | n6126 ;
  assign n6128 = n1365 | n2222 ;
  assign n6129 = n2663 | n6128 ;
  assign n6130 = n189 | n841 ;
  assign n6131 = n1737 | n6130 ;
  assign n6132 = n6129 | n6131 ;
  assign n6133 = n1253 | n1770 ;
  assign n6134 = n2550 | n6133 ;
  assign n6135 = n6132 | n6134 ;
  assign n6136 = n3355 | n4475 ;
  assign n6137 = n97 | n2211 ;
  assign n6138 = n6136 | n6137 ;
  assign n6139 = n113 | n641 ;
  assign n6140 = n896 | n1264 ;
  assign n6141 = n6139 | n6140 ;
  assign n6142 = n1593 | n2269 ;
  assign n6143 = n6141 | n6142 ;
  assign n6144 = n6138 | n6143 ;
  assign n6145 = n6135 | n6144 ;
  assign n6146 = n4966 | n6145 ;
  assign n6147 = n6127 | n6146 ;
  assign n6148 = ( n6103 & n6113 ) | ( n6103 & n6147 ) | ( n6113 & n6147 ) ;
  assign n6149 = ~n2888 & n3273 ;
  assign n6150 = n2735 & n3270 ;
  assign n6151 = n2820 & n3274 ;
  assign n6152 = n6150 | n6151 ;
  assign n6153 = n6149 | n6152 ;
  assign n6154 = n390 | n6153 ;
  assign n6155 = n3129 | n3239 ;
  assign n6156 = ~n3128 & n3240 ;
  assign n6157 = ( ~n2735 & n6155 ) | ( ~n2735 & n6156 ) | ( n6155 & n6156 ) ;
  assign n6158 = ( n6153 & n6154 ) | ( n6153 & ~n6157 ) | ( n6154 & ~n6157 ) ;
  assign n6159 = n734 | n3547 ;
  assign n6160 = n308 | n6159 ;
  assign n6161 = n146 | n6160 ;
  assign n6162 = n233 | n586 ;
  assign n6163 = n192 | n6162 ;
  assign n6164 = n2084 | n6163 ;
  assign n6165 = n6161 | n6164 ;
  assign n6166 = n2378 | n2946 ;
  assign n6167 = n923 | n2222 ;
  assign n6168 = n6166 | n6167 ;
  assign n6169 = n5643 | n6168 ;
  assign n6170 = n750 | n5034 ;
  assign n6171 = n1075 | n6170 ;
  assign n6172 = n6169 | n6171 ;
  assign n6173 = n6165 | n6172 ;
  assign n6174 = n4424 | n6173 ;
  assign n6175 = n4455 | n6174 ;
  assign n6176 = n835 | n1019 ;
  assign n6177 = n3100 | n6176 ;
  assign n6178 = n4470 | n6177 ;
  assign n6179 = n4411 | n6178 ;
  assign n6180 = n358 | n688 ;
  assign n6181 = n1560 | n1745 ;
  assign n6182 = n6180 | n6181 ;
  assign n6183 = n3059 | n4781 ;
  assign n6184 = n435 | n470 ;
  assign n6185 = n6183 | n6184 ;
  assign n6186 = n6182 | n6185 ;
  assign n6187 = n6179 | n6186 ;
  assign n6188 = n2329 | n6187 ;
  assign n6189 = n6175 | n6188 ;
  assign n6190 = ( n6148 & n6158 ) | ( n6148 & n6189 ) | ( n6158 & n6189 ) ;
  assign n6191 = ~n2467 & n4039 ;
  assign n6192 = x29 & n6191 ;
  assign n6193 = ~n2521 & n3501 ;
  assign n6194 = ~n2608 & n3536 ;
  assign n6195 = n6193 | n6194 ;
  assign n6196 = n3541 | n6195 ;
  assign n6197 = ( ~n5693 & n6195 ) | ( ~n5693 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6198 = x29 & ~n6197 ;
  assign n6199 = ( ~x29 & n6191 ) | ( ~x29 & n6197 ) | ( n6191 & n6197 ) ;
  assign n6200 = ( ~n6192 & n6198 ) | ( ~n6192 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = ( ~x2 & n5605 ) | ( ~x2 & n5634 ) | ( n5605 & n5634 ) ;
  assign n6202 = ( x2 & ~n5605 ) | ( x2 & n5634 ) | ( ~n5605 & n5634 ) ;
  assign n6203 = ( ~n5634 & n6201 ) | ( ~n5634 & n6202 ) | ( n6201 & n6202 ) ;
  assign n6204 = ( n6190 & n6200 ) | ( n6190 & n6203 ) | ( n6200 & n6203 ) ;
  assign n6205 = ( ~n5634 & n5652 ) | ( ~n5634 & n6202 ) | ( n5652 & n6202 ) ;
  assign n6206 = ( n5634 & n5652 ) | ( n5634 & n6202 ) | ( n5652 & n6202 ) ;
  assign n6207 = ( n5634 & n6205 ) | ( n5634 & ~n6206 ) | ( n6205 & ~n6206 ) ;
  assign n6208 = n2735 & n3273 ;
  assign n6209 = ~n2608 & n3270 ;
  assign n6210 = n2642 & n3274 ;
  assign n6211 = n6209 | n6210 ;
  assign n6212 = n6208 | n6211 ;
  assign n6213 = n390 | n6212 ;
  assign n6214 = n3131 & n3241 ;
  assign n6215 = ~n3130 & n3242 ;
  assign n6216 = ( n2608 & ~n6214 ) | ( n2608 & n6215 ) | ( ~n6214 & n6215 ) ;
  assign n6217 = ( n6212 & n6213 ) | ( n6212 & ~n6216 ) | ( n6213 & ~n6216 ) ;
  assign n6218 = ( n6204 & n6207 ) | ( n6204 & n6217 ) | ( n6207 & n6217 ) ;
  assign n6219 = ~n2521 & n3242 ;
  assign n6220 = ( n2521 & n3131 ) | ( n2521 & n3242 ) | ( n3131 & n3242 ) ;
  assign n6221 = ( n3132 & n6219 ) | ( n3132 & ~n6220 ) | ( n6219 & ~n6220 ) ;
  assign n6222 = ~n2608 & n3274 ;
  assign n6223 = ~n2521 & n3270 ;
  assign n6224 = n6222 | n6223 ;
  assign n6225 = n2642 & n3273 ;
  assign n6226 = n6224 | n6225 ;
  assign n6227 = n390 | n6226 ;
  assign n6228 = ( n6221 & n6226 ) | ( n6221 & n6227 ) | ( n6226 & n6227 ) ;
  assign n6229 = ( n5655 & n5658 ) | ( n5655 & n5682 ) | ( n5658 & n5682 ) ;
  assign n6230 = ( n5682 & n5684 ) | ( n5682 & ~n6229 ) | ( n5684 & ~n6229 ) ;
  assign n6231 = ( n6218 & n6228 ) | ( n6218 & ~n6230 ) | ( n6228 & ~n6230 ) ;
  assign n6232 = ~n2364 & n3501 ;
  assign n6233 = x29 & n6232 ;
  assign n6234 = ~n2282 & n4039 ;
  assign n6235 = n2398 & n3536 ;
  assign n6236 = n6234 | n6235 ;
  assign n6237 = n3541 | n6236 ;
  assign n6238 = ( ~n5494 & n6236 ) | ( ~n5494 & n6237 ) | ( n6236 & n6237 ) ;
  assign n6239 = x29 & ~n6238 ;
  assign n6240 = ( ~x29 & n6232 ) | ( ~x29 & n6238 ) | ( n6232 & n6238 ) ;
  assign n6241 = ( ~n6233 & n6239 ) | ( ~n6233 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6242 = ( ~n5684 & n5694 ) | ( ~n5684 & n5696 ) | ( n5694 & n5696 ) ;
  assign n6243 = ( n5684 & ~n5697 ) | ( n5684 & n6242 ) | ( ~n5697 & n6242 ) ;
  assign n6244 = ( n6231 & n6241 ) | ( n6231 & n6243 ) | ( n6241 & n6243 ) ;
  assign n6245 = ~n2041 & n4200 ;
  assign n6246 = x26 & n6245 ;
  assign n6247 = n1943 & n4215 ;
  assign n6248 = n2083 & n2102 ;
  assign n6249 = n6247 | n6248 ;
  assign n6250 = n4203 | n6249 ;
  assign n6251 = ( ~n4985 & n6249 ) | ( ~n4985 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6252 = x26 & ~n6251 ;
  assign n6253 = ( ~x26 & n6245 ) | ( ~x26 & n6251 ) | ( n6245 & n6251 ) ;
  assign n6254 = ( ~n6246 & n6252 ) | ( ~n6246 & n6253 ) | ( n6252 & n6253 ) ;
  assign n6255 = ( ~n5697 & n5707 ) | ( ~n5697 & n5709 ) | ( n5707 & n5709 ) ;
  assign n6256 = ( ~n5707 & n5710 ) | ( ~n5707 & n6255 ) | ( n5710 & n6255 ) ;
  assign n6257 = ( n6244 & n6254 ) | ( n6244 & ~n6256 ) | ( n6254 & ~n6256 ) ;
  assign n6258 = n1687 & n4637 ;
  assign n6259 = n1792 & n4584 ;
  assign n6260 = n1600 & n4649 ;
  assign n6261 = n6259 | n6260 ;
  assign n6262 = n6258 | n6261 ;
  assign n6263 = x23 & n6262 ;
  assign n6264 = n4591 & n4674 ;
  assign n6265 = x23 & ~n6264 ;
  assign n6266 = ( ~x23 & n6262 ) | ( ~x23 & n6264 ) | ( n6262 & n6264 ) ;
  assign n6267 = ( ~n6263 & n6265 ) | ( ~n6263 & n6266 ) | ( n6265 & n6266 ) ;
  assign n6268 = x26 & x29 ;
  assign n6269 = n3535 & ~n6268 ;
  assign n6270 = ~n5845 & n6269 ;
  assign n6271 = n5845 & ~n6269 ;
  assign n6272 = n6270 | n6271 ;
  assign n6273 = ( n5828 & n5835 ) | ( n5828 & n6272 ) | ( n5835 & n6272 ) ;
  assign n6274 = ( ~n5828 & n5835 ) | ( ~n5828 & n6272 ) | ( n5835 & n6272 ) ;
  assign n6275 = ( n5828 & ~n6273 ) | ( n5828 & n6274 ) | ( ~n6273 & n6274 ) ;
  assign n6276 = ( n6257 & n6267 ) | ( n6257 & n6275 ) | ( n6267 & n6275 ) ;
  assign n6277 = ( ~n5816 & n5826 ) | ( ~n5816 & n5849 ) | ( n5826 & n5849 ) ;
  assign n6278 = ( n5816 & ~n5850 ) | ( n5816 & n6277 ) | ( ~n5850 & n6277 ) ;
  assign n6279 = n1600 & n4637 ;
  assign n6280 = x23 & n6279 ;
  assign n6281 = ~n1529 & n4649 ;
  assign n6282 = n1687 & n4584 ;
  assign n6283 = n6281 | n6282 ;
  assign n6284 = n4591 | n6283 ;
  assign n6285 = ( ~n4531 & n6283 ) | ( ~n4531 & n6284 ) | ( n6283 & n6284 ) ;
  assign n6286 = x23 & ~n6285 ;
  assign n6287 = ( ~x23 & n6279 ) | ( ~x23 & n6285 ) | ( n6279 & n6285 ) ;
  assign n6288 = ( ~n6280 & n6286 ) | ( ~n6280 & n6287 ) | ( n6286 & n6287 ) ;
  assign n6289 = ( n6276 & n6278 ) | ( n6276 & n6288 ) | ( n6278 & n6288 ) ;
  assign n6290 = n1316 & n4874 ;
  assign n6291 = ~n1207 & n5232 ;
  assign n6292 = n6290 | n6291 ;
  assign n6293 = ~n1118 & n4878 ;
  assign n6294 = n6292 | n6293 ;
  assign n6295 = n4879 | n6294 ;
  assign n6296 = ( n3841 & n6294 ) | ( n3841 & n6295 ) | ( n6294 & n6295 ) ;
  assign n6297 = x20 & ~n6296 ;
  assign n6298 = ~x20 & n6296 ;
  assign n6299 = n6297 | n6298 ;
  assign n6300 = ( n5850 & ~n5852 ) | ( n5850 & n5862 ) | ( ~n5852 & n5862 ) ;
  assign n6301 = ( n5852 & ~n5863 ) | ( n5852 & n6300 ) | ( ~n5863 & n6300 ) ;
  assign n6302 = ( n6289 & n6299 ) | ( n6289 & n6301 ) | ( n6299 & n6301 ) ;
  assign n6303 = ~n721 & n5584 ;
  assign n6304 = x17 & n6303 ;
  assign n6305 = n859 & n5413 ;
  assign n6306 = n564 & n5417 ;
  assign n6307 = n6305 | n6306 ;
  assign n6308 = n5418 | n6307 ;
  assign n6309 = ( ~n3268 & n6307 ) | ( ~n3268 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = x17 & ~n6309 ;
  assign n6311 = ( ~x17 & n6303 ) | ( ~x17 & n6309 ) | ( n6303 & n6309 ) ;
  assign n6312 = ( ~n6304 & n6310 ) | ( ~n6304 & n6311 ) | ( n6310 & n6311 ) ;
  assign n6313 = ( ~n5863 & n5865 ) | ( ~n5863 & n5875 ) | ( n5865 & n5875 ) ;
  assign n6314 = ( n5863 & ~n5876 ) | ( n5863 & n6313 ) | ( ~n5876 & n6313 ) ;
  assign n6315 = ( n6302 & n6312 ) | ( n6302 & n6314 ) | ( n6312 & n6314 ) ;
  assign n6316 = ~n3487 & n5417 ;
  assign n6317 = ~n721 & n5413 ;
  assign n6318 = n564 & n5584 ;
  assign n6319 = n6317 | n6318 ;
  assign n6320 = n6316 | n6319 ;
  assign n6321 = n5418 | n6320 ;
  assign n6322 = ( ~n3492 & n6320 ) | ( ~n3492 & n6321 ) | ( n6320 & n6321 ) ;
  assign n6323 = x17 & ~n6322 ;
  assign n6324 = ~x17 & n6322 ;
  assign n6325 = n6323 | n6324 ;
  assign n6326 = ( ~n5876 & n5878 ) | ( ~n5876 & n5888 ) | ( n5878 & n5888 ) ;
  assign n6327 = ( n5876 & ~n5889 ) | ( n5876 & n6326 ) | ( ~n5889 & n6326 ) ;
  assign n6328 = ( n6315 & n6325 ) | ( n6315 & n6327 ) | ( n6325 & n6327 ) ;
  assign n6329 = ( ~n5889 & n5899 ) | ( ~n5889 & n5901 ) | ( n5899 & n5901 ) ;
  assign n6330 = ( n5889 & ~n5902 ) | ( n5889 & n6329 ) | ( ~n5902 & n6329 ) ;
  assign n6331 = n5904 & ~n5906 ;
  assign n6332 = ~n5911 & n6331 ;
  assign n6333 = ~n3516 & n6332 ;
  assign n6334 = x14 & n6333 ;
  assign n6335 = ~n3533 & n5909 ;
  assign n6336 = n5915 | n6335 ;
  assign n6337 = ( n3609 & n6335 ) | ( n3609 & n6336 ) | ( n6335 & n6336 ) ;
  assign n6338 = x14 & ~n6337 ;
  assign n6339 = ( ~x14 & n6333 ) | ( ~x14 & n6337 ) | ( n6333 & n6337 ) ;
  assign n6340 = ( ~n6334 & n6338 ) | ( ~n6334 & n6339 ) | ( n6338 & n6339 ) ;
  assign n6341 = ( n6328 & n6330 ) | ( n6328 & n6340 ) | ( n6330 & n6340 ) ;
  assign n6342 = ( ~n6231 & n6241 ) | ( ~n6231 & n6243 ) | ( n6241 & n6243 ) ;
  assign n6343 = ( n6231 & ~n6244 ) | ( n6231 & n6342 ) | ( ~n6244 & n6342 ) ;
  assign n6344 = ~n2041 & n4215 ;
  assign n6345 = n2083 & n2187 ;
  assign n6346 = n6344 | n6345 ;
  assign n6347 = n2102 & n4200 ;
  assign n6348 = n6346 | n6347 ;
  assign n6349 = x26 & n6348 ;
  assign n6350 = n4203 & ~n4997 ;
  assign n6351 = x26 & ~n6350 ;
  assign n6352 = ( ~x26 & n6348 ) | ( ~x26 & n6350 ) | ( n6348 & n6350 ) ;
  assign n6353 = ( ~n6349 & n6351 ) | ( ~n6349 & n6352 ) | ( n6351 & n6352 ) ;
  assign n6354 = n2102 & n4215 ;
  assign n6355 = n2187 & n4200 ;
  assign n6356 = n6354 | n6355 ;
  assign n6357 = n2083 & ~n2282 ;
  assign n6358 = n6356 | n6357 ;
  assign n6359 = n4203 | n6358 ;
  assign n6360 = ( ~n5331 & n6358 ) | ( ~n5331 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6361 = x26 & ~n6360 ;
  assign n6362 = ~x26 & n6360 ;
  assign n6363 = n6361 | n6362 ;
  assign n6364 = ~n2364 & n4039 ;
  assign n6365 = n2398 & n3501 ;
  assign n6366 = n6364 | n6365 ;
  assign n6367 = n3541 | n6366 ;
  assign n6368 = ( n5713 & n6366 ) | ( n5713 & n6367 ) | ( n6366 & n6367 ) ;
  assign n6369 = ~n2467 & n3536 ;
  assign n6370 = n6368 | n6369 ;
  assign n6371 = x29 & ~n6370 ;
  assign n6372 = ~x29 & n6370 ;
  assign n6373 = n6371 | n6372 ;
  assign n6374 = ( n6218 & n6228 ) | ( n6218 & n6230 ) | ( n6228 & n6230 ) ;
  assign n6375 = ( n6230 & n6231 ) | ( n6230 & ~n6374 ) | ( n6231 & ~n6374 ) ;
  assign n6376 = ( n6363 & n6373 ) | ( n6363 & ~n6375 ) | ( n6373 & ~n6375 ) ;
  assign n6377 = ( n6343 & n6353 ) | ( n6343 & n6376 ) | ( n6353 & n6376 ) ;
  assign n6378 = n1687 & n4649 ;
  assign n6379 = n1792 & n4637 ;
  assign n6380 = n6378 | n6379 ;
  assign n6381 = ~n1841 & n4584 ;
  assign n6382 = n6380 | n6381 ;
  assign n6383 = x23 & n6382 ;
  assign n6384 = n4331 & n4591 ;
  assign n6385 = x23 & ~n6384 ;
  assign n6386 = ( ~x23 & n6382 ) | ( ~x23 & n6384 ) | ( n6382 & n6384 ) ;
  assign n6387 = ( ~n6383 & n6385 ) | ( ~n6383 & n6386 ) | ( n6385 & n6386 ) ;
  assign n6388 = ( ~n6244 & n6254 ) | ( ~n6244 & n6256 ) | ( n6254 & n6256 ) ;
  assign n6389 = ( ~n6254 & n6257 ) | ( ~n6254 & n6388 ) | ( n6257 & n6388 ) ;
  assign n6390 = ( n6377 & n6387 ) | ( n6377 & ~n6389 ) | ( n6387 & ~n6389 ) ;
  assign n6391 = n1398 & n5232 ;
  assign n6392 = n4874 | n6391 ;
  assign n6393 = ( ~n1529 & n6391 ) | ( ~n1529 & n6392 ) | ( n6391 & n6392 ) ;
  assign n6394 = n1316 & n4878 ;
  assign n6395 = n6393 | n6394 ;
  assign n6396 = n4879 | n6395 ;
  assign n6397 = ( n4084 & n6395 ) | ( n4084 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = x20 & ~n6397 ;
  assign n6399 = ~x20 & n6397 ;
  assign n6400 = n6398 | n6399 ;
  assign n6401 = ( ~n6257 & n6267 ) | ( ~n6257 & n6275 ) | ( n6267 & n6275 ) ;
  assign n6402 = ( n6257 & ~n6276 ) | ( n6257 & n6401 ) | ( ~n6276 & n6401 ) ;
  assign n6403 = ( n6390 & n6400 ) | ( n6390 & n6402 ) | ( n6400 & n6402 ) ;
  assign n6404 = ( ~n6276 & n6278 ) | ( ~n6276 & n6288 ) | ( n6278 & n6288 ) ;
  assign n6405 = ( n6276 & ~n6289 ) | ( n6276 & n6404 ) | ( ~n6289 & n6404 ) ;
  assign n6406 = n1398 & n4874 ;
  assign n6407 = n5232 | n6406 ;
  assign n6408 = ( n1316 & n6406 ) | ( n1316 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6409 = ~n1207 & n4878 ;
  assign n6410 = n6408 | n6409 ;
  assign n6411 = n4879 | n6410 ;
  assign n6412 = ( ~n4157 & n6410 ) | ( ~n4157 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6413 = x20 & ~n6412 ;
  assign n6414 = ~x20 & n6412 ;
  assign n6415 = n6413 | n6414 ;
  assign n6416 = ( n6403 & n6405 ) | ( n6403 & n6415 ) | ( n6405 & n6415 ) ;
  assign n6417 = ( ~n6289 & n6299 ) | ( ~n6289 & n6301 ) | ( n6299 & n6301 ) ;
  assign n6418 = ( n6289 & ~n6302 ) | ( n6289 & n6417 ) | ( ~n6302 & n6417 ) ;
  assign n6419 = n859 & n5584 ;
  assign n6420 = ~n721 & n5417 ;
  assign n6421 = n6419 | n6420 ;
  assign n6422 = n995 & n5413 ;
  assign n6423 = n6421 | n6422 ;
  assign n6424 = n5418 | n6423 ;
  assign n6425 = ( ~n3829 & n6423 ) | ( ~n3829 & n6424 ) | ( n6423 & n6424 ) ;
  assign n6426 = x17 & ~n6425 ;
  assign n6427 = ~x17 & n6425 ;
  assign n6428 = n6426 | n6427 ;
  assign n6429 = ( n6416 & n6418 ) | ( n6416 & n6428 ) | ( n6418 & n6428 ) ;
  assign n6430 = ( ~n6302 & n6312 ) | ( ~n6302 & n6314 ) | ( n6312 & n6314 ) ;
  assign n6431 = ( n6302 & ~n6315 ) | ( n6302 & n6430 ) | ( ~n6315 & n6430 ) ;
  assign n6432 = ~n3487 & n5909 ;
  assign n6433 = x14 & n6432 ;
  assign n6434 = ~n3601 & n6332 ;
  assign n6435 = ~n3533 & n5914 ;
  assign n6436 = n6434 | n6435 ;
  assign n6437 = n5915 | n6436 ;
  assign n6438 = ( ~n4223 & n6436 ) | ( ~n4223 & n6437 ) | ( n6436 & n6437 ) ;
  assign n6439 = x14 & ~n6438 ;
  assign n6440 = ( ~x14 & n6432 ) | ( ~x14 & n6438 ) | ( n6432 & n6438 ) ;
  assign n6441 = ( ~n6433 & n6439 ) | ( ~n6433 & n6440 ) | ( n6439 & n6440 ) ;
  assign n6442 = ( n6429 & n6431 ) | ( n6429 & n6441 ) | ( n6431 & n6441 ) ;
  assign n6443 = ~n3516 & n5914 ;
  assign n6444 = n5909 | n6443 ;
  assign n6445 = ( ~n3601 & n6443 ) | ( ~n3601 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6446 = ~n3533 & n6332 ;
  assign n6447 = n6445 | n6446 ;
  assign n6448 = n5915 | n6447 ;
  assign n6449 = ( ~n4058 & n6447 ) | ( ~n4058 & n6448 ) | ( n6447 & n6448 ) ;
  assign n6450 = x14 & ~n6449 ;
  assign n6451 = ~x14 & n6449 ;
  assign n6452 = n6450 | n6451 ;
  assign n6453 = ( ~n6315 & n6325 ) | ( ~n6315 & n6327 ) | ( n6325 & n6327 ) ;
  assign n6454 = ( n6315 & ~n6328 ) | ( n6315 & n6453 ) | ( ~n6328 & n6453 ) ;
  assign n6455 = ( n6442 & n6452 ) | ( n6442 & n6454 ) | ( n6452 & n6454 ) ;
  assign n6456 = ( ~n6204 & n6207 ) | ( ~n6204 & n6217 ) | ( n6207 & n6217 ) ;
  assign n6457 = ( n6204 & ~n6218 ) | ( n6204 & n6456 ) | ( ~n6218 & n6456 ) ;
  assign n6458 = n2083 & ~n2364 ;
  assign n6459 = n2187 & n4215 ;
  assign n6460 = n6458 | n6459 ;
  assign n6461 = ~n2282 & n4200 ;
  assign n6462 = n6460 | n6461 ;
  assign n6463 = x26 & n6462 ;
  assign n6464 = n4203 & n5137 ;
  assign n6465 = x26 & ~n6464 ;
  assign n6466 = ( ~x26 & n6462 ) | ( ~x26 & n6464 ) | ( n6462 & n6464 ) ;
  assign n6467 = ( ~n6463 & n6465 ) | ( ~n6463 & n6466 ) | ( n6465 & n6466 ) ;
  assign n6468 = ~n2467 & n3501 ;
  assign n6469 = ~n2521 & n3536 ;
  assign n6470 = n2398 & n4039 ;
  assign n6471 = n6469 | n6470 ;
  assign n6472 = n6468 | n6471 ;
  assign n6473 = x29 & n6472 ;
  assign n6474 = n3541 & n5452 ;
  assign n6475 = x29 & ~n6474 ;
  assign n6476 = ( ~x29 & n6472 ) | ( ~x29 & n6474 ) | ( n6472 & n6474 ) ;
  assign n6477 = ( ~n6473 & n6475 ) | ( ~n6473 & n6476 ) | ( n6475 & n6476 ) ;
  assign n6478 = ( n6457 & n6467 ) | ( n6457 & n6477 ) | ( n6467 & n6477 ) ;
  assign n6479 = ~n2041 & n4584 ;
  assign n6480 = x23 & n6479 ;
  assign n6481 = ~n1841 & n4649 ;
  assign n6482 = n1943 & n4637 ;
  assign n6483 = n6481 | n6482 ;
  assign n6484 = n4591 | n6483 ;
  assign n6485 = ( ~n4753 & n6483 ) | ( ~n4753 & n6484 ) | ( n6483 & n6484 ) ;
  assign n6486 = x23 & ~n6485 ;
  assign n6487 = ( ~x23 & n6479 ) | ( ~x23 & n6485 ) | ( n6479 & n6485 ) ;
  assign n6488 = ( ~n6480 & n6486 ) | ( ~n6480 & n6487 ) | ( n6486 & n6487 ) ;
  assign n6489 = ~n6269 & n6368 ;
  assign n6490 = n6269 | n6368 ;
  assign n6491 = ( ~n6370 & n6489 ) | ( ~n6370 & n6490 ) | ( n6489 & n6490 ) ;
  assign n6492 = ( n6360 & ~n6375 ) | ( n6360 & n6491 ) | ( ~n6375 & n6491 ) ;
  assign n6493 = ( n6360 & n6375 ) | ( n6360 & n6491 ) | ( n6375 & n6491 ) ;
  assign n6494 = ( n6375 & n6492 ) | ( n6375 & ~n6493 ) | ( n6492 & ~n6493 ) ;
  assign n6495 = ( n6478 & n6488 ) | ( n6478 & ~n6494 ) | ( n6488 & ~n6494 ) ;
  assign n6496 = n1792 & n4649 ;
  assign n6497 = x23 & n6496 ;
  assign n6498 = ~n1841 & n4637 ;
  assign n6499 = n1943 & n4584 ;
  assign n6500 = n6498 | n6499 ;
  assign n6501 = n4591 | n6500 ;
  assign n6502 = ( ~n4831 & n6500 ) | ( ~n4831 & n6501 ) | ( n6500 & n6501 ) ;
  assign n6503 = x23 & ~n6502 ;
  assign n6504 = ( ~x23 & n6496 ) | ( ~x23 & n6502 ) | ( n6496 & n6502 ) ;
  assign n6505 = ( ~n6497 & n6503 ) | ( ~n6497 & n6504 ) | ( n6503 & n6504 ) ;
  assign n6506 = ( ~n6343 & n6353 ) | ( ~n6343 & n6376 ) | ( n6353 & n6376 ) ;
  assign n6507 = ( n6343 & ~n6377 ) | ( n6343 & n6506 ) | ( ~n6377 & n6506 ) ;
  assign n6508 = ( n6495 & n6505 ) | ( n6495 & n6507 ) | ( n6505 & n6507 ) ;
  assign n6509 = ~n1529 & n5232 ;
  assign n6510 = n1600 & n4874 ;
  assign n6511 = n1398 & n4878 ;
  assign n6512 = n6510 | n6511 ;
  assign n6513 = n6509 | n6512 ;
  assign n6514 = n4879 | n6513 ;
  assign n6515 = ( ~n4324 & n6513 ) | ( ~n4324 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6516 = x20 & ~n6515 ;
  assign n6517 = ~x20 & n6515 ;
  assign n6518 = n6516 | n6517 ;
  assign n6519 = ( ~n6377 & n6387 ) | ( ~n6377 & n6389 ) | ( n6387 & n6389 ) ;
  assign n6520 = ( ~n6387 & n6390 ) | ( ~n6387 & n6519 ) | ( n6390 & n6519 ) ;
  assign n6521 = ( n6508 & n6518 ) | ( n6508 & ~n6520 ) | ( n6518 & ~n6520 ) ;
  assign n6522 = n995 & n5417 ;
  assign n6523 = ~n1207 & n5413 ;
  assign n6524 = n6522 | n6523 ;
  assign n6525 = ~n1118 & n5584 ;
  assign n6526 = n6524 | n6525 ;
  assign n6527 = n5418 | n6526 ;
  assign n6528 = ( n4173 & n6526 ) | ( n4173 & n6527 ) | ( n6526 & n6527 ) ;
  assign n6529 = x17 & ~n6528 ;
  assign n6530 = ~x17 & n6528 ;
  assign n6531 = n6529 | n6530 ;
  assign n6532 = ( ~n6390 & n6400 ) | ( ~n6390 & n6402 ) | ( n6400 & n6402 ) ;
  assign n6533 = ( n6390 & ~n6403 ) | ( n6390 & n6532 ) | ( ~n6403 & n6532 ) ;
  assign n6534 = ( n6521 & n6531 ) | ( n6521 & n6533 ) | ( n6531 & n6533 ) ;
  assign n6535 = ( ~n6403 & n6405 ) | ( ~n6403 & n6415 ) | ( n6405 & n6415 ) ;
  assign n6536 = ( n6403 & ~n6416 ) | ( n6403 & n6535 ) | ( ~n6416 & n6535 ) ;
  assign n6537 = n995 & n5584 ;
  assign n6538 = x17 & n6537 ;
  assign n6539 = n859 & n5417 ;
  assign n6540 = ~n1118 & n5413 ;
  assign n6541 = n6539 | n6540 ;
  assign n6542 = n5418 | n6541 ;
  assign n6543 = ( ~n4034 & n6541 ) | ( ~n4034 & n6542 ) | ( n6541 & n6542 ) ;
  assign n6544 = x17 & ~n6543 ;
  assign n6545 = ( ~x17 & n6537 ) | ( ~x17 & n6543 ) | ( n6537 & n6543 ) ;
  assign n6546 = ( ~n6538 & n6544 ) | ( ~n6538 & n6545 ) | ( n6544 & n6545 ) ;
  assign n6547 = ( n6534 & n6536 ) | ( n6534 & n6546 ) | ( n6536 & n6546 ) ;
  assign n6548 = ~n3601 & n5914 ;
  assign n6549 = n564 & n5909 ;
  assign n6550 = n6548 | n6549 ;
  assign n6551 = ~n3487 & n6332 ;
  assign n6552 = n6550 | n6551 ;
  assign n6553 = n5915 | n6552 ;
  assign n6554 = ( n3674 & n6552 ) | ( n3674 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = x14 & ~n6554 ;
  assign n6556 = ~x14 & n6554 ;
  assign n6557 = n6555 | n6556 ;
  assign n6558 = ( ~n6416 & n6418 ) | ( ~n6416 & n6428 ) | ( n6418 & n6428 ) ;
  assign n6559 = ( n6416 & ~n6429 ) | ( n6416 & n6558 ) | ( ~n6429 & n6558 ) ;
  assign n6560 = ( n6547 & n6557 ) | ( n6547 & n6559 ) | ( n6557 & n6559 ) ;
  assign n6561 = x8 & x9 ;
  assign n6562 = x10 & n6561 ;
  assign n6563 = ~x11 & n6562 ;
  assign n6564 = x8 | x9 ;
  assign n6565 = x10 | n6564 ;
  assign n6566 = x10 | x11 ;
  assign n6567 = ( n6563 & ~n6565 ) | ( n6563 & n6566 ) | ( ~n6565 & n6566 ) ;
  assign n6568 = ~n6561 & n6564 ;
  assign n6569 = x10 & x11 ;
  assign n6570 = ( ~n6566 & n6568 ) | ( ~n6566 & n6569 ) | ( n6568 & n6569 ) ;
  assign n6571 = n6568 & ~n6570 ;
  assign n6572 = ( ~n3516 & n3608 ) | ( ~n3516 & n6571 ) | ( n3608 & n6571 ) ;
  assign n6573 = ( ~n3607 & n6567 ) | ( ~n3607 & n6572 ) | ( n6567 & n6572 ) ;
  assign n6574 = x11 & ~n6573 ;
  assign n6575 = ~x11 & n6573 ;
  assign n6576 = n6574 | n6575 ;
  assign n6577 = ( ~n6429 & n6431 ) | ( ~n6429 & n6441 ) | ( n6431 & n6441 ) ;
  assign n6578 = ( n6429 & ~n6442 ) | ( n6429 & n6577 ) | ( ~n6442 & n6577 ) ;
  assign n6579 = ( n6560 & n6576 ) | ( n6560 & n6578 ) | ( n6576 & n6578 ) ;
  assign n6580 = n3123 & n3536 ;
  assign n6581 = ~n2977 & n3501 ;
  assign n6582 = n6580 | n6581 ;
  assign n6583 = ~n2944 & n4039 ;
  assign n6584 = n6582 | n6583 ;
  assign n6585 = x29 & n6584 ;
  assign n6586 = n3541 & ~n5926 ;
  assign n6587 = x29 & ~n6586 ;
  assign n6588 = ( ~x29 & n6584 ) | ( ~x29 & n6586 ) | ( n6584 & n6586 ) ;
  assign n6589 = ( ~n6585 & n6587 ) | ( ~n6585 & n6588 ) | ( n6587 & n6588 ) ;
  assign n6590 = n389 & n3233 ;
  assign n6591 = ( x29 & x30 ) | ( x29 & ~n3049 ) | ( x30 & ~n3049 ) ;
  assign n6592 = ( x31 & ~n3232 ) | ( x31 & n6591 ) | ( ~n3232 & n6591 ) ;
  assign n6593 = x31 & n6591 ;
  assign n6594 = ( n6590 & n6592 ) | ( n6590 & ~n6593 ) | ( n6592 & ~n6593 ) ;
  assign n6595 = n3541 & n5965 ;
  assign n6596 = n3123 & n4039 ;
  assign n6597 = ~n3049 & n3501 ;
  assign n6598 = n6596 | n6597 ;
  assign n6599 = ~n3232 & n3536 ;
  assign n6600 = n6598 | n6599 ;
  assign n6601 = n6595 | n6600 ;
  assign n6602 = ~n3232 & n3500 ;
  assign n6603 = ~n3049 & n3500 ;
  assign n6604 = n3232 & ~n6603 ;
  assign n6605 = n3501 | n3541 ;
  assign n6606 = ( n3232 & n6603 ) | ( n3232 & ~n6605 ) | ( n6603 & ~n6605 ) ;
  assign n6607 = ~n6603 & n6605 ;
  assign n6608 = ( ~n6604 & n6606 ) | ( ~n6604 & n6607 ) | ( n6606 & n6607 ) ;
  assign n6609 = n6602 | n6608 ;
  assign n6610 = x29 & ~n6609 ;
  assign n6611 = ~n6601 & n6610 ;
  assign n6612 = n57 & ~n3232 ;
  assign n6613 = n6611 | n6612 ;
  assign n6614 = n3123 & n3501 ;
  assign n6615 = ~n3049 & n3536 ;
  assign n6616 = n6614 | n6615 ;
  assign n6617 = ~n2977 & n4039 ;
  assign n6618 = n6616 | n6617 ;
  assign n6619 = n3541 | n6618 ;
  assign n6620 = ( n6000 & n6618 ) | ( n6000 & n6619 ) | ( n6618 & n6619 ) ;
  assign n6621 = n42 & ~n3232 ;
  assign n6622 = n6620 & n6621 ;
  assign n6623 = n6620 & ~n6621 ;
  assign n6624 = ( n6613 & n6622 ) | ( n6613 & ~n6623 ) | ( n6622 & ~n6623 ) ;
  assign n6625 = ( n6589 & n6594 ) | ( n6589 & n6624 ) | ( n6594 & n6624 ) ;
  assign n6626 = ~n2888 & n4039 ;
  assign n6627 = ~n2977 & n3536 ;
  assign n6628 = ~n2944 & n3501 ;
  assign n6629 = n6627 | n6628 ;
  assign n6630 = n6626 | n6629 ;
  assign n6631 = x29 & n6630 ;
  assign n6632 = n3541 & ~n6055 ;
  assign n6633 = x29 & ~n6632 ;
  assign n6634 = ( ~x29 & n6630 ) | ( ~x29 & n6632 ) | ( n6630 & n6632 ) ;
  assign n6635 = ( ~n6631 & n6633 ) | ( ~n6631 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6636 = ~n5972 & n5995 ;
  assign n6637 = n5996 | n6636 ;
  assign n6638 = ( n6625 & n6635 ) | ( n6625 & ~n6637 ) | ( n6635 & ~n6637 ) ;
  assign n6639 = ~n2888 & n3501 ;
  assign n6640 = n2820 & n4039 ;
  assign n6641 = ~n2944 & n3536 ;
  assign n6642 = n6640 | n6641 ;
  assign n6643 = n6639 | n6642 ;
  assign n6644 = n3541 | n6643 ;
  assign n6645 = ( n6106 & n6643 ) | ( n6106 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = x29 & ~n6645 ;
  assign n6647 = ~x29 & n6645 ;
  assign n6648 = n6646 | n6647 ;
  assign n6649 = ( n5996 & ~n6007 ) | ( n5996 & n6049 ) | ( ~n6007 & n6049 ) ;
  assign n6650 = ( ~n5996 & n6050 ) | ( ~n5996 & n6649 ) | ( n6050 & n6649 ) ;
  assign n6651 = ( n6638 & n6648 ) | ( n6638 & ~n6650 ) | ( n6648 & ~n6650 ) ;
  assign n6652 = n2735 & n4039 ;
  assign n6653 = n2820 & n3501 ;
  assign n6654 = n6652 | n6653 ;
  assign n6655 = ~n2888 & n3536 ;
  assign n6656 = n6654 | n6655 ;
  assign n6657 = n3541 | n6656 ;
  assign n6658 = ( ~n6157 & n6656 ) | ( ~n6157 & n6657 ) | ( n6656 & n6657 ) ;
  assign n6659 = x29 & ~n6658 ;
  assign n6660 = ~x29 & n6658 ;
  assign n6661 = n6659 | n6660 ;
  assign n6662 = ( ~n5933 & n5963 ) | ( ~n5933 & n6050 ) | ( n5963 & n6050 ) ;
  assign n6663 = ( n5933 & ~n6051 ) | ( n5933 & n6662 ) | ( ~n6051 & n6662 ) ;
  assign n6664 = ( n6651 & n6661 ) | ( n6651 & n6663 ) | ( n6661 & n6663 ) ;
  assign n6665 = ( n6051 & ~n6062 ) | ( n6051 & n6102 ) | ( ~n6062 & n6102 ) ;
  assign n6666 = ( ~n6051 & n6103 ) | ( ~n6051 & n6665 ) | ( n6103 & n6665 ) ;
  assign n6667 = n2820 & n3536 ;
  assign n6668 = n2642 & n4039 ;
  assign n6669 = n6667 | n6668 ;
  assign n6670 = n2735 & n3501 ;
  assign n6671 = n6669 | n6670 ;
  assign n6672 = x29 & n6671 ;
  assign n6673 = n3541 & n5598 ;
  assign n6674 = x29 & ~n6673 ;
  assign n6675 = ( ~x29 & n6671 ) | ( ~x29 & n6673 ) | ( n6671 & n6673 ) ;
  assign n6676 = ( ~n6672 & n6674 ) | ( ~n6672 & n6675 ) | ( n6674 & n6675 ) ;
  assign n6677 = ( n6664 & ~n6666 ) | ( n6664 & n6676 ) | ( ~n6666 & n6676 ) ;
  assign n6678 = n2642 & n3501 ;
  assign n6679 = ~n2608 & n4039 ;
  assign n6680 = n6678 | n6679 ;
  assign n6681 = n2735 & n3536 ;
  assign n6682 = n6680 | n6681 ;
  assign n6683 = n3541 | n6682 ;
  assign n6684 = ( ~n6216 & n6682 ) | ( ~n6216 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6685 = x29 & ~n6684 ;
  assign n6686 = ~x29 & n6684 ;
  assign n6687 = n6685 | n6686 ;
  assign n6688 = ( ~n6103 & n6113 ) | ( ~n6103 & n6147 ) | ( n6113 & n6147 ) ;
  assign n6689 = ( n6103 & ~n6148 ) | ( n6103 & n6688 ) | ( ~n6148 & n6688 ) ;
  assign n6690 = ( n6677 & n6687 ) | ( n6677 & n6689 ) | ( n6687 & n6689 ) ;
  assign n6691 = n2642 & n3536 ;
  assign n6692 = ~n2608 & n3501 ;
  assign n6693 = n6691 | n6692 ;
  assign n6694 = ~n2521 & n4039 ;
  assign n6695 = n6693 | n6694 ;
  assign n6696 = x29 & n6695 ;
  assign n6697 = n3541 & n6221 ;
  assign n6698 = x29 & ~n6697 ;
  assign n6699 = ( ~x29 & n6695 ) | ( ~x29 & n6697 ) | ( n6695 & n6697 ) ;
  assign n6700 = ( ~n6696 & n6698 ) | ( ~n6696 & n6699 ) | ( n6698 & n6699 ) ;
  assign n6701 = ( ~n6148 & n6158 ) | ( ~n6148 & n6189 ) | ( n6158 & n6189 ) ;
  assign n6702 = ( n6148 & ~n6190 ) | ( n6148 & n6701 ) | ( ~n6190 & n6701 ) ;
  assign n6703 = ( n6690 & n6700 ) | ( n6690 & n6702 ) | ( n6700 & n6702 ) ;
  assign n6704 = ( ~n6190 & n6200 ) | ( ~n6190 & n6203 ) | ( n6200 & n6203 ) ;
  assign n6705 = ( n6190 & ~n6204 ) | ( n6190 & n6704 ) | ( ~n6204 & n6704 ) ;
  assign n6706 = ~n2364 & n4200 ;
  assign n6707 = ~n2282 & n4215 ;
  assign n6708 = n6706 | n6707 ;
  assign n6709 = n2083 & n2398 ;
  assign n6710 = n6708 | n6709 ;
  assign n6711 = n4203 | n6710 ;
  assign n6712 = ( ~n5494 & n6710 ) | ( ~n5494 & n6711 ) | ( n6710 & n6711 ) ;
  assign n6713 = x26 & ~n6712 ;
  assign n6714 = ~x26 & n6712 ;
  assign n6715 = n6713 | n6714 ;
  assign n6716 = ( n6703 & n6705 ) | ( n6703 & n6715 ) | ( n6705 & n6715 ) ;
  assign n6717 = ~n2041 & n4637 ;
  assign n6718 = x23 & n6717 ;
  assign n6719 = n1943 & n4649 ;
  assign n6720 = n2102 & n4584 ;
  assign n6721 = n6719 | n6720 ;
  assign n6722 = n4591 | n6721 ;
  assign n6723 = ( ~n4985 & n6721 ) | ( ~n4985 & n6722 ) | ( n6721 & n6722 ) ;
  assign n6724 = x23 & ~n6723 ;
  assign n6725 = ( ~x23 & n6717 ) | ( ~x23 & n6723 ) | ( n6717 & n6723 ) ;
  assign n6726 = ( ~n6718 & n6724 ) | ( ~n6718 & n6725 ) | ( n6724 & n6725 ) ;
  assign n6727 = ( ~n6457 & n6467 ) | ( ~n6457 & n6477 ) | ( n6467 & n6477 ) ;
  assign n6728 = ( n6457 & ~n6478 ) | ( n6457 & n6727 ) | ( ~n6478 & n6727 ) ;
  assign n6729 = ( n6716 & n6726 ) | ( n6716 & n6728 ) | ( n6726 & n6728 ) ;
  assign n6730 = ( n6478 & ~n6488 ) | ( n6478 & n6494 ) | ( ~n6488 & n6494 ) ;
  assign n6731 = ( ~n6478 & n6495 ) | ( ~n6478 & n6730 ) | ( n6495 & n6730 ) ;
  assign n6732 = n1687 & n5232 ;
  assign n6733 = n1792 & n4874 ;
  assign n6734 = n1600 & n4878 ;
  assign n6735 = n6733 | n6734 ;
  assign n6736 = n6732 | n6735 ;
  assign n6737 = n4879 | n6736 ;
  assign n6738 = ( n4674 & n6736 ) | ( n4674 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6739 = x20 & ~n6738 ;
  assign n6740 = ~x20 & n6738 ;
  assign n6741 = n6739 | n6740 ;
  assign n6742 = ( n6729 & ~n6731 ) | ( n6729 & n6741 ) | ( ~n6731 & n6741 ) ;
  assign n6743 = ( ~n6495 & n6505 ) | ( ~n6495 & n6507 ) | ( n6505 & n6507 ) ;
  assign n6744 = ( n6495 & ~n6508 ) | ( n6495 & n6743 ) | ( ~n6508 & n6743 ) ;
  assign n6745 = ~n1529 & n4878 ;
  assign n6746 = n1687 & n4874 ;
  assign n6747 = n6745 | n6746 ;
  assign n6748 = n1600 & n5232 ;
  assign n6749 = n6747 | n6748 ;
  assign n6750 = n4879 | n6749 ;
  assign n6751 = ( ~n4531 & n6749 ) | ( ~n4531 & n6750 ) | ( n6749 & n6750 ) ;
  assign n6752 = x20 & ~n6751 ;
  assign n6753 = ~x20 & n6751 ;
  assign n6754 = n6752 | n6753 ;
  assign n6755 = ( n6742 & n6744 ) | ( n6742 & n6754 ) | ( n6744 & n6754 ) ;
  assign n6756 = n1316 & n5413 ;
  assign n6757 = ~n1207 & n5584 ;
  assign n6758 = n6756 | n6757 ;
  assign n6759 = ~n1118 & n5417 ;
  assign n6760 = n6758 | n6759 ;
  assign n6761 = n5418 | n6760 ;
  assign n6762 = ( n3841 & n6760 ) | ( n3841 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6763 = x17 & ~n6762 ;
  assign n6764 = ~x17 & n6762 ;
  assign n6765 = n6763 | n6764 ;
  assign n6766 = ( ~n6508 & n6518 ) | ( ~n6508 & n6520 ) | ( n6518 & n6520 ) ;
  assign n6767 = ( ~n6518 & n6521 ) | ( ~n6518 & n6766 ) | ( n6521 & n6766 ) ;
  assign n6768 = ( n6755 & n6765 ) | ( n6755 & ~n6767 ) | ( n6765 & ~n6767 ) ;
  assign n6769 = ( ~n6521 & n6531 ) | ( ~n6521 & n6533 ) | ( n6531 & n6533 ) ;
  assign n6770 = ( n6521 & ~n6534 ) | ( n6521 & n6769 ) | ( ~n6534 & n6769 ) ;
  assign n6771 = ~n721 & n6332 ;
  assign n6772 = x14 & n6771 ;
  assign n6773 = n564 & n5914 ;
  assign n6774 = n859 & n5909 ;
  assign n6775 = n6773 | n6774 ;
  assign n6776 = n5915 | n6775 ;
  assign n6777 = ( ~n3268 & n6775 ) | ( ~n3268 & n6776 ) | ( n6775 & n6776 ) ;
  assign n6778 = x14 & ~n6777 ;
  assign n6779 = ( ~x14 & n6771 ) | ( ~x14 & n6777 ) | ( n6771 & n6777 ) ;
  assign n6780 = ( ~n6772 & n6778 ) | ( ~n6772 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = ( n6768 & n6770 ) | ( n6768 & n6780 ) | ( n6770 & n6780 ) ;
  assign n6782 = ~n3487 & n5914 ;
  assign n6783 = ~n721 & n5909 ;
  assign n6784 = n564 & n6332 ;
  assign n6785 = n6783 | n6784 ;
  assign n6786 = n6782 | n6785 ;
  assign n6787 = n5915 | n6786 ;
  assign n6788 = ( ~n3492 & n6786 ) | ( ~n3492 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6789 = x14 & ~n6788 ;
  assign n6790 = ~x14 & n6788 ;
  assign n6791 = n6789 | n6790 ;
  assign n6792 = ( ~n6534 & n6536 ) | ( ~n6534 & n6546 ) | ( n6536 & n6546 ) ;
  assign n6793 = ( n6534 & ~n6547 ) | ( n6534 & n6792 ) | ( ~n6547 & n6792 ) ;
  assign n6794 = ( n6781 & n6791 ) | ( n6781 & n6793 ) | ( n6791 & n6793 ) ;
  assign n6795 = ~n6562 & n6565 ;
  assign n6796 = ~n6568 & n6795 ;
  assign n6797 = ~n3516 & n6796 ;
  assign n6798 = x11 & n6797 ;
  assign n6799 = ~n3533 & n6567 ;
  assign n6800 = n6571 | n6799 ;
  assign n6801 = ( n3609 & n6799 ) | ( n3609 & n6800 ) | ( n6799 & n6800 ) ;
  assign n6802 = x11 & ~n6801 ;
  assign n6803 = ( ~x11 & n6797 ) | ( ~x11 & n6801 ) | ( n6797 & n6801 ) ;
  assign n6804 = ( ~n6798 & n6802 ) | ( ~n6798 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6805 = ( ~n6547 & n6557 ) | ( ~n6547 & n6559 ) | ( n6557 & n6559 ) ;
  assign n6806 = ( n6547 & ~n6560 ) | ( n6547 & n6805 ) | ( ~n6560 & n6805 ) ;
  assign n6807 = ( n6794 & n6804 ) | ( n6794 & n6806 ) | ( n6804 & n6806 ) ;
  assign n6808 = ~n2944 & n4215 ;
  assign n6809 = ~n2977 & n4200 ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = n2083 & n3123 ;
  assign n6812 = n6810 | n6811 ;
  assign n6813 = n4203 | n6812 ;
  assign n6814 = ( ~n5926 & n6812 ) | ( ~n5926 & n6813 ) | ( n6812 & n6813 ) ;
  assign n6815 = x26 & ~n6814 ;
  assign n6816 = ~x26 & n6814 ;
  assign n6817 = n6815 | n6816 ;
  assign n6818 = ( x29 & n6602 ) | ( x29 & ~n6608 ) | ( n6602 & ~n6608 ) ;
  assign n6819 = x29 & ~n6608 ;
  assign n6820 = ( n6609 & ~n6818 ) | ( n6609 & n6819 ) | ( ~n6818 & n6819 ) ;
  assign n6821 = n3123 & n4200 ;
  assign n6822 = ~n2977 & n4215 ;
  assign n6823 = n6821 | n6822 ;
  assign n6824 = n2083 & ~n3049 ;
  assign n6825 = n6823 | n6824 ;
  assign n6826 = x26 & n6825 ;
  assign n6827 = n4203 & n6000 ;
  assign n6828 = x26 & ~n6827 ;
  assign n6829 = ( ~x26 & n6825 ) | ( ~x26 & n6827 ) | ( n6825 & n6827 ) ;
  assign n6830 = ( ~n6826 & n6828 ) | ( ~n6826 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6831 = n4203 & n5965 ;
  assign n6832 = n3123 & n4215 ;
  assign n6833 = ~n3049 & n4200 ;
  assign n6834 = n6832 | n6833 ;
  assign n6835 = n2083 & ~n3232 ;
  assign n6836 = n6834 | n6835 ;
  assign n6837 = n6831 | n6836 ;
  assign n6838 = n263 | n3232 ;
  assign n6839 = x25 | n72 ;
  assign n6840 = ~n6838 & n6839 ;
  assign n6841 = ~n3049 & n4202 ;
  assign n6842 = x26 & ~n6841 ;
  assign n6843 = ~n6840 & n6842 ;
  assign n6844 = ~n6837 & n6843 ;
  assign n6845 = ( n6602 & n6830 ) | ( n6602 & ~n6844 ) | ( n6830 & ~n6844 ) ;
  assign n6846 = n6602 & ~n6844 ;
  assign n6847 = ( n6602 & ~n6830 ) | ( n6602 & n6844 ) | ( ~n6830 & n6844 ) ;
  assign n6848 = ( n6845 & ~n6846 ) | ( n6845 & n6847 ) | ( ~n6846 & n6847 ) ;
  assign n6849 = ( n6602 & n6830 ) | ( n6602 & ~n6848 ) | ( n6830 & ~n6848 ) ;
  assign n6850 = ( n6817 & n6820 ) | ( n6817 & n6849 ) | ( n6820 & n6849 ) ;
  assign n6851 = ~n2888 & n4215 ;
  assign n6852 = n2083 & ~n2977 ;
  assign n6853 = ~n2944 & n4200 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = n6851 | n6854 ;
  assign n6856 = x26 & n6855 ;
  assign n6857 = n4203 & ~n6055 ;
  assign n6858 = x26 & ~n6857 ;
  assign n6859 = ( ~x26 & n6855 ) | ( ~x26 & n6857 ) | ( n6855 & n6857 ) ;
  assign n6860 = ( ~n6856 & n6858 ) | ( ~n6856 & n6859 ) | ( n6858 & n6859 ) ;
  assign n6861 = x29 & n6609 ;
  assign n6862 = ~n6601 & n6861 ;
  assign n6863 = n6601 & ~n6861 ;
  assign n6864 = n6862 | n6863 ;
  assign n6865 = ( n6850 & n6860 ) | ( n6850 & n6864 ) | ( n6860 & n6864 ) ;
  assign n6866 = n2083 & ~n2944 ;
  assign n6867 = n2820 & n4215 ;
  assign n6868 = n6866 | n6867 ;
  assign n6869 = ~n2888 & n4200 ;
  assign n6870 = n6868 | n6869 ;
  assign n6871 = n4203 | n6870 ;
  assign n6872 = ( n6106 & n6870 ) | ( n6106 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = x26 & ~n6872 ;
  assign n6874 = ~x26 & n6872 ;
  assign n6875 = n6873 | n6874 ;
  assign n6876 = n389 & ~n3232 ;
  assign n6877 = x29 & ~n6611 ;
  assign n6878 = ( n6620 & n6876 ) | ( n6620 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6879 = ( ~n6620 & n6876 ) | ( ~n6620 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6880 = ( n6620 & ~n6878 ) | ( n6620 & n6879 ) | ( ~n6878 & n6879 ) ;
  assign n6881 = ( n6865 & n6875 ) | ( n6865 & n6880 ) | ( n6875 & n6880 ) ;
  assign n6882 = n2820 & n4200 ;
  assign n6883 = x26 & n6882 ;
  assign n6884 = n2735 & n4215 ;
  assign n6885 = n2083 & ~n2888 ;
  assign n6886 = n6884 | n6885 ;
  assign n6887 = n4203 | n6886 ;
  assign n6888 = ( ~n6157 & n6886 ) | ( ~n6157 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6889 = x26 & ~n6888 ;
  assign n6890 = ( ~x26 & n6882 ) | ( ~x26 & n6888 ) | ( n6882 & n6888 ) ;
  assign n6891 = ( ~n6883 & n6889 ) | ( ~n6883 & n6890 ) | ( n6889 & n6890 ) ;
  assign n6892 = ( ~n6589 & n6594 ) | ( ~n6589 & n6624 ) | ( n6594 & n6624 ) ;
  assign n6893 = ( n6589 & ~n6625 ) | ( n6589 & n6892 ) | ( ~n6625 & n6892 ) ;
  assign n6894 = ( n6881 & n6891 ) | ( n6881 & n6893 ) | ( n6891 & n6893 ) ;
  assign n6895 = ( n6625 & ~n6635 ) | ( n6625 & n6637 ) | ( ~n6635 & n6637 ) ;
  assign n6896 = ( ~n6625 & n6638 ) | ( ~n6625 & n6895 ) | ( n6638 & n6895 ) ;
  assign n6897 = n2083 & n2820 ;
  assign n6898 = n2642 & n4215 ;
  assign n6899 = n6897 | n6898 ;
  assign n6900 = n2735 & n4200 ;
  assign n6901 = n6899 | n6900 ;
  assign n6902 = n4203 | n6901 ;
  assign n6903 = ( n5598 & n6901 ) | ( n5598 & n6902 ) | ( n6901 & n6902 ) ;
  assign n6904 = x26 & ~n6903 ;
  assign n6905 = ~x26 & n6903 ;
  assign n6906 = n6904 | n6905 ;
  assign n6907 = ( n6894 & ~n6896 ) | ( n6894 & n6906 ) | ( ~n6896 & n6906 ) ;
  assign n6908 = ( n6638 & ~n6648 ) | ( n6638 & n6650 ) | ( ~n6648 & n6650 ) ;
  assign n6909 = ( ~n6638 & n6651 ) | ( ~n6638 & n6908 ) | ( n6651 & n6908 ) ;
  assign n6910 = n2083 & n2735 ;
  assign n6911 = n2642 & n4200 ;
  assign n6912 = ~n2608 & n4215 ;
  assign n6913 = n6911 | n6912 ;
  assign n6914 = n6910 | n6913 ;
  assign n6915 = x26 & n6914 ;
  assign n6916 = n4203 & ~n6216 ;
  assign n6917 = x26 & ~n6916 ;
  assign n6918 = ( ~x26 & n6914 ) | ( ~x26 & n6916 ) | ( n6914 & n6916 ) ;
  assign n6919 = ( ~n6915 & n6917 ) | ( ~n6915 & n6918 ) | ( n6917 & n6918 ) ;
  assign n6920 = ( n6907 & ~n6909 ) | ( n6907 & n6919 ) | ( ~n6909 & n6919 ) ;
  assign n6921 = ( ~n6651 & n6661 ) | ( ~n6651 & n6663 ) | ( n6661 & n6663 ) ;
  assign n6922 = ( n6651 & ~n6664 ) | ( n6651 & n6921 ) | ( ~n6664 & n6921 ) ;
  assign n6923 = n2083 & n2642 ;
  assign n6924 = ~n2608 & n4200 ;
  assign n6925 = n6923 | n6924 ;
  assign n6926 = ~n2521 & n4215 ;
  assign n6927 = n6925 | n6926 ;
  assign n6928 = x26 & n6927 ;
  assign n6929 = n4203 & n6221 ;
  assign n6930 = x26 & ~n6929 ;
  assign n6931 = ( ~x26 & n6927 ) | ( ~x26 & n6929 ) | ( n6927 & n6929 ) ;
  assign n6932 = ( ~n6928 & n6930 ) | ( ~n6928 & n6931 ) | ( n6930 & n6931 ) ;
  assign n6933 = ( n6920 & n6922 ) | ( n6920 & n6932 ) | ( n6922 & n6932 ) ;
  assign n6934 = ~n2467 & n4215 ;
  assign n6935 = x26 & n6934 ;
  assign n6936 = ~n2521 & n4200 ;
  assign n6937 = n2083 & ~n2608 ;
  assign n6938 = n6936 | n6937 ;
  assign n6939 = n4203 | n6938 ;
  assign n6940 = ( ~n5693 & n6938 ) | ( ~n5693 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6941 = x26 & ~n6940 ;
  assign n6942 = ( ~x26 & n6934 ) | ( ~x26 & n6940 ) | ( n6934 & n6940 ) ;
  assign n6943 = ( ~n6935 & n6941 ) | ( ~n6935 & n6942 ) | ( n6941 & n6942 ) ;
  assign n6944 = ( n6664 & n6666 ) | ( n6664 & ~n6676 ) | ( n6666 & ~n6676 ) ;
  assign n6945 = ( ~n6664 & n6677 ) | ( ~n6664 & n6944 ) | ( n6677 & n6944 ) ;
  assign n6946 = ( n6933 & n6943 ) | ( n6933 & ~n6945 ) | ( n6943 & ~n6945 ) ;
  assign n6947 = ( ~n6677 & n6687 ) | ( ~n6677 & n6689 ) | ( n6687 & n6689 ) ;
  assign n6948 = ( n6677 & ~n6690 ) | ( n6677 & n6947 ) | ( ~n6690 & n6947 ) ;
  assign n6949 = ~n2467 & n4200 ;
  assign n6950 = n2398 & n4215 ;
  assign n6951 = n2083 & ~n2521 ;
  assign n6952 = n6950 | n6951 ;
  assign n6953 = n6949 | n6952 ;
  assign n6954 = n4203 | n6953 ;
  assign n6955 = ( n5452 & n6953 ) | ( n5452 & n6954 ) | ( n6953 & n6954 ) ;
  assign n6956 = x26 & ~n6955 ;
  assign n6957 = ~x26 & n6955 ;
  assign n6958 = n6956 | n6957 ;
  assign n6959 = ( n6946 & n6948 ) | ( n6946 & n6958 ) | ( n6948 & n6958 ) ;
  assign n6960 = ( ~n6690 & n6700 ) | ( ~n6690 & n6702 ) | ( n6700 & n6702 ) ;
  assign n6961 = ( n6690 & ~n6703 ) | ( n6690 & n6960 ) | ( ~n6703 & n6960 ) ;
  assign n6962 = ~n2364 & n4215 ;
  assign n6963 = n2083 & ~n2467 ;
  assign n6964 = n6962 | n6963 ;
  assign n6965 = n2398 & n4200 ;
  assign n6966 = n6964 | n6965 ;
  assign n6967 = x26 & n6966 ;
  assign n6968 = n4203 & n5713 ;
  assign n6969 = x26 & ~n6968 ;
  assign n6970 = ( ~x26 & n6966 ) | ( ~x26 & n6968 ) | ( n6966 & n6968 ) ;
  assign n6971 = ( ~n6967 & n6969 ) | ( ~n6967 & n6970 ) | ( n6969 & n6970 ) ;
  assign n6972 = ( n6959 & n6961 ) | ( n6959 & n6971 ) | ( n6961 & n6971 ) ;
  assign n6973 = ( ~n6703 & n6705 ) | ( ~n6703 & n6715 ) | ( n6705 & n6715 ) ;
  assign n6974 = ( n6703 & ~n6716 ) | ( n6703 & n6973 ) | ( ~n6716 & n6973 ) ;
  assign n6975 = n2102 & n4637 ;
  assign n6976 = n2187 & n4584 ;
  assign n6977 = n6975 | n6976 ;
  assign n6978 = ~n2041 & n4649 ;
  assign n6979 = n6977 | n6978 ;
  assign n6980 = x23 & n6979 ;
  assign n6981 = n4591 & ~n4997 ;
  assign n6982 = x23 & ~n6981 ;
  assign n6983 = ( ~x23 & n6979 ) | ( ~x23 & n6981 ) | ( n6979 & n6981 ) ;
  assign n6984 = ( ~n6980 & n6982 ) | ( ~n6980 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6985 = ( n6972 & n6974 ) | ( n6972 & n6984 ) | ( n6974 & n6984 ) ;
  assign n6986 = ( ~n6716 & n6726 ) | ( ~n6716 & n6728 ) | ( n6726 & n6728 ) ;
  assign n6987 = ( n6716 & ~n6729 ) | ( n6716 & n6986 ) | ( ~n6729 & n6986 ) ;
  assign n6988 = ~n1841 & n4874 ;
  assign n6989 = n1792 & n5232 ;
  assign n6990 = n6988 | n6989 ;
  assign n6991 = n1687 & n4878 ;
  assign n6992 = n6990 | n6991 ;
  assign n6993 = n4879 | n6992 ;
  assign n6994 = ( n4331 & n6992 ) | ( n4331 & n6993 ) | ( n6992 & n6993 ) ;
  assign n6995 = x20 & ~n6994 ;
  assign n6996 = ~x20 & n6994 ;
  assign n6997 = n6995 | n6996 ;
  assign n6998 = ( n6985 & n6987 ) | ( n6985 & n6997 ) | ( n6987 & n6997 ) ;
  assign n6999 = ( n6729 & n6731 ) | ( n6729 & ~n6741 ) | ( n6731 & ~n6741 ) ;
  assign n7000 = ( ~n6729 & n6742 ) | ( ~n6729 & n6999 ) | ( n6742 & n6999 ) ;
  assign n7001 = ~n1529 & n5413 ;
  assign n7002 = n1316 & n5417 ;
  assign n7003 = n7001 | n7002 ;
  assign n7004 = n1398 & n5584 ;
  assign n7005 = n7003 | n7004 ;
  assign n7006 = n5418 | n7005 ;
  assign n7007 = ( n4084 & n7005 ) | ( n4084 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7008 = x17 & ~n7007 ;
  assign n7009 = ~x17 & n7007 ;
  assign n7010 = n7008 | n7009 ;
  assign n7011 = ( n6998 & ~n7000 ) | ( n6998 & n7010 ) | ( ~n7000 & n7010 ) ;
  assign n7012 = ( ~n6742 & n6744 ) | ( ~n6742 & n6754 ) | ( n6744 & n6754 ) ;
  assign n7013 = ( n6742 & ~n6755 ) | ( n6742 & n7012 ) | ( ~n6755 & n7012 ) ;
  assign n7014 = n1316 & n5584 ;
  assign n7015 = ~n1207 & n5417 ;
  assign n7016 = n1398 & n5413 ;
  assign n7017 = n7015 | n7016 ;
  assign n7018 = n7014 | n7017 ;
  assign n7019 = n5418 | n7018 ;
  assign n7020 = ( ~n4157 & n7018 ) | ( ~n4157 & n7019 ) | ( n7018 & n7019 ) ;
  assign n7021 = x17 & ~n7020 ;
  assign n7022 = ~x17 & n7020 ;
  assign n7023 = n7021 | n7022 ;
  assign n7024 = ( n7011 & n7013 ) | ( n7011 & n7023 ) | ( n7013 & n7023 ) ;
  assign n7025 = ( n6755 & ~n6765 ) | ( n6755 & n6767 ) | ( ~n6765 & n6767 ) ;
  assign n7026 = ( ~n6755 & n6768 ) | ( ~n6755 & n7025 ) | ( n6768 & n7025 ) ;
  assign n7027 = n995 & n5909 ;
  assign n7028 = x14 & n7027 ;
  assign n7029 = n859 & n6332 ;
  assign n7030 = ~n721 & n5914 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = n5915 | n7031 ;
  assign n7033 = ( ~n3829 & n7031 ) | ( ~n3829 & n7032 ) | ( n7031 & n7032 ) ;
  assign n7034 = x14 & ~n7033 ;
  assign n7035 = ( ~x14 & n7027 ) | ( ~x14 & n7033 ) | ( n7027 & n7033 ) ;
  assign n7036 = ( ~n7028 & n7034 ) | ( ~n7028 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7037 = ( n7024 & ~n7026 ) | ( n7024 & n7036 ) | ( ~n7026 & n7036 ) ;
  assign n7038 = ~n3487 & n6567 ;
  assign n7039 = ~n3601 & n6796 ;
  assign n7040 = n3533 & n6570 ;
  assign n7041 = ( n6570 & n7039 ) | ( n6570 & ~n7040 ) | ( n7039 & ~n7040 ) ;
  assign n7042 = n7038 | n7041 ;
  assign n7043 = n6571 | n7042 ;
  assign n7044 = ( ~n4223 & n7042 ) | ( ~n4223 & n7043 ) | ( n7042 & n7043 ) ;
  assign n7045 = x11 & ~n7044 ;
  assign n7046 = ~x11 & n7044 ;
  assign n7047 = n7045 | n7046 ;
  assign n7048 = ( ~n6768 & n6770 ) | ( ~n6768 & n6780 ) | ( n6770 & n6780 ) ;
  assign n7049 = ( n6768 & ~n6781 ) | ( n6768 & n7048 ) | ( ~n6781 & n7048 ) ;
  assign n7050 = ( n7037 & n7047 ) | ( n7037 & n7049 ) | ( n7047 & n7049 ) ;
  assign n7051 = ~n3533 & n6796 ;
  assign n7052 = x11 & n7051 ;
  assign n7053 = ~n3516 & n6570 ;
  assign n7054 = n6567 | n7053 ;
  assign n7055 = ( ~n3601 & n7053 ) | ( ~n3601 & n7054 ) | ( n7053 & n7054 ) ;
  assign n7056 = n6571 | n7055 ;
  assign n7057 = ( ~n4058 & n7055 ) | ( ~n4058 & n7056 ) | ( n7055 & n7056 ) ;
  assign n7058 = x11 & ~n7057 ;
  assign n7059 = ( ~x11 & n7051 ) | ( ~x11 & n7057 ) | ( n7051 & n7057 ) ;
  assign n7060 = ( ~n7052 & n7058 ) | ( ~n7052 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7061 = ( ~n6781 & n6791 ) | ( ~n6781 & n6793 ) | ( n6791 & n6793 ) ;
  assign n7062 = ( n6781 & ~n6794 ) | ( n6781 & n7061 ) | ( ~n6794 & n7061 ) ;
  assign n7063 = ( n7050 & n7060 ) | ( n7050 & n7062 ) | ( n7060 & n7062 ) ;
  assign n7064 = n4199 | n6841 ;
  assign n7065 = ( ~n4199 & n6838 ) | ( ~n4199 & n6841 ) | ( n6838 & n6841 ) ;
  assign n7066 = n6838 | n6841 ;
  assign n7067 = ( n7064 & n7065 ) | ( n7064 & ~n7066 ) | ( n7065 & ~n7066 ) ;
  assign n7068 = n3123 & n4584 ;
  assign n7069 = ~n2977 & n4637 ;
  assign n7070 = n7068 | n7069 ;
  assign n7071 = ~n2944 & n4649 ;
  assign n7072 = n7070 | n7071 ;
  assign n7073 = x23 & n7072 ;
  assign n7074 = n4591 & ~n5926 ;
  assign n7075 = x23 & ~n7074 ;
  assign n7076 = ( ~x23 & n7072 ) | ( ~x23 & n7074 ) | ( n7072 & n7074 ) ;
  assign n7077 = ( ~n7073 & n7075 ) | ( ~n7073 & n7076 ) | ( n7075 & n7076 ) ;
  assign n7078 = n3123 & n4637 ;
  assign n7079 = ~n2977 & n4649 ;
  assign n7080 = n7078 | n7079 ;
  assign n7081 = ~n3049 & n4584 ;
  assign n7082 = n7080 | n7081 ;
  assign n7083 = x23 & n7082 ;
  assign n7084 = n4591 & n6000 ;
  assign n7085 = x23 & ~n7084 ;
  assign n7086 = ( ~x23 & n7082 ) | ( ~x23 & n7084 ) | ( n7082 & n7084 ) ;
  assign n7087 = ( ~n7083 & n7085 ) | ( ~n7083 & n7086 ) | ( n7085 & n7086 ) ;
  assign n7088 = ~n3232 & n4590 ;
  assign n7089 = ( n3049 & n3232 ) | ( n3049 & n4587 ) | ( n3232 & n4587 ) ;
  assign n7090 = ( ~n4587 & n4590 ) | ( ~n4587 & n7089 ) | ( n4590 & n7089 ) ;
  assign n7091 = ~n3232 & n7089 ;
  assign n7092 = ( ~n3049 & n7090 ) | ( ~n3049 & n7091 ) | ( n7090 & n7091 ) ;
  assign n7093 = ~n3232 & n4637 ;
  assign n7094 = n7092 | n7093 ;
  assign n7095 = n7088 | n7094 ;
  assign n7096 = n4591 & n5965 ;
  assign n7097 = n3123 & n4649 ;
  assign n7098 = ~n3049 & n4637 ;
  assign n7099 = n7097 | n7098 ;
  assign n7100 = ~n3232 & n4584 ;
  assign n7101 = n7099 | n7100 ;
  assign n7102 = n7096 | n7101 ;
  assign n7103 = x23 & ~n7102 ;
  assign n7104 = ~n7095 & n7103 ;
  assign n7105 = ~n3232 & n4202 ;
  assign n7106 = ( n7087 & n7104 ) | ( n7087 & n7105 ) | ( n7104 & n7105 ) ;
  assign n7107 = n7087 | n7104 ;
  assign n7108 = ( ~n7087 & n7104 ) | ( ~n7087 & n7105 ) | ( n7104 & n7105 ) ;
  assign n7109 = ( ~n7106 & n7107 ) | ( ~n7106 & n7108 ) | ( n7107 & n7108 ) ;
  assign n7110 = ( n7087 & n7106 ) | ( n7087 & ~n7109 ) | ( n7106 & ~n7109 ) ;
  assign n7111 = ( n7067 & n7077 ) | ( n7067 & n7110 ) | ( n7077 & n7110 ) ;
  assign n7112 = ~n2888 & n4649 ;
  assign n7113 = ~n2977 & n4584 ;
  assign n7114 = ~n2944 & n4637 ;
  assign n7115 = n7113 | n7114 ;
  assign n7116 = n7112 | n7115 ;
  assign n7117 = n4591 | n7116 ;
  assign n7118 = ( ~n6055 & n7116 ) | ( ~n6055 & n7117 ) | ( n7116 & n7117 ) ;
  assign n7119 = x23 & ~n7118 ;
  assign n7120 = ~x23 & n7118 ;
  assign n7121 = n7119 | n7120 ;
  assign n7122 = x26 & ~n6843 ;
  assign n7123 = ~n6837 & n7122 ;
  assign n7124 = n6837 & ~n7122 ;
  assign n7125 = n7123 | n7124 ;
  assign n7126 = ( n7111 & n7121 ) | ( n7111 & n7125 ) | ( n7121 & n7125 ) ;
  assign n7127 = ~n2944 & n4584 ;
  assign n7128 = n2820 & n4649 ;
  assign n7129 = n7127 | n7128 ;
  assign n7130 = ~n2888 & n4637 ;
  assign n7131 = n7129 | n7130 ;
  assign n7132 = n4591 | n7131 ;
  assign n7133 = ( n6106 & n7131 ) | ( n6106 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7134 = x23 & ~n7133 ;
  assign n7135 = ~x23 & n7133 ;
  assign n7136 = n7134 | n7135 ;
  assign n7137 = ( n6848 & n7126 ) | ( n6848 & n7136 ) | ( n7126 & n7136 ) ;
  assign n7138 = ( ~n6817 & n6820 ) | ( ~n6817 & n6849 ) | ( n6820 & n6849 ) ;
  assign n7139 = ( n6817 & ~n6850 ) | ( n6817 & n7138 ) | ( ~n6850 & n7138 ) ;
  assign n7140 = n2735 & n4649 ;
  assign n7141 = n2820 & n4637 ;
  assign n7142 = n7140 | n7141 ;
  assign n7143 = ~n2888 & n4584 ;
  assign n7144 = n7142 | n7143 ;
  assign n7145 = n4591 | n7144 ;
  assign n7146 = ( ~n6157 & n7144 ) | ( ~n6157 & n7145 ) | ( n7144 & n7145 ) ;
  assign n7147 = x23 & ~n7146 ;
  assign n7148 = ~x23 & n7146 ;
  assign n7149 = n7147 | n7148 ;
  assign n7150 = ( n7137 & n7139 ) | ( n7137 & n7149 ) | ( n7139 & n7149 ) ;
  assign n7151 = ( ~n6850 & n6860 ) | ( ~n6850 & n6864 ) | ( n6860 & n6864 ) ;
  assign n7152 = ( n6850 & ~n6865 ) | ( n6850 & n7151 ) | ( ~n6865 & n7151 ) ;
  assign n7153 = n2820 & n4584 ;
  assign n7154 = n2642 & n4649 ;
  assign n7155 = n7153 | n7154 ;
  assign n7156 = n2735 & n4637 ;
  assign n7157 = n7155 | n7156 ;
  assign n7158 = n4591 | n7157 ;
  assign n7159 = ( n5598 & n7157 ) | ( n5598 & n7158 ) | ( n7157 & n7158 ) ;
  assign n7160 = x23 & ~n7159 ;
  assign n7161 = ~x23 & n7159 ;
  assign n7162 = n7160 | n7161 ;
  assign n7163 = ( n7150 & n7152 ) | ( n7150 & n7162 ) | ( n7152 & n7162 ) ;
  assign n7164 = ( ~n6865 & n6875 ) | ( ~n6865 & n6880 ) | ( n6875 & n6880 ) ;
  assign n7165 = ( n6865 & ~n6881 ) | ( n6865 & n7164 ) | ( ~n6881 & n7164 ) ;
  assign n7166 = n2735 & n4584 ;
  assign n7167 = n2642 & n4637 ;
  assign n7168 = ~n2608 & n4649 ;
  assign n7169 = n7167 | n7168 ;
  assign n7170 = n7166 | n7169 ;
  assign n7171 = x23 & n7170 ;
  assign n7172 = n4591 & ~n6216 ;
  assign n7173 = x23 & ~n7172 ;
  assign n7174 = ( ~x23 & n7170 ) | ( ~x23 & n7172 ) | ( n7170 & n7172 ) ;
  assign n7175 = ( ~n7171 & n7173 ) | ( ~n7171 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7176 = ( n7163 & n7165 ) | ( n7163 & n7175 ) | ( n7165 & n7175 ) ;
  assign n7177 = n2642 & n4584 ;
  assign n7178 = ~n2521 & n4649 ;
  assign n7179 = n7177 | n7178 ;
  assign n7180 = ~n2608 & n4637 ;
  assign n7181 = n7179 | n7180 ;
  assign n7182 = n4591 | n7181 ;
  assign n7183 = ( n6221 & n7181 ) | ( n6221 & n7182 ) | ( n7181 & n7182 ) ;
  assign n7184 = x23 & ~n7183 ;
  assign n7185 = ~x23 & n7183 ;
  assign n7186 = n7184 | n7185 ;
  assign n7187 = ( ~n6881 & n6891 ) | ( ~n6881 & n6893 ) | ( n6891 & n6893 ) ;
  assign n7188 = ( n6881 & ~n6894 ) | ( n6881 & n7187 ) | ( ~n6894 & n7187 ) ;
  assign n7189 = ( n7176 & n7186 ) | ( n7176 & n7188 ) | ( n7186 & n7188 ) ;
  assign n7190 = ~n2467 & n4649 ;
  assign n7191 = ~n2521 & n4637 ;
  assign n7192 = ~n2608 & n4584 ;
  assign n7193 = n7191 | n7192 ;
  assign n7194 = n7190 | n7193 ;
  assign n7195 = n4591 | n7194 ;
  assign n7196 = ( ~n5693 & n7194 ) | ( ~n5693 & n7195 ) | ( n7194 & n7195 ) ;
  assign n7197 = x23 & ~n7196 ;
  assign n7198 = ~x23 & n7196 ;
  assign n7199 = n7197 | n7198 ;
  assign n7200 = ( n6894 & n6896 ) | ( n6894 & n6906 ) | ( n6896 & n6906 ) ;
  assign n7201 = ( n6896 & n6907 ) | ( n6896 & ~n7200 ) | ( n6907 & ~n7200 ) ;
  assign n7202 = ( n7189 & n7199 ) | ( n7189 & ~n7201 ) | ( n7199 & ~n7201 ) ;
  assign n7203 = ~n2467 & n4637 ;
  assign n7204 = ~n2521 & n4584 ;
  assign n7205 = n2398 & n4649 ;
  assign n7206 = n7204 | n7205 ;
  assign n7207 = n7203 | n7206 ;
  assign n7208 = x23 & n7207 ;
  assign n7209 = n4591 & n5452 ;
  assign n7210 = x23 & ~n7209 ;
  assign n7211 = ( ~x23 & n7207 ) | ( ~x23 & n7209 ) | ( n7207 & n7209 ) ;
  assign n7212 = ( ~n7208 & n7210 ) | ( ~n7208 & n7211 ) | ( n7210 & n7211 ) ;
  assign n7213 = ( n6907 & n6909 ) | ( n6907 & ~n6919 ) | ( n6909 & ~n6919 ) ;
  assign n7214 = ( ~n6907 & n6920 ) | ( ~n6907 & n7213 ) | ( n6920 & n7213 ) ;
  assign n7215 = ( n7202 & n7212 ) | ( n7202 & ~n7214 ) | ( n7212 & ~n7214 ) ;
  assign n7216 = ( ~n6920 & n6922 ) | ( ~n6920 & n6932 ) | ( n6922 & n6932 ) ;
  assign n7217 = ( n6920 & ~n6933 ) | ( n6920 & n7216 ) | ( ~n6933 & n7216 ) ;
  assign n7218 = ~n2364 & n4649 ;
  assign n7219 = n2398 & n4637 ;
  assign n7220 = n7218 | n7219 ;
  assign n7221 = ~n2467 & n4584 ;
  assign n7222 = n7220 | n7221 ;
  assign n7223 = x23 & n7222 ;
  assign n7224 = n4591 & n5713 ;
  assign n7225 = x23 & ~n7224 ;
  assign n7226 = ( ~x23 & n7222 ) | ( ~x23 & n7224 ) | ( n7222 & n7224 ) ;
  assign n7227 = ( ~n7223 & n7225 ) | ( ~n7223 & n7226 ) | ( n7225 & n7226 ) ;
  assign n7228 = ( n7215 & n7217 ) | ( n7215 & n7227 ) | ( n7217 & n7227 ) ;
  assign n7229 = ~n2364 & n4637 ;
  assign n7230 = ~n2282 & n4649 ;
  assign n7231 = n7229 | n7230 ;
  assign n7232 = n2398 & n4584 ;
  assign n7233 = n7231 | n7232 ;
  assign n7234 = n4591 | n7233 ;
  assign n7235 = ( ~n5494 & n7233 ) | ( ~n5494 & n7234 ) | ( n7233 & n7234 ) ;
  assign n7236 = x23 & ~n7235 ;
  assign n7237 = ~x23 & n7235 ;
  assign n7238 = n7236 | n7237 ;
  assign n7239 = ( n6933 & ~n6943 ) | ( n6933 & n6945 ) | ( ~n6943 & n6945 ) ;
  assign n7240 = ( ~n6933 & n6946 ) | ( ~n6933 & n7239 ) | ( n6946 & n7239 ) ;
  assign n7241 = ( n7228 & n7238 ) | ( n7228 & ~n7240 ) | ( n7238 & ~n7240 ) ;
  assign n7242 = ( ~n6946 & n6948 ) | ( ~n6946 & n6958 ) | ( n6948 & n6958 ) ;
  assign n7243 = ( n6946 & ~n6959 ) | ( n6946 & n7242 ) | ( ~n6959 & n7242 ) ;
  assign n7244 = ~n2364 & n4584 ;
  assign n7245 = x23 & n7244 ;
  assign n7246 = n2187 & n4649 ;
  assign n7247 = ~n2282 & n4637 ;
  assign n7248 = n7246 | n7247 ;
  assign n7249 = n4591 | n7248 ;
  assign n7250 = ( n5137 & n7248 ) | ( n5137 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7251 = x23 & ~n7250 ;
  assign n7252 = ( ~x23 & n7244 ) | ( ~x23 & n7250 ) | ( n7244 & n7250 ) ;
  assign n7253 = ( ~n7245 & n7251 ) | ( ~n7245 & n7252 ) | ( n7251 & n7252 ) ;
  assign n7254 = ( n7241 & n7243 ) | ( n7241 & n7253 ) | ( n7243 & n7253 ) ;
  assign n7255 = n2102 & n4649 ;
  assign n7256 = n2187 & n4637 ;
  assign n7257 = n7255 | n7256 ;
  assign n7258 = ~n2282 & n4584 ;
  assign n7259 = n7257 | n7258 ;
  assign n7260 = n4591 | n7259 ;
  assign n7261 = ( ~n5331 & n7259 ) | ( ~n5331 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = x23 & ~n7261 ;
  assign n7263 = ~x23 & n7261 ;
  assign n7264 = n7262 | n7263 ;
  assign n7265 = ( ~n6959 & n6961 ) | ( ~n6959 & n6971 ) | ( n6961 & n6971 ) ;
  assign n7266 = ( n6959 & ~n6972 ) | ( n6959 & n7265 ) | ( ~n6972 & n7265 ) ;
  assign n7267 = ( n7254 & n7264 ) | ( n7254 & n7266 ) | ( n7264 & n7266 ) ;
  assign n7268 = ( ~n6972 & n6974 ) | ( ~n6972 & n6984 ) | ( n6974 & n6984 ) ;
  assign n7269 = ( n6972 & ~n6985 ) | ( n6972 & n7268 ) | ( ~n6985 & n7268 ) ;
  assign n7270 = ~n1841 & n5232 ;
  assign n7271 = n1943 & n4874 ;
  assign n7272 = n7270 | n7271 ;
  assign n7273 = n1792 & n4878 ;
  assign n7274 = n7272 | n7273 ;
  assign n7275 = n4879 | n7274 ;
  assign n7276 = ( ~n4831 & n7274 ) | ( ~n4831 & n7275 ) | ( n7274 & n7275 ) ;
  assign n7277 = x20 & ~n7276 ;
  assign n7278 = ~x20 & n7276 ;
  assign n7279 = n7277 | n7278 ;
  assign n7280 = ( n7267 & n7269 ) | ( n7267 & n7279 ) | ( n7269 & n7279 ) ;
  assign n7281 = ( ~n6985 & n6987 ) | ( ~n6985 & n6997 ) | ( n6987 & n6997 ) ;
  assign n7282 = ( n6985 & ~n6998 ) | ( n6985 & n7281 ) | ( ~n6998 & n7281 ) ;
  assign n7283 = n1398 & n5417 ;
  assign n7284 = n5584 | n7283 ;
  assign n7285 = ( ~n1529 & n7283 ) | ( ~n1529 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = n1600 & n5413 ;
  assign n7287 = n7285 | n7286 ;
  assign n7288 = n5418 | n7287 ;
  assign n7289 = ( ~n4324 & n7287 ) | ( ~n4324 & n7288 ) | ( n7287 & n7288 ) ;
  assign n7290 = x17 & ~n7289 ;
  assign n7291 = ~x17 & n7289 ;
  assign n7292 = n7290 | n7291 ;
  assign n7293 = ( n7280 & n7282 ) | ( n7280 & n7292 ) | ( n7282 & n7292 ) ;
  assign n7294 = ( n6998 & n7000 ) | ( n6998 & ~n7010 ) | ( n7000 & ~n7010 ) ;
  assign n7295 = ( ~n6998 & n7011 ) | ( ~n6998 & n7294 ) | ( n7011 & n7294 ) ;
  assign n7296 = n995 & n5914 ;
  assign n7297 = ~n1207 & n5909 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = ~n1118 & n6332 ;
  assign n7300 = n7298 | n7299 ;
  assign n7301 = n5915 | n7300 ;
  assign n7302 = ( n4173 & n7300 ) | ( n4173 & n7301 ) | ( n7300 & n7301 ) ;
  assign n7303 = x14 & ~n7302 ;
  assign n7304 = ~x14 & n7302 ;
  assign n7305 = n7303 | n7304 ;
  assign n7306 = ( n7293 & ~n7295 ) | ( n7293 & n7305 ) | ( ~n7295 & n7305 ) ;
  assign n7307 = ( ~n7011 & n7013 ) | ( ~n7011 & n7023 ) | ( n7013 & n7023 ) ;
  assign n7308 = ( n7011 & ~n7024 ) | ( n7011 & n7307 ) | ( ~n7024 & n7307 ) ;
  assign n7309 = n859 & n5914 ;
  assign n7310 = n995 & n6332 ;
  assign n7311 = n7309 | n7310 ;
  assign n7312 = ~n1118 & n5909 ;
  assign n7313 = n7311 | n7312 ;
  assign n7314 = n5915 | n7313 ;
  assign n7315 = ( ~n4034 & n7313 ) | ( ~n4034 & n7314 ) | ( n7313 & n7314 ) ;
  assign n7316 = x14 & ~n7315 ;
  assign n7317 = ~x14 & n7315 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = ( n7306 & n7308 ) | ( n7306 & n7318 ) | ( n7308 & n7318 ) ;
  assign n7320 = ( n7024 & n7026 ) | ( n7024 & ~n7036 ) | ( n7026 & ~n7036 ) ;
  assign n7321 = ( ~n7024 & n7037 ) | ( ~n7024 & n7320 ) | ( n7037 & n7320 ) ;
  assign n7322 = ~n3601 & n6570 ;
  assign n7323 = n564 & n6567 ;
  assign n7324 = n7322 | n7323 ;
  assign n7325 = ~n3487 & n6796 ;
  assign n7326 = n7324 | n7325 ;
  assign n7327 = n6571 | n7326 ;
  assign n7328 = ( n3674 & n7326 ) | ( n3674 & n7327 ) | ( n7326 & n7327 ) ;
  assign n7329 = x11 & ~n7328 ;
  assign n7330 = ~x11 & n7328 ;
  assign n7331 = n7329 | n7330 ;
  assign n7332 = ( n7319 & ~n7321 ) | ( n7319 & n7331 ) | ( ~n7321 & n7331 ) ;
  assign n7333 = ( ~n7037 & n7047 ) | ( ~n7037 & n7049 ) | ( n7047 & n7049 ) ;
  assign n7334 = ( n7037 & ~n7050 ) | ( n7037 & n7333 ) | ( ~n7050 & n7333 ) ;
  assign n7335 = x5 | x6 ;
  assign n7336 = x7 | n7335 ;
  assign n7337 = x8 & ~n7336 ;
  assign n7338 = x5 & x6 ;
  assign n7339 = x7 & ~x8 ;
  assign n7340 = n7338 & n7339 ;
  assign n7341 = n7337 | n7340 ;
  assign n7342 = n7335 & ~n7338 ;
  assign n7343 = x7 & x8 ;
  assign n7344 = x7 | x8 ;
  assign n7345 = ( n7342 & n7343 ) | ( n7342 & ~n7344 ) | ( n7343 & ~n7344 ) ;
  assign n7346 = n7342 & ~n7345 ;
  assign n7347 = ( ~n3516 & n3608 ) | ( ~n3516 & n7346 ) | ( n3608 & n7346 ) ;
  assign n7348 = ( ~n3607 & n7341 ) | ( ~n3607 & n7347 ) | ( n7341 & n7347 ) ;
  assign n7349 = x8 & ~n7348 ;
  assign n7350 = ~x8 & n7348 ;
  assign n7351 = n7349 | n7350 ;
  assign n7352 = ( n7332 & n7334 ) | ( n7332 & n7351 ) | ( n7334 & n7351 ) ;
  assign n7353 = n3123 & n5232 ;
  assign n7354 = ~n2977 & n4878 ;
  assign n7355 = n7353 | n7354 ;
  assign n7356 = ~n3049 & n4874 ;
  assign n7357 = n7355 | n7356 ;
  assign n7358 = x20 & n7357 ;
  assign n7359 = n4879 & n6000 ;
  assign n7360 = x20 & ~n7359 ;
  assign n7361 = ( ~x20 & n7357 ) | ( ~x20 & n7359 ) | ( n7357 & n7359 ) ;
  assign n7362 = ( ~n7358 & n7360 ) | ( ~n7358 & n7361 ) | ( n7360 & n7361 ) ;
  assign n7363 = n3233 & n4875 ;
  assign n7364 = n4879 | n5232 ;
  assign n7365 = ( n3049 & n5232 ) | ( n3049 & n7364 ) | ( n5232 & n7364 ) ;
  assign n7366 = ~n3232 & n7365 ;
  assign n7367 = n3049 | n4878 ;
  assign n7368 = ( ~n3049 & n7366 ) | ( ~n3049 & n7367 ) | ( n7366 & n7367 ) ;
  assign n7369 = n7363 | n7368 ;
  assign n7370 = ~n3232 & n4875 ;
  assign n7371 = x20 & ~n7370 ;
  assign n7372 = ~n7369 & n7371 ;
  assign n7373 = n4879 & n5965 ;
  assign n7374 = n3123 & n4878 ;
  assign n7375 = ~n3049 & n5232 ;
  assign n7376 = n7374 | n7375 ;
  assign n7377 = ~n3232 & n4874 ;
  assign n7378 = n7376 | n7377 ;
  assign n7379 = n7373 | n7378 ;
  assign n7380 = n7372 & ~n7379 ;
  assign n7381 = n7088 | n7380 ;
  assign n7382 = n7362 & n7381 ;
  assign n7383 = ~n2977 & n5232 ;
  assign n7384 = x20 & n7383 ;
  assign n7385 = ~n2944 & n4878 ;
  assign n7386 = n3123 & n4874 ;
  assign n7387 = n7385 | n7386 ;
  assign n7388 = n4879 | n7387 ;
  assign n7389 = ( ~n5926 & n7387 ) | ( ~n5926 & n7388 ) | ( n7387 & n7388 ) ;
  assign n7390 = x20 & ~n7389 ;
  assign n7391 = ( ~x20 & n7383 ) | ( ~x20 & n7389 ) | ( n7383 & n7389 ) ;
  assign n7392 = ( ~n7384 & n7390 ) | ( ~n7384 & n7391 ) | ( n7390 & n7391 ) ;
  assign n7393 = ( ~x23 & n3232 ) | ( ~x23 & n7094 ) | ( n3232 & n7094 ) ;
  assign n7394 = x23 & ~n7092 ;
  assign n7395 = ( n7095 & n7393 ) | ( n7095 & n7394 ) | ( n7393 & n7394 ) ;
  assign n7396 = ( n7382 & n7392 ) | ( n7382 & n7395 ) | ( n7392 & n7395 ) ;
  assign n7397 = ~n2888 & n4878 ;
  assign n7398 = ~n2977 & n4874 ;
  assign n7399 = ~n2944 & n5232 ;
  assign n7400 = n7398 | n7399 ;
  assign n7401 = n7397 | n7400 ;
  assign n7402 = x20 & n7401 ;
  assign n7403 = n4879 & ~n6055 ;
  assign n7404 = x20 & ~n7403 ;
  assign n7405 = ( ~x20 & n7401 ) | ( ~x20 & n7403 ) | ( n7401 & n7403 ) ;
  assign n7406 = ( ~n7402 & n7404 ) | ( ~n7402 & n7405 ) | ( n7404 & n7405 ) ;
  assign n7407 = ( x23 & n7102 ) | ( x23 & n7104 ) | ( n7102 & n7104 ) ;
  assign n7408 = ( x23 & ~n7095 ) | ( x23 & n7103 ) | ( ~n7095 & n7103 ) ;
  assign n7409 = ( n7102 & ~n7407 ) | ( n7102 & n7408 ) | ( ~n7407 & n7408 ) ;
  assign n7410 = ( n7396 & n7406 ) | ( n7396 & n7409 ) | ( n7406 & n7409 ) ;
  assign n7411 = ~n2888 & n5232 ;
  assign n7412 = ~n2944 & n4874 ;
  assign n7413 = n2820 & n4878 ;
  assign n7414 = n7412 | n7413 ;
  assign n7415 = n7411 | n7414 ;
  assign n7416 = x20 & n7415 ;
  assign n7417 = n4879 & n6106 ;
  assign n7418 = x20 & ~n7417 ;
  assign n7419 = ( ~x20 & n7415 ) | ( ~x20 & n7417 ) | ( n7415 & n7417 ) ;
  assign n7420 = ( ~n7416 & n7418 ) | ( ~n7416 & n7419 ) | ( n7418 & n7419 ) ;
  assign n7421 = ( n7109 & n7410 ) | ( n7109 & n7420 ) | ( n7410 & n7420 ) ;
  assign n7422 = n2735 & n4878 ;
  assign n7423 = n2820 & n5232 ;
  assign n7424 = n7422 | n7423 ;
  assign n7425 = ~n2888 & n4874 ;
  assign n7426 = n7424 | n7425 ;
  assign n7427 = n4879 | n7426 ;
  assign n7428 = ( ~n6157 & n7426 ) | ( ~n6157 & n7427 ) | ( n7426 & n7427 ) ;
  assign n7429 = x20 & ~n7428 ;
  assign n7430 = ~x20 & n7428 ;
  assign n7431 = n7429 | n7430 ;
  assign n7432 = ( n7067 & n7077 ) | ( n7067 & ~n7110 ) | ( n7077 & ~n7110 ) ;
  assign n7433 = ( n7110 & ~n7111 ) | ( n7110 & n7432 ) | ( ~n7111 & n7432 ) ;
  assign n7434 = ( n7421 & n7431 ) | ( n7421 & n7433 ) | ( n7431 & n7433 ) ;
  assign n7435 = ( ~n7111 & n7121 ) | ( ~n7111 & n7125 ) | ( n7121 & n7125 ) ;
  assign n7436 = ( n7111 & ~n7126 ) | ( n7111 & n7435 ) | ( ~n7126 & n7435 ) ;
  assign n7437 = n2735 & n5232 ;
  assign n7438 = n2642 & n4878 ;
  assign n7439 = n7437 | n7438 ;
  assign n7440 = n2820 & n4874 ;
  assign n7441 = n7439 | n7440 ;
  assign n7442 = n4879 | n7441 ;
  assign n7443 = ( n5598 & n7441 ) | ( n5598 & n7442 ) | ( n7441 & n7442 ) ;
  assign n7444 = x20 & ~n7443 ;
  assign n7445 = ~x20 & n7443 ;
  assign n7446 = n7444 | n7445 ;
  assign n7447 = ( n7434 & n7436 ) | ( n7434 & n7446 ) | ( n7436 & n7446 ) ;
  assign n7448 = ( n6848 & ~n7126 ) | ( n6848 & n7136 ) | ( ~n7126 & n7136 ) ;
  assign n7449 = ( n7126 & ~n7137 ) | ( n7126 & n7448 ) | ( ~n7137 & n7448 ) ;
  assign n7450 = n2735 & n4874 ;
  assign n7451 = ~n2608 & n4878 ;
  assign n7452 = n2642 & n5232 ;
  assign n7453 = n7451 | n7452 ;
  assign n7454 = n7450 | n7453 ;
  assign n7455 = x20 & n7454 ;
  assign n7456 = n4879 & ~n6216 ;
  assign n7457 = x20 & ~n7456 ;
  assign n7458 = ( ~x20 & n7454 ) | ( ~x20 & n7456 ) | ( n7454 & n7456 ) ;
  assign n7459 = ( ~n7455 & n7457 ) | ( ~n7455 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7460 = ( n7447 & n7449 ) | ( n7447 & n7459 ) | ( n7449 & n7459 ) ;
  assign n7461 = ( ~n7137 & n7139 ) | ( ~n7137 & n7149 ) | ( n7139 & n7149 ) ;
  assign n7462 = ( n7137 & ~n7150 ) | ( n7137 & n7461 ) | ( ~n7150 & n7461 ) ;
  assign n7463 = n2642 & n4874 ;
  assign n7464 = ~n2521 & n4878 ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = ~n2608 & n5232 ;
  assign n7467 = n7465 | n7466 ;
  assign n7468 = x20 & n7467 ;
  assign n7469 = n4879 & n6221 ;
  assign n7470 = x20 & ~n7469 ;
  assign n7471 = ( ~x20 & n7467 ) | ( ~x20 & n7469 ) | ( n7467 & n7469 ) ;
  assign n7472 = ( ~n7468 & n7470 ) | ( ~n7468 & n7471 ) | ( n7470 & n7471 ) ;
  assign n7473 = ( n7460 & n7462 ) | ( n7460 & n7472 ) | ( n7462 & n7472 ) ;
  assign n7474 = ( ~n7150 & n7152 ) | ( ~n7150 & n7162 ) | ( n7152 & n7162 ) ;
  assign n7475 = ( n7150 & ~n7163 ) | ( n7150 & n7474 ) | ( ~n7163 & n7474 ) ;
  assign n7476 = ~n2467 & n4878 ;
  assign n7477 = ~n2521 & n5232 ;
  assign n7478 = ~n2608 & n4874 ;
  assign n7479 = n7477 | n7478 ;
  assign n7480 = n7476 | n7479 ;
  assign n7481 = n4879 | n7480 ;
  assign n7482 = ( ~n5693 & n7480 ) | ( ~n5693 & n7481 ) | ( n7480 & n7481 ) ;
  assign n7483 = x20 & ~n7482 ;
  assign n7484 = ~x20 & n7482 ;
  assign n7485 = n7483 | n7484 ;
  assign n7486 = ( n7473 & n7475 ) | ( n7473 & n7485 ) | ( n7475 & n7485 ) ;
  assign n7487 = ( ~n7163 & n7165 ) | ( ~n7163 & n7175 ) | ( n7165 & n7175 ) ;
  assign n7488 = ( n7163 & ~n7176 ) | ( n7163 & n7487 ) | ( ~n7176 & n7487 ) ;
  assign n7489 = ~n2467 & n5232 ;
  assign n7490 = n2398 & n4878 ;
  assign n7491 = ~n2521 & n4874 ;
  assign n7492 = n7490 | n7491 ;
  assign n7493 = n7489 | n7492 ;
  assign n7494 = n4879 | n7493 ;
  assign n7495 = ( n5452 & n7493 ) | ( n5452 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7496 = x20 & ~n7495 ;
  assign n7497 = ~x20 & n7495 ;
  assign n7498 = n7496 | n7497 ;
  assign n7499 = ( n7486 & n7488 ) | ( n7486 & n7498 ) | ( n7488 & n7498 ) ;
  assign n7500 = ( ~n7176 & n7186 ) | ( ~n7176 & n7188 ) | ( n7186 & n7188 ) ;
  assign n7501 = ( n7176 & ~n7189 ) | ( n7176 & n7500 ) | ( ~n7189 & n7500 ) ;
  assign n7502 = ~n2467 & n4874 ;
  assign n7503 = ~n2364 & n4878 ;
  assign n7504 = n7502 | n7503 ;
  assign n7505 = n2398 & n5232 ;
  assign n7506 = n7504 | n7505 ;
  assign n7507 = x20 & n7506 ;
  assign n7508 = n4879 & n5713 ;
  assign n7509 = x20 & ~n7508 ;
  assign n7510 = ( ~x20 & n7506 ) | ( ~x20 & n7508 ) | ( n7506 & n7508 ) ;
  assign n7511 = ( ~n7507 & n7509 ) | ( ~n7507 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = ( n7499 & n7501 ) | ( n7499 & n7511 ) | ( n7501 & n7511 ) ;
  assign n7513 = ~n2364 & n5232 ;
  assign n7514 = n2398 & n4874 ;
  assign n7515 = n7513 | n7514 ;
  assign n7516 = ~n2282 & n4878 ;
  assign n7517 = n7515 | n7516 ;
  assign n7518 = x20 & n7517 ;
  assign n7519 = n4879 & ~n5494 ;
  assign n7520 = x20 & ~n7519 ;
  assign n7521 = ( ~x20 & n7517 ) | ( ~x20 & n7519 ) | ( n7517 & n7519 ) ;
  assign n7522 = ( ~n7518 & n7520 ) | ( ~n7518 & n7521 ) | ( n7520 & n7521 ) ;
  assign n7523 = ( n7189 & ~n7199 ) | ( n7189 & n7201 ) | ( ~n7199 & n7201 ) ;
  assign n7524 = ( ~n7189 & n7202 ) | ( ~n7189 & n7523 ) | ( n7202 & n7523 ) ;
  assign n7525 = ( n7512 & n7522 ) | ( n7512 & ~n7524 ) | ( n7522 & ~n7524 ) ;
  assign n7526 = ( n7202 & ~n7212 ) | ( n7202 & n7214 ) | ( ~n7212 & n7214 ) ;
  assign n7527 = ( ~n7202 & n7215 ) | ( ~n7202 & n7526 ) | ( n7215 & n7526 ) ;
  assign n7528 = ~n2364 & n4874 ;
  assign n7529 = x20 & n7528 ;
  assign n7530 = n2187 & n4878 ;
  assign n7531 = ~n2282 & n5232 ;
  assign n7532 = n7530 | n7531 ;
  assign n7533 = n4879 | n7532 ;
  assign n7534 = ( n5137 & n7532 ) | ( n5137 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = x20 & ~n7534 ;
  assign n7536 = ( ~x20 & n7528 ) | ( ~x20 & n7534 ) | ( n7528 & n7534 ) ;
  assign n7537 = ( ~n7529 & n7535 ) | ( ~n7529 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7538 = ( n7525 & ~n7527 ) | ( n7525 & n7537 ) | ( ~n7527 & n7537 ) ;
  assign n7539 = ( ~n7215 & n7217 ) | ( ~n7215 & n7227 ) | ( n7217 & n7227 ) ;
  assign n7540 = ( n7215 & ~n7228 ) | ( n7215 & n7539 ) | ( ~n7228 & n7539 ) ;
  assign n7541 = n2102 & n4878 ;
  assign n7542 = n2187 & n5232 ;
  assign n7543 = n7541 | n7542 ;
  assign n7544 = ~n2282 & n4874 ;
  assign n7545 = n7543 | n7544 ;
  assign n7546 = x20 & n7545 ;
  assign n7547 = n4879 & ~n5331 ;
  assign n7548 = x20 & ~n7547 ;
  assign n7549 = ( ~x20 & n7545 ) | ( ~x20 & n7547 ) | ( n7545 & n7547 ) ;
  assign n7550 = ( ~n7546 & n7548 ) | ( ~n7546 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7551 = ( n7538 & n7540 ) | ( n7538 & n7550 ) | ( n7540 & n7550 ) ;
  assign n7552 = ~n2041 & n4878 ;
  assign n7553 = n2102 & n5232 ;
  assign n7554 = n7552 | n7553 ;
  assign n7555 = n2187 & n4874 ;
  assign n7556 = n7554 | n7555 ;
  assign n7557 = n4879 | n7556 ;
  assign n7558 = ( ~n4997 & n7556 ) | ( ~n4997 & n7557 ) | ( n7556 & n7557 ) ;
  assign n7559 = x20 & ~n7558 ;
  assign n7560 = ~x20 & n7558 ;
  assign n7561 = n7559 | n7560 ;
  assign n7562 = ( n7228 & n7238 ) | ( n7228 & n7240 ) | ( n7238 & n7240 ) ;
  assign n7563 = ( n7240 & n7241 ) | ( n7240 & ~n7562 ) | ( n7241 & ~n7562 ) ;
  assign n7564 = ( n7551 & n7561 ) | ( n7551 & ~n7563 ) | ( n7561 & ~n7563 ) ;
  assign n7565 = ( ~n7241 & n7243 ) | ( ~n7241 & n7253 ) | ( n7243 & n7253 ) ;
  assign n7566 = ( n7241 & ~n7254 ) | ( n7241 & n7565 ) | ( ~n7254 & n7565 ) ;
  assign n7567 = ~n2041 & n5232 ;
  assign n7568 = x20 & n7567 ;
  assign n7569 = n1943 & n4878 ;
  assign n7570 = n2102 & n4874 ;
  assign n7571 = n7569 | n7570 ;
  assign n7572 = n4879 | n7571 ;
  assign n7573 = ( ~n4985 & n7571 ) | ( ~n4985 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = x20 & ~n7573 ;
  assign n7575 = ( ~x20 & n7567 ) | ( ~x20 & n7573 ) | ( n7567 & n7573 ) ;
  assign n7576 = ( ~n7568 & n7574 ) | ( ~n7568 & n7575 ) | ( n7574 & n7575 ) ;
  assign n7577 = ( n7564 & n7566 ) | ( n7564 & n7576 ) | ( n7566 & n7576 ) ;
  assign n7578 = ( ~n7254 & n7264 ) | ( ~n7254 & n7266 ) | ( n7264 & n7266 ) ;
  assign n7579 = ( n7254 & ~n7267 ) | ( n7254 & n7578 ) | ( ~n7267 & n7578 ) ;
  assign n7580 = ~n1841 & n4878 ;
  assign n7581 = n1943 & n5232 ;
  assign n7582 = n7580 | n7581 ;
  assign n7583 = ~n2041 & n4874 ;
  assign n7584 = n7582 | n7583 ;
  assign n7585 = n4879 | n7584 ;
  assign n7586 = ( ~n4753 & n7584 ) | ( ~n4753 & n7585 ) | ( n7584 & n7585 ) ;
  assign n7587 = x20 & ~n7586 ;
  assign n7588 = ~x20 & n7586 ;
  assign n7589 = n7587 | n7588 ;
  assign n7590 = ( n7577 & n7579 ) | ( n7577 & n7589 ) | ( n7579 & n7589 ) ;
  assign n7591 = ( ~n7267 & n7269 ) | ( ~n7267 & n7279 ) | ( n7269 & n7279 ) ;
  assign n7592 = ( n7267 & ~n7280 ) | ( n7267 & n7591 ) | ( ~n7280 & n7591 ) ;
  assign n7593 = ~n1529 & n5417 ;
  assign n7594 = n1687 & n5413 ;
  assign n7595 = n7593 | n7594 ;
  assign n7596 = n1600 & n5584 ;
  assign n7597 = n7595 | n7596 ;
  assign n7598 = n5418 | n7597 ;
  assign n7599 = ( ~n4531 & n7597 ) | ( ~n4531 & n7598 ) | ( n7597 & n7598 ) ;
  assign n7600 = x17 & ~n7599 ;
  assign n7601 = ~x17 & n7599 ;
  assign n7602 = n7600 | n7601 ;
  assign n7603 = ( n7590 & n7592 ) | ( n7590 & n7602 ) | ( n7592 & n7602 ) ;
  assign n7604 = ( ~n7280 & n7282 ) | ( ~n7280 & n7292 ) | ( n7282 & n7292 ) ;
  assign n7605 = ( n7280 & ~n7293 ) | ( n7280 & n7604 ) | ( ~n7293 & n7604 ) ;
  assign n7606 = n1316 & n5909 ;
  assign n7607 = ~n1207 & n6332 ;
  assign n7608 = n7606 | n7607 ;
  assign n7609 = ~n1118 & n5914 ;
  assign n7610 = n7608 | n7609 ;
  assign n7611 = n5915 | n7610 ;
  assign n7612 = ( n3841 & n7610 ) | ( n3841 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = x14 & ~n7612 ;
  assign n7614 = ~x14 & n7612 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = ( n7603 & n7605 ) | ( n7603 & n7615 ) | ( n7605 & n7615 ) ;
  assign n7617 = ( n7293 & n7295 ) | ( n7293 & ~n7305 ) | ( n7295 & ~n7305 ) ;
  assign n7618 = ( ~n7293 & n7306 ) | ( ~n7293 & n7617 ) | ( n7306 & n7617 ) ;
  assign n7619 = ~n721 & n6796 ;
  assign n7620 = x11 & n7619 ;
  assign n7621 = n859 & n6567 ;
  assign n7622 = n564 & n6570 ;
  assign n7623 = n7621 | n7622 ;
  assign n7624 = n6571 | n7623 ;
  assign n7625 = ( ~n3268 & n7623 ) | ( ~n3268 & n7624 ) | ( n7623 & n7624 ) ;
  assign n7626 = x11 & ~n7625 ;
  assign n7627 = ( ~x11 & n7619 ) | ( ~x11 & n7625 ) | ( n7619 & n7625 ) ;
  assign n7628 = ( ~n7620 & n7626 ) | ( ~n7620 & n7627 ) | ( n7626 & n7627 ) ;
  assign n7629 = ( n7616 & ~n7618 ) | ( n7616 & n7628 ) | ( ~n7618 & n7628 ) ;
  assign n7630 = ( ~n7306 & n7308 ) | ( ~n7306 & n7318 ) | ( n7308 & n7318 ) ;
  assign n7631 = ( n7306 & ~n7319 ) | ( n7306 & n7630 ) | ( ~n7319 & n7630 ) ;
  assign n7632 = ~n3487 & n6570 ;
  assign n7633 = ~n721 & n6567 ;
  assign n7634 = n564 & n6796 ;
  assign n7635 = n7633 | n7634 ;
  assign n7636 = n7632 | n7635 ;
  assign n7637 = n6571 | n7636 ;
  assign n7638 = ( ~n3492 & n7636 ) | ( ~n3492 & n7637 ) | ( n7636 & n7637 ) ;
  assign n7639 = x11 & ~n7638 ;
  assign n7640 = ~x11 & n7638 ;
  assign n7641 = n7639 | n7640 ;
  assign n7642 = ( n7629 & n7631 ) | ( n7629 & n7641 ) | ( n7631 & n7641 ) ;
  assign n7643 = ( x7 & n7335 ) | ( x7 & n7342 ) | ( n7335 & n7342 ) ;
  assign n7644 = n7336 & ~n7643 ;
  assign n7645 = ~n3516 & n7644 ;
  assign n7646 = x8 & n7645 ;
  assign n7647 = ~n3533 & n7341 ;
  assign n7648 = n7346 | n7647 ;
  assign n7649 = ( n3609 & n7647 ) | ( n3609 & n7648 ) | ( n7647 & n7648 ) ;
  assign n7650 = x8 & ~n7649 ;
  assign n7651 = ( ~x8 & n7645 ) | ( ~x8 & n7649 ) | ( n7645 & n7649 ) ;
  assign n7652 = ( ~n7646 & n7650 ) | ( ~n7646 & n7651 ) | ( n7650 & n7651 ) ;
  assign n7653 = ( n7319 & n7321 ) | ( n7319 & ~n7331 ) | ( n7321 & ~n7331 ) ;
  assign n7654 = ( ~n7319 & n7332 ) | ( ~n7319 & n7653 ) | ( n7332 & n7653 ) ;
  assign n7655 = ( n7642 & n7652 ) | ( n7642 & ~n7654 ) | ( n7652 & ~n7654 ) ;
  assign n7656 = ~n2977 & n5584 ;
  assign n7657 = ~n2944 & n5417 ;
  assign n7658 = n7656 | n7657 ;
  assign n7659 = n3123 & n5413 ;
  assign n7660 = n7658 | n7659 ;
  assign n7661 = x17 & n7660 ;
  assign n7662 = n5418 & ~n5926 ;
  assign n7663 = x17 & ~n7662 ;
  assign n7664 = ( ~x17 & n7660 ) | ( ~x17 & n7662 ) | ( n7660 & n7662 ) ;
  assign n7665 = ( ~n7661 & n7663 ) | ( ~n7661 & n7664 ) | ( n7663 & n7664 ) ;
  assign n7666 = x20 & n7370 ;
  assign n7667 = ~n7369 & n7666 ;
  assign n7668 = n7369 & ~n7666 ;
  assign n7669 = n7667 | n7668 ;
  assign n7670 = ~n2977 & n5417 ;
  assign n7671 = ~n3049 & n5413 ;
  assign n7672 = n7670 | n7671 ;
  assign n7673 = n3123 & n5584 ;
  assign n7674 = n7672 | n7673 ;
  assign n7675 = x17 & n7674 ;
  assign n7676 = n5418 & n6000 ;
  assign n7677 = x17 & ~n7676 ;
  assign n7678 = ( ~x17 & n7674 ) | ( ~x17 & n7676 ) | ( n7674 & n7676 ) ;
  assign n7679 = ( ~n7675 & n7677 ) | ( ~n7675 & n7678 ) | ( n7677 & n7678 ) ;
  assign n7680 = n5418 & n5965 ;
  assign n7681 = n3123 & n5417 ;
  assign n7682 = ~n3049 & n5584 ;
  assign n7683 = n7681 | n7682 ;
  assign n7684 = ~n3232 & n5413 ;
  assign n7685 = n7683 | n7684 ;
  assign n7686 = n7680 | n7685 ;
  assign n7687 = n5418 | n5584 ;
  assign n7688 = ( n3049 & n5584 ) | ( n3049 & n7687 ) | ( n5584 & n7687 ) ;
  assign n7689 = ~n3232 & n7688 ;
  assign n7690 = n3232 | n5417 ;
  assign n7691 = ~n3049 & n5414 ;
  assign n7692 = n7690 & n7691 ;
  assign n7693 = n7689 | n7692 ;
  assign n7694 = ~n3232 & n5414 ;
  assign n7695 = x17 & ~n7694 ;
  assign n7696 = ~n7693 & n7695 ;
  assign n7697 = ~n7686 & n7696 ;
  assign n7698 = ( n7370 & n7679 ) | ( n7370 & ~n7697 ) | ( n7679 & ~n7697 ) ;
  assign n7699 = n7370 & ~n7697 ;
  assign n7700 = ( n7370 & ~n7679 ) | ( n7370 & n7697 ) | ( ~n7679 & n7697 ) ;
  assign n7701 = ( n7698 & ~n7699 ) | ( n7698 & n7700 ) | ( ~n7699 & n7700 ) ;
  assign n7702 = ( n7370 & n7679 ) | ( n7370 & ~n7701 ) | ( n7679 & ~n7701 ) ;
  assign n7703 = ( n7665 & n7669 ) | ( n7665 & n7702 ) | ( n7669 & n7702 ) ;
  assign n7704 = ~n2888 & n5417 ;
  assign n7705 = ~n2977 & n5413 ;
  assign n7706 = ~n2944 & n5584 ;
  assign n7707 = n7705 | n7706 ;
  assign n7708 = n7704 | n7707 ;
  assign n7709 = x17 & n7708 ;
  assign n7710 = n5418 & ~n6055 ;
  assign n7711 = x17 & ~n7710 ;
  assign n7712 = ( ~x17 & n7708 ) | ( ~x17 & n7710 ) | ( n7708 & n7710 ) ;
  assign n7713 = ( ~n7709 & n7711 ) | ( ~n7709 & n7712 ) | ( n7711 & n7712 ) ;
  assign n7714 = x20 & ~n7372 ;
  assign n7715 = ~n7379 & n7714 ;
  assign n7716 = n7379 & ~n7714 ;
  assign n7717 = n7715 | n7716 ;
  assign n7718 = ( n7703 & n7713 ) | ( n7703 & n7717 ) | ( n7713 & n7717 ) ;
  assign n7719 = n2820 & n5417 ;
  assign n7720 = x17 & n7719 ;
  assign n7721 = n5418 & n6106 ;
  assign n7722 = ~n2944 & n5413 ;
  assign n7723 = ~n2888 & n5584 ;
  assign n7724 = n7722 | n7723 ;
  assign n7725 = n7721 | n7724 ;
  assign n7726 = x17 & ~n7725 ;
  assign n7727 = ( ~x17 & n7719 ) | ( ~x17 & n7725 ) | ( n7719 & n7725 ) ;
  assign n7728 = ( ~n7720 & n7726 ) | ( ~n7720 & n7727 ) | ( n7726 & n7727 ) ;
  assign n7729 = ( n7088 & n7362 ) | ( n7088 & ~n7380 ) | ( n7362 & ~n7380 ) ;
  assign n7730 = ( n7380 & ~n7382 ) | ( n7380 & n7729 ) | ( ~n7382 & n7729 ) ;
  assign n7731 = ( n7718 & n7728 ) | ( n7718 & n7730 ) | ( n7728 & n7730 ) ;
  assign n7732 = ~n2888 & n5413 ;
  assign n7733 = n2735 & n5417 ;
  assign n7734 = n2820 & n5584 ;
  assign n7735 = n7733 | n7734 ;
  assign n7736 = n7732 | n7735 ;
  assign n7737 = x17 & n7736 ;
  assign n7738 = n5418 & ~n6157 ;
  assign n7739 = x17 & ~n7738 ;
  assign n7740 = ( ~x17 & n7736 ) | ( ~x17 & n7738 ) | ( n7736 & n7738 ) ;
  assign n7741 = ( ~n7737 & n7739 ) | ( ~n7737 & n7740 ) | ( n7739 & n7740 ) ;
  assign n7742 = ( n7382 & ~n7392 ) | ( n7382 & n7395 ) | ( ~n7392 & n7395 ) ;
  assign n7743 = ( n7392 & ~n7396 ) | ( n7392 & n7742 ) | ( ~n7396 & n7742 ) ;
  assign n7744 = ( n7731 & n7741 ) | ( n7731 & n7743 ) | ( n7741 & n7743 ) ;
  assign n7745 = ( ~n7396 & n7406 ) | ( ~n7396 & n7409 ) | ( n7406 & n7409 ) ;
  assign n7746 = ( n7396 & ~n7410 ) | ( n7396 & n7745 ) | ( ~n7410 & n7745 ) ;
  assign n7747 = n2820 & n5413 ;
  assign n7748 = n2642 & n5417 ;
  assign n7749 = n7747 | n7748 ;
  assign n7750 = n2735 & n5584 ;
  assign n7751 = n7749 | n7750 ;
  assign n7752 = x17 & n7751 ;
  assign n7753 = n5418 & n5598 ;
  assign n7754 = x17 & ~n7753 ;
  assign n7755 = ( ~x17 & n7751 ) | ( ~x17 & n7753 ) | ( n7751 & n7753 ) ;
  assign n7756 = ( ~n7752 & n7754 ) | ( ~n7752 & n7755 ) | ( n7754 & n7755 ) ;
  assign n7757 = ( n7744 & n7746 ) | ( n7744 & n7756 ) | ( n7746 & n7756 ) ;
  assign n7758 = ( n7109 & ~n7410 ) | ( n7109 & n7420 ) | ( ~n7410 & n7420 ) ;
  assign n7759 = ( n7410 & ~n7421 ) | ( n7410 & n7758 ) | ( ~n7421 & n7758 ) ;
  assign n7760 = n2735 & n5413 ;
  assign n7761 = n2642 & n5584 ;
  assign n7762 = ~n2608 & n5417 ;
  assign n7763 = n7761 | n7762 ;
  assign n7764 = n7760 | n7763 ;
  assign n7765 = x17 & n7764 ;
  assign n7766 = n5418 & ~n6216 ;
  assign n7767 = x17 & ~n7766 ;
  assign n7768 = ( ~x17 & n7764 ) | ( ~x17 & n7766 ) | ( n7764 & n7766 ) ;
  assign n7769 = ( ~n7765 & n7767 ) | ( ~n7765 & n7768 ) | ( n7767 & n7768 ) ;
  assign n7770 = ( n7757 & n7759 ) | ( n7757 & n7769 ) | ( n7759 & n7769 ) ;
  assign n7771 = ( ~n7421 & n7431 ) | ( ~n7421 & n7433 ) | ( n7431 & n7433 ) ;
  assign n7772 = ( n7421 & ~n7434 ) | ( n7421 & n7771 ) | ( ~n7434 & n7771 ) ;
  assign n7773 = n2642 & n5413 ;
  assign n7774 = ~n2608 & n5584 ;
  assign n7775 = n7773 | n7774 ;
  assign n7776 = ~n2521 & n5417 ;
  assign n7777 = n7775 | n7776 ;
  assign n7778 = x17 & n7777 ;
  assign n7779 = n5418 & n6221 ;
  assign n7780 = x17 & ~n7779 ;
  assign n7781 = ( ~x17 & n7777 ) | ( ~x17 & n7779 ) | ( n7777 & n7779 ) ;
  assign n7782 = ( ~n7778 & n7780 ) | ( ~n7778 & n7781 ) | ( n7780 & n7781 ) ;
  assign n7783 = ( n7770 & n7772 ) | ( n7770 & n7782 ) | ( n7772 & n7782 ) ;
  assign n7784 = ~n2467 & n5417 ;
  assign n7785 = ~n2521 & n5584 ;
  assign n7786 = ~n2608 & n5413 ;
  assign n7787 = n7785 | n7786 ;
  assign n7788 = n7784 | n7787 ;
  assign n7789 = x17 & n7788 ;
  assign n7790 = n5418 & ~n5693 ;
  assign n7791 = ( ~x17 & n7788 ) | ( ~x17 & n7790 ) | ( n7788 & n7790 ) ;
  assign n7792 = x17 & ~n7790 ;
  assign n7793 = ( ~n7789 & n7791 ) | ( ~n7789 & n7792 ) | ( n7791 & n7792 ) ;
  assign n7794 = ( ~n7434 & n7436 ) | ( ~n7434 & n7446 ) | ( n7436 & n7446 ) ;
  assign n7795 = ( n7434 & ~n7447 ) | ( n7434 & n7794 ) | ( ~n7447 & n7794 ) ;
  assign n7796 = ( n7783 & n7793 ) | ( n7783 & n7795 ) | ( n7793 & n7795 ) ;
  assign n7797 = ( ~n7447 & n7449 ) | ( ~n7447 & n7459 ) | ( n7449 & n7459 ) ;
  assign n7798 = ( n7447 & ~n7460 ) | ( n7447 & n7797 ) | ( ~n7460 & n7797 ) ;
  assign n7799 = ~n2467 & n5584 ;
  assign n7800 = ~n2521 & n5413 ;
  assign n7801 = n2398 & n5417 ;
  assign n7802 = n7800 | n7801 ;
  assign n7803 = n7799 | n7802 ;
  assign n7804 = x17 & n7803 ;
  assign n7805 = n5418 & n5452 ;
  assign n7806 = x17 & ~n7805 ;
  assign n7807 = ( ~x17 & n7803 ) | ( ~x17 & n7805 ) | ( n7803 & n7805 ) ;
  assign n7808 = ( ~n7804 & n7806 ) | ( ~n7804 & n7807 ) | ( n7806 & n7807 ) ;
  assign n7809 = ( n7796 & n7798 ) | ( n7796 & n7808 ) | ( n7798 & n7808 ) ;
  assign n7810 = ( ~n7460 & n7462 ) | ( ~n7460 & n7472 ) | ( n7462 & n7472 ) ;
  assign n7811 = ( n7460 & ~n7473 ) | ( n7460 & n7810 ) | ( ~n7473 & n7810 ) ;
  assign n7812 = ~n2467 & n5413 ;
  assign n7813 = ~n2364 & n5417 ;
  assign n7814 = n7812 | n7813 ;
  assign n7815 = n2398 & n5584 ;
  assign n7816 = n7814 | n7815 ;
  assign n7817 = x17 & n7816 ;
  assign n7818 = n5418 & n5713 ;
  assign n7819 = x17 & ~n7818 ;
  assign n7820 = ( ~x17 & n7816 ) | ( ~x17 & n7818 ) | ( n7816 & n7818 ) ;
  assign n7821 = ( ~n7817 & n7819 ) | ( ~n7817 & n7820 ) | ( n7819 & n7820 ) ;
  assign n7822 = ( n7809 & n7811 ) | ( n7809 & n7821 ) | ( n7811 & n7821 ) ;
  assign n7823 = ( ~n7473 & n7475 ) | ( ~n7473 & n7485 ) | ( n7475 & n7485 ) ;
  assign n7824 = ( n7473 & ~n7486 ) | ( n7473 & n7823 ) | ( ~n7486 & n7823 ) ;
  assign n7825 = ~n2282 & n5417 ;
  assign n7826 = ~n2364 & n5584 ;
  assign n7827 = n7825 | n7826 ;
  assign n7828 = n2398 & n5413 ;
  assign n7829 = n7827 | n7828 ;
  assign n7830 = x17 & n7829 ;
  assign n7831 = n5418 & ~n5494 ;
  assign n7832 = x17 & ~n7831 ;
  assign n7833 = ( ~x17 & n7829 ) | ( ~x17 & n7831 ) | ( n7829 & n7831 ) ;
  assign n7834 = ( ~n7830 & n7832 ) | ( ~n7830 & n7833 ) | ( n7832 & n7833 ) ;
  assign n7835 = ( n7822 & n7824 ) | ( n7822 & n7834 ) | ( n7824 & n7834 ) ;
  assign n7836 = ( ~n7486 & n7488 ) | ( ~n7486 & n7498 ) | ( n7488 & n7498 ) ;
  assign n7837 = ( n7486 & ~n7499 ) | ( n7486 & n7836 ) | ( ~n7499 & n7836 ) ;
  assign n7838 = ~n2364 & n5413 ;
  assign n7839 = n2187 & n5417 ;
  assign n7840 = n7838 | n7839 ;
  assign n7841 = ~n2282 & n5584 ;
  assign n7842 = n7840 | n7841 ;
  assign n7843 = x17 & n7842 ;
  assign n7844 = n5137 & n5418 ;
  assign n7845 = x17 & ~n7844 ;
  assign n7846 = ( ~x17 & n7842 ) | ( ~x17 & n7844 ) | ( n7842 & n7844 ) ;
  assign n7847 = ( ~n7843 & n7845 ) | ( ~n7843 & n7846 ) | ( n7845 & n7846 ) ;
  assign n7848 = ( n7835 & n7837 ) | ( n7835 & n7847 ) | ( n7837 & n7847 ) ;
  assign n7849 = ( ~n7499 & n7501 ) | ( ~n7499 & n7511 ) | ( n7501 & n7511 ) ;
  assign n7850 = ( n7499 & ~n7512 ) | ( n7499 & n7849 ) | ( ~n7512 & n7849 ) ;
  assign n7851 = n2102 & n5417 ;
  assign n7852 = n2187 & n5584 ;
  assign n7853 = n7851 | n7852 ;
  assign n7854 = ~n2282 & n5413 ;
  assign n7855 = n7853 | n7854 ;
  assign n7856 = x17 & n7855 ;
  assign n7857 = ~n5331 & n5418 ;
  assign n7858 = ( ~x17 & n7855 ) | ( ~x17 & n7857 ) | ( n7855 & n7857 ) ;
  assign n7859 = x17 & ~n7857 ;
  assign n7860 = ( ~n7856 & n7858 ) | ( ~n7856 & n7859 ) | ( n7858 & n7859 ) ;
  assign n7861 = ( n7848 & n7850 ) | ( n7848 & n7860 ) | ( n7850 & n7860 ) ;
  assign n7862 = ~n2041 & n5417 ;
  assign n7863 = n2102 & n5584 ;
  assign n7864 = n7862 | n7863 ;
  assign n7865 = n2187 & n5413 ;
  assign n7866 = n7864 | n7865 ;
  assign n7867 = n5418 | n7866 ;
  assign n7868 = ( ~n4997 & n7866 ) | ( ~n4997 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = x17 & ~n7868 ;
  assign n7870 = ~x17 & n7868 ;
  assign n7871 = n7869 | n7870 ;
  assign n7872 = ( n7512 & n7522 ) | ( n7512 & n7524 ) | ( n7522 & n7524 ) ;
  assign n7873 = ( n7524 & n7525 ) | ( n7524 & ~n7872 ) | ( n7525 & ~n7872 ) ;
  assign n7874 = ( n7861 & n7871 ) | ( n7861 & ~n7873 ) | ( n7871 & ~n7873 ) ;
  assign n7875 = ~n2041 & n5584 ;
  assign n7876 = n1943 & n5417 ;
  assign n7877 = n7875 | n7876 ;
  assign n7878 = n2102 & n5413 ;
  assign n7879 = n7877 | n7878 ;
  assign n7880 = n5418 | n7879 ;
  assign n7881 = ( ~n4985 & n7879 ) | ( ~n4985 & n7880 ) | ( n7879 & n7880 ) ;
  assign n7882 = x17 & ~n7881 ;
  assign n7883 = ~x17 & n7881 ;
  assign n7884 = n7882 | n7883 ;
  assign n7885 = ( n7525 & n7527 ) | ( n7525 & n7537 ) | ( n7527 & n7537 ) ;
  assign n7886 = ( n7527 & n7538 ) | ( n7527 & ~n7885 ) | ( n7538 & ~n7885 ) ;
  assign n7887 = ( n7874 & n7884 ) | ( n7874 & ~n7886 ) | ( n7884 & ~n7886 ) ;
  assign n7888 = ~n2041 & n5413 ;
  assign n7889 = n1943 & n5584 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = ~n1841 & n5417 ;
  assign n7892 = n7890 | n7891 ;
  assign n7893 = n5418 | n7892 ;
  assign n7894 = ( ~n4753 & n7892 ) | ( ~n4753 & n7893 ) | ( n7892 & n7893 ) ;
  assign n7895 = x17 & ~n7894 ;
  assign n7896 = ~x17 & n7894 ;
  assign n7897 = n7895 | n7896 ;
  assign n7898 = ( ~n7538 & n7540 ) | ( ~n7538 & n7550 ) | ( n7540 & n7550 ) ;
  assign n7899 = ( n7538 & ~n7551 ) | ( n7538 & n7898 ) | ( ~n7551 & n7898 ) ;
  assign n7900 = ( n7887 & n7897 ) | ( n7887 & n7899 ) | ( n7897 & n7899 ) ;
  assign n7901 = n1943 & n5413 ;
  assign n7902 = ~n1841 & n5584 ;
  assign n7903 = n7901 | n7902 ;
  assign n7904 = n1792 & n5417 ;
  assign n7905 = n7903 | n7904 ;
  assign n7906 = n5418 | n7905 ;
  assign n7907 = ( ~n4831 & n7905 ) | ( ~n4831 & n7906 ) | ( n7905 & n7906 ) ;
  assign n7908 = x17 & ~n7907 ;
  assign n7909 = ~x17 & n7907 ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = ( n7551 & ~n7561 ) | ( n7551 & n7563 ) | ( ~n7561 & n7563 ) ;
  assign n7912 = ( ~n7551 & n7564 ) | ( ~n7551 & n7911 ) | ( n7564 & n7911 ) ;
  assign n7913 = ( n7900 & n7910 ) | ( n7900 & ~n7912 ) | ( n7910 & ~n7912 ) ;
  assign n7914 = ~n1841 & n5413 ;
  assign n7915 = n1792 & n5584 ;
  assign n7916 = n7914 | n7915 ;
  assign n7917 = n1687 & n5417 ;
  assign n7918 = n7916 | n7917 ;
  assign n7919 = n5418 | n7918 ;
  assign n7920 = ( n4331 & n7918 ) | ( n4331 & n7919 ) | ( n7918 & n7919 ) ;
  assign n7921 = x17 & ~n7920 ;
  assign n7922 = ~x17 & n7920 ;
  assign n7923 = n7921 | n7922 ;
  assign n7924 = ( ~n7564 & n7566 ) | ( ~n7564 & n7576 ) | ( n7566 & n7576 ) ;
  assign n7925 = ( n7564 & ~n7577 ) | ( n7564 & n7924 ) | ( ~n7577 & n7924 ) ;
  assign n7926 = ( n7913 & n7923 ) | ( n7913 & n7925 ) | ( n7923 & n7925 ) ;
  assign n7927 = ( ~n7577 & n7579 ) | ( ~n7577 & n7589 ) | ( n7579 & n7589 ) ;
  assign n7928 = ( n7577 & ~n7590 ) | ( n7577 & n7927 ) | ( ~n7590 & n7927 ) ;
  assign n7929 = n1687 & n5584 ;
  assign n7930 = n1792 & n5413 ;
  assign n7931 = n1600 & n5417 ;
  assign n7932 = n7930 | n7931 ;
  assign n7933 = n7929 | n7932 ;
  assign n7934 = n5418 | n7933 ;
  assign n7935 = ( n4674 & n7933 ) | ( n4674 & n7934 ) | ( n7933 & n7934 ) ;
  assign n7936 = x17 & ~n7935 ;
  assign n7937 = ~x17 & n7935 ;
  assign n7938 = n7936 | n7937 ;
  assign n7939 = ( n7926 & n7928 ) | ( n7926 & n7938 ) | ( n7928 & n7938 ) ;
  assign n7940 = ( ~n7590 & n7592 ) | ( ~n7590 & n7602 ) | ( n7592 & n7602 ) ;
  assign n7941 = ( n7590 & ~n7603 ) | ( n7590 & n7940 ) | ( ~n7603 & n7940 ) ;
  assign n7942 = n1316 & n6332 ;
  assign n7943 = ~n1207 & n5914 ;
  assign n7944 = n1398 & n5909 ;
  assign n7945 = n7943 | n7944 ;
  assign n7946 = n7942 | n7945 ;
  assign n7947 = n5915 | n7946 ;
  assign n7948 = ( ~n4157 & n7946 ) | ( ~n4157 & n7947 ) | ( n7946 & n7947 ) ;
  assign n7949 = x14 & ~n7948 ;
  assign n7950 = ~x14 & n7948 ;
  assign n7951 = n7949 | n7950 ;
  assign n7952 = ( n7939 & n7941 ) | ( n7939 & n7951 ) | ( n7941 & n7951 ) ;
  assign n7953 = n859 & n6796 ;
  assign n7954 = ~n721 & n6570 ;
  assign n7955 = n7953 | n7954 ;
  assign n7956 = n995 & n6567 ;
  assign n7957 = n7955 | n7956 ;
  assign n7958 = n6571 | n7957 ;
  assign n7959 = ( ~n3829 & n7957 ) | ( ~n3829 & n7958 ) | ( n7957 & n7958 ) ;
  assign n7960 = x11 & ~n7959 ;
  assign n7961 = ~x11 & n7959 ;
  assign n7962 = n7960 | n7961 ;
  assign n7963 = ( ~n7603 & n7605 ) | ( ~n7603 & n7615 ) | ( n7605 & n7615 ) ;
  assign n7964 = ( n7603 & ~n7616 ) | ( n7603 & n7963 ) | ( ~n7616 & n7963 ) ;
  assign n7965 = ( n7952 & n7962 ) | ( n7952 & n7964 ) | ( n7962 & n7964 ) ;
  assign n7966 = ~n3487 & n7341 ;
  assign n7967 = ~n3601 & n7644 ;
  assign n7968 = n3533 & n7345 ;
  assign n7969 = ( n7345 & n7967 ) | ( n7345 & ~n7968 ) | ( n7967 & ~n7968 ) ;
  assign n7970 = n7966 | n7969 ;
  assign n7971 = n7346 | n7970 ;
  assign n7972 = ( ~n4223 & n7970 ) | ( ~n4223 & n7971 ) | ( n7970 & n7971 ) ;
  assign n7973 = x8 & ~n7972 ;
  assign n7974 = ~x8 & n7972 ;
  assign n7975 = n7973 | n7974 ;
  assign n7976 = ( n7616 & n7618 ) | ( n7616 & n7628 ) | ( n7618 & n7628 ) ;
  assign n7977 = ( n7618 & n7629 ) | ( n7618 & ~n7976 ) | ( n7629 & ~n7976 ) ;
  assign n7978 = ( n7965 & n7975 ) | ( n7965 & ~n7977 ) | ( n7975 & ~n7977 ) ;
  assign n7979 = ~n3516 & n7345 ;
  assign n7980 = n7341 | n7979 ;
  assign n7981 = ( ~n3601 & n7979 ) | ( ~n3601 & n7980 ) | ( n7979 & n7980 ) ;
  assign n7982 = ~n3533 & n7644 ;
  assign n7983 = n7981 | n7982 ;
  assign n7984 = n7346 | n7983 ;
  assign n7985 = ( ~n4058 & n7983 ) | ( ~n4058 & n7984 ) | ( n7983 & n7984 ) ;
  assign n7986 = x8 & ~n7985 ;
  assign n7987 = ~x8 & n7985 ;
  assign n7988 = n7986 | n7987 ;
  assign n7989 = ( ~n7629 & n7631 ) | ( ~n7629 & n7641 ) | ( n7631 & n7641 ) ;
  assign n7990 = ( n7629 & ~n7642 ) | ( n7629 & n7989 ) | ( ~n7642 & n7989 ) ;
  assign n7991 = ( n7978 & n7988 ) | ( n7978 & n7990 ) | ( n7988 & n7990 ) ;
  assign n7992 = n5915 & n5965 ;
  assign n7993 = ~n3232 & n5909 ;
  assign n7994 = ~n3049 & n6332 ;
  assign n7995 = n7993 | n7994 ;
  assign n7996 = n3123 & n5914 ;
  assign n7997 = n7995 | n7996 ;
  assign n7998 = n7992 | n7997 ;
  assign n7999 = ~n3232 & n5911 ;
  assign n8000 = n3233 & n5911 ;
  assign n8001 = n5915 | n6332 ;
  assign n8002 = ( n3049 & n6332 ) | ( n3049 & n8001 ) | ( n6332 & n8001 ) ;
  assign n8003 = ~n3232 & n8002 ;
  assign n8004 = n3049 | n5914 ;
  assign n8005 = ( ~n3049 & n8003 ) | ( ~n3049 & n8004 ) | ( n8003 & n8004 ) ;
  assign n8006 = n8000 | n8005 ;
  assign n8007 = n7999 | n8006 ;
  assign n8008 = x14 & ~n8007 ;
  assign n8009 = ~n7998 & n8008 ;
  assign n8010 = x14 & ~n8009 ;
  assign n8011 = n5915 & n6000 ;
  assign n8012 = n3123 & n6332 ;
  assign n8013 = ~n2977 & n5914 ;
  assign n8014 = n8012 | n8013 ;
  assign n8015 = ~n3049 & n5909 ;
  assign n8016 = n8014 | n8015 ;
  assign n8017 = n8011 | n8016 ;
  assign n8018 = ( n7694 & ~n8010 ) | ( n7694 & n8017 ) | ( ~n8010 & n8017 ) ;
  assign n8019 = ( n7694 & n8010 ) | ( n7694 & ~n8017 ) | ( n8010 & ~n8017 ) ;
  assign n8020 = ( ~n7694 & n8018 ) | ( ~n7694 & n8019 ) | ( n8018 & n8019 ) ;
  assign n8021 = ( n7694 & n8009 ) | ( n7694 & ~n8020 ) | ( n8009 & ~n8020 ) ;
  assign n8022 = n3123 & n5909 ;
  assign n8023 = ~n2977 & n6332 ;
  assign n8024 = n8022 | n8023 ;
  assign n8025 = ~n2944 & n5914 ;
  assign n8026 = n8024 | n8025 ;
  assign n8027 = x14 & n8026 ;
  assign n8028 = n5915 & ~n5926 ;
  assign n8029 = x14 & ~n8028 ;
  assign n8030 = ( ~x14 & n8026 ) | ( ~x14 & n8028 ) | ( n8026 & n8028 ) ;
  assign n8031 = ( ~n8027 & n8029 ) | ( ~n8027 & n8030 ) | ( n8029 & n8030 ) ;
  assign n8032 = x17 & n7694 ;
  assign n8033 = ~n7693 & n8032 ;
  assign n8034 = n7693 & ~n8032 ;
  assign n8035 = n8033 | n8034 ;
  assign n8036 = ( n8021 & n8031 ) | ( n8021 & n8035 ) | ( n8031 & n8035 ) ;
  assign n8037 = ~n2888 & n5914 ;
  assign n8038 = ~n2977 & n5909 ;
  assign n8039 = ~n2944 & n6332 ;
  assign n8040 = n8038 | n8039 ;
  assign n8041 = n8037 | n8040 ;
  assign n8042 = x14 & n8041 ;
  assign n8043 = n5915 & ~n6055 ;
  assign n8044 = x14 & ~n8043 ;
  assign n8045 = ( ~x14 & n8041 ) | ( ~x14 & n8043 ) | ( n8041 & n8043 ) ;
  assign n8046 = ( ~n8042 & n8044 ) | ( ~n8042 & n8045 ) | ( n8044 & n8045 ) ;
  assign n8047 = x17 & ~n7696 ;
  assign n8048 = ~n7686 & n8047 ;
  assign n8049 = n7686 & ~n8047 ;
  assign n8050 = n8048 | n8049 ;
  assign n8051 = ( n8036 & n8046 ) | ( n8036 & n8050 ) | ( n8046 & n8050 ) ;
  assign n8052 = ~n2888 & n6332 ;
  assign n8053 = n2820 & n5914 ;
  assign n8054 = ~n2944 & n5909 ;
  assign n8055 = n8053 | n8054 ;
  assign n8056 = n8052 | n8055 ;
  assign n8057 = x14 & n8056 ;
  assign n8058 = n5915 & n6106 ;
  assign n8059 = ( ~x14 & n8056 ) | ( ~x14 & n8058 ) | ( n8056 & n8058 ) ;
  assign n8060 = x14 & ~n8058 ;
  assign n8061 = ( ~n8057 & n8059 ) | ( ~n8057 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8062 = ( n7701 & n8051 ) | ( n7701 & n8061 ) | ( n8051 & n8061 ) ;
  assign n8063 = n2735 & n5914 ;
  assign n8064 = n2820 & n6332 ;
  assign n8065 = n8063 | n8064 ;
  assign n8066 = ~n2888 & n5909 ;
  assign n8067 = n8065 | n8066 ;
  assign n8068 = x14 & n8067 ;
  assign n8069 = n5915 & ~n6157 ;
  assign n8070 = ( ~x14 & n8067 ) | ( ~x14 & n8069 ) | ( n8067 & n8069 ) ;
  assign n8071 = x14 & ~n8069 ;
  assign n8072 = ( ~n8068 & n8070 ) | ( ~n8068 & n8071 ) | ( n8070 & n8071 ) ;
  assign n8073 = ( ~n7665 & n7669 ) | ( ~n7665 & n7702 ) | ( n7669 & n7702 ) ;
  assign n8074 = ( n7665 & ~n7703 ) | ( n7665 & n8073 ) | ( ~n7703 & n8073 ) ;
  assign n8075 = ( n8062 & n8072 ) | ( n8062 & n8074 ) | ( n8072 & n8074 ) ;
  assign n8076 = ( ~n7703 & n7713 ) | ( ~n7703 & n7717 ) | ( n7713 & n7717 ) ;
  assign n8077 = ( n7703 & ~n7718 ) | ( n7703 & n8076 ) | ( ~n7718 & n8076 ) ;
  assign n8078 = n2735 & n6332 ;
  assign n8079 = n2642 & n5914 ;
  assign n8080 = n8078 | n8079 ;
  assign n8081 = n2820 & n5909 ;
  assign n8082 = n8080 | n8081 ;
  assign n8083 = x14 & n8082 ;
  assign n8084 = n5598 & n5915 ;
  assign n8085 = ( ~x14 & n8082 ) | ( ~x14 & n8084 ) | ( n8082 & n8084 ) ;
  assign n8086 = x14 & ~n8084 ;
  assign n8087 = ( ~n8083 & n8085 ) | ( ~n8083 & n8086 ) | ( n8085 & n8086 ) ;
  assign n8088 = ( n8075 & n8077 ) | ( n8075 & n8087 ) | ( n8077 & n8087 ) ;
  assign n8089 = n2735 & n5909 ;
  assign n8090 = n2642 & n6332 ;
  assign n8091 = ~n2608 & n5914 ;
  assign n8092 = n8090 | n8091 ;
  assign n8093 = n8089 | n8092 ;
  assign n8094 = x14 & n8093 ;
  assign n8095 = n5915 & ~n6216 ;
  assign n8096 = x14 & ~n8095 ;
  assign n8097 = ( ~x14 & n8093 ) | ( ~x14 & n8095 ) | ( n8093 & n8095 ) ;
  assign n8098 = ( ~n8094 & n8096 ) | ( ~n8094 & n8097 ) | ( n8096 & n8097 ) ;
  assign n8099 = ( ~n7718 & n7728 ) | ( ~n7718 & n7730 ) | ( n7728 & n7730 ) ;
  assign n8100 = ( n7718 & ~n7731 ) | ( n7718 & n8099 ) | ( ~n7731 & n8099 ) ;
  assign n8101 = ( n8088 & n8098 ) | ( n8088 & n8100 ) | ( n8098 & n8100 ) ;
  assign n8102 = n2642 & n5909 ;
  assign n8103 = ~n2608 & n6332 ;
  assign n8104 = n8102 | n8103 ;
  assign n8105 = ~n2521 & n5914 ;
  assign n8106 = n8104 | n8105 ;
  assign n8107 = x14 & n8106 ;
  assign n8108 = n5915 & n6221 ;
  assign n8109 = x14 & ~n8108 ;
  assign n8110 = ( ~x14 & n8106 ) | ( ~x14 & n8108 ) | ( n8106 & n8108 ) ;
  assign n8111 = ( ~n8107 & n8109 ) | ( ~n8107 & n8110 ) | ( n8109 & n8110 ) ;
  assign n8112 = ( ~n7731 & n7741 ) | ( ~n7731 & n7743 ) | ( n7741 & n7743 ) ;
  assign n8113 = ( n7731 & ~n7744 ) | ( n7731 & n8112 ) | ( ~n7744 & n8112 ) ;
  assign n8114 = ( n8101 & n8111 ) | ( n8101 & n8113 ) | ( n8111 & n8113 ) ;
  assign n8115 = ~n2467 & n5914 ;
  assign n8116 = ~n2521 & n6332 ;
  assign n8117 = ~n2608 & n5909 ;
  assign n8118 = n8116 | n8117 ;
  assign n8119 = n8115 | n8118 ;
  assign n8120 = x14 & n8119 ;
  assign n8121 = ~n5693 & n5915 ;
  assign n8122 = x14 & ~n8121 ;
  assign n8123 = ( ~x14 & n8119 ) | ( ~x14 & n8121 ) | ( n8119 & n8121 ) ;
  assign n8124 = ( ~n8120 & n8122 ) | ( ~n8120 & n8123 ) | ( n8122 & n8123 ) ;
  assign n8125 = ( ~n7744 & n7746 ) | ( ~n7744 & n7756 ) | ( n7746 & n7756 ) ;
  assign n8126 = ( n7744 & ~n7757 ) | ( n7744 & n8125 ) | ( ~n7757 & n8125 ) ;
  assign n8127 = ( n8114 & n8124 ) | ( n8114 & n8126 ) | ( n8124 & n8126 ) ;
  assign n8128 = ( ~n7757 & n7759 ) | ( ~n7757 & n7769 ) | ( n7759 & n7769 ) ;
  assign n8129 = ( n7757 & ~n7770 ) | ( n7757 & n8128 ) | ( ~n7770 & n8128 ) ;
  assign n8130 = ~n2467 & n6332 ;
  assign n8131 = ~n2521 & n5909 ;
  assign n8132 = n2398 & n5914 ;
  assign n8133 = n8131 | n8132 ;
  assign n8134 = n8130 | n8133 ;
  assign n8135 = x14 & n8134 ;
  assign n8136 = n5452 & n5915 ;
  assign n8137 = x14 & ~n8136 ;
  assign n8138 = ( ~x14 & n8134 ) | ( ~x14 & n8136 ) | ( n8134 & n8136 ) ;
  assign n8139 = ( ~n8135 & n8137 ) | ( ~n8135 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8140 = ( n8127 & n8129 ) | ( n8127 & n8139 ) | ( n8129 & n8139 ) ;
  assign n8141 = ( ~n7770 & n7772 ) | ( ~n7770 & n7782 ) | ( n7772 & n7782 ) ;
  assign n8142 = ( n7770 & ~n7783 ) | ( n7770 & n8141 ) | ( ~n7783 & n8141 ) ;
  assign n8143 = ~n2364 & n5914 ;
  assign n8144 = n2398 & n6332 ;
  assign n8145 = n8143 | n8144 ;
  assign n8146 = ~n2467 & n5909 ;
  assign n8147 = n8145 | n8146 ;
  assign n8148 = n5915 | n8147 ;
  assign n8149 = ( n5713 & n8147 ) | ( n5713 & n8148 ) | ( n8147 & n8148 ) ;
  assign n8150 = x14 & ~n8149 ;
  assign n8151 = ~x14 & n8149 ;
  assign n8152 = n8150 | n8151 ;
  assign n8153 = ( n8140 & n8142 ) | ( n8140 & n8152 ) | ( n8142 & n8152 ) ;
  assign n8154 = n2398 & n5909 ;
  assign n8155 = x14 & n8154 ;
  assign n8156 = ~n2364 & n6332 ;
  assign n8157 = ~n2282 & n5914 ;
  assign n8158 = n8156 | n8157 ;
  assign n8159 = n5915 | n8158 ;
  assign n8160 = ( ~n5494 & n8158 ) | ( ~n5494 & n8159 ) | ( n8158 & n8159 ) ;
  assign n8161 = x14 & ~n8160 ;
  assign n8162 = ( ~x14 & n8154 ) | ( ~x14 & n8160 ) | ( n8154 & n8160 ) ;
  assign n8163 = ( ~n8155 & n8161 ) | ( ~n8155 & n8162 ) | ( n8161 & n8162 ) ;
  assign n8164 = ( ~n7783 & n7793 ) | ( ~n7783 & n7795 ) | ( n7793 & n7795 ) ;
  assign n8165 = ( n7783 & ~n7796 ) | ( n7783 & n8164 ) | ( ~n7796 & n8164 ) ;
  assign n8166 = ( n8153 & n8163 ) | ( n8153 & n8165 ) | ( n8163 & n8165 ) ;
  assign n8167 = ( ~n7796 & n7798 ) | ( ~n7796 & n7808 ) | ( n7798 & n7808 ) ;
  assign n8168 = ( n7796 & ~n7809 ) | ( n7796 & n8167 ) | ( ~n7809 & n8167 ) ;
  assign n8169 = n2187 & n5914 ;
  assign n8170 = x14 & n8169 ;
  assign n8171 = ~n2364 & n5909 ;
  assign n8172 = ~n2282 & n6332 ;
  assign n8173 = n8171 | n8172 ;
  assign n8174 = n5915 | n8173 ;
  assign n8175 = ( n5137 & n8173 ) | ( n5137 & n8174 ) | ( n8173 & n8174 ) ;
  assign n8176 = x14 & ~n8175 ;
  assign n8177 = ( ~x14 & n8169 ) | ( ~x14 & n8175 ) | ( n8169 & n8175 ) ;
  assign n8178 = ( ~n8170 & n8176 ) | ( ~n8170 & n8177 ) | ( n8176 & n8177 ) ;
  assign n8179 = ( n8166 & n8168 ) | ( n8166 & n8178 ) | ( n8168 & n8178 ) ;
  assign n8180 = n2102 & n5914 ;
  assign n8181 = ~n2282 & n5909 ;
  assign n8182 = n8180 | n8181 ;
  assign n8183 = n2187 & n6332 ;
  assign n8184 = n8182 | n8183 ;
  assign n8185 = n5915 | n8184 ;
  assign n8186 = ( ~n5331 & n8184 ) | ( ~n5331 & n8185 ) | ( n8184 & n8185 ) ;
  assign n8187 = x14 & ~n8186 ;
  assign n8188 = ~x14 & n8186 ;
  assign n8189 = n8187 | n8188 ;
  assign n8190 = ( ~n7809 & n7811 ) | ( ~n7809 & n7821 ) | ( n7811 & n7821 ) ;
  assign n8191 = ( n7809 & ~n7822 ) | ( n7809 & n8190 ) | ( ~n7822 & n8190 ) ;
  assign n8192 = ( n8179 & n8189 ) | ( n8179 & n8191 ) | ( n8189 & n8191 ) ;
  assign n8193 = ( ~n7822 & n7824 ) | ( ~n7822 & n7834 ) | ( n7824 & n7834 ) ;
  assign n8194 = ( n7822 & ~n7835 ) | ( n7822 & n8193 ) | ( ~n7835 & n8193 ) ;
  assign n8195 = ~n2041 & n5914 ;
  assign n8196 = n2187 & n5909 ;
  assign n8197 = n8195 | n8196 ;
  assign n8198 = n2102 & n6332 ;
  assign n8199 = n8197 | n8198 ;
  assign n8200 = n5915 | n8199 ;
  assign n8201 = ( ~n4997 & n8199 ) | ( ~n4997 & n8200 ) | ( n8199 & n8200 ) ;
  assign n8202 = x14 & ~n8201 ;
  assign n8203 = ~x14 & n8201 ;
  assign n8204 = n8202 | n8203 ;
  assign n8205 = ( n8192 & n8194 ) | ( n8192 & n8204 ) | ( n8194 & n8204 ) ;
  assign n8206 = ( ~n7835 & n7837 ) | ( ~n7835 & n7847 ) | ( n7837 & n7847 ) ;
  assign n8207 = ( n7835 & ~n7848 ) | ( n7835 & n8206 ) | ( ~n7848 & n8206 ) ;
  assign n8208 = ~n2041 & n6332 ;
  assign n8209 = n1943 & n5914 ;
  assign n8210 = n8208 | n8209 ;
  assign n8211 = n2102 & n5909 ;
  assign n8212 = n8210 | n8211 ;
  assign n8213 = n5915 | n8212 ;
  assign n8214 = ( ~n4985 & n8212 ) | ( ~n4985 & n8213 ) | ( n8212 & n8213 ) ;
  assign n8215 = x14 & ~n8214 ;
  assign n8216 = ~x14 & n8214 ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = ( n8205 & n8207 ) | ( n8205 & n8217 ) | ( n8207 & n8217 ) ;
  assign n8219 = ~n2041 & n5909 ;
  assign n8220 = n1943 & n6332 ;
  assign n8221 = n8219 | n8220 ;
  assign n8222 = ~n1841 & n5914 ;
  assign n8223 = n8221 | n8222 ;
  assign n8224 = n5915 | n8223 ;
  assign n8225 = ( ~n4753 & n8223 ) | ( ~n4753 & n8224 ) | ( n8223 & n8224 ) ;
  assign n8226 = x14 & ~n8225 ;
  assign n8227 = ~x14 & n8225 ;
  assign n8228 = n8226 | n8227 ;
  assign n8229 = ( ~n7848 & n7850 ) | ( ~n7848 & n7860 ) | ( n7850 & n7860 ) ;
  assign n8230 = ( n7848 & ~n7861 ) | ( n7848 & n8229 ) | ( ~n7861 & n8229 ) ;
  assign n8231 = ( n8218 & n8228 ) | ( n8218 & n8230 ) | ( n8228 & n8230 ) ;
  assign n8232 = n1943 & n5909 ;
  assign n8233 = n1792 & n5914 ;
  assign n8234 = n8232 | n8233 ;
  assign n8235 = ~n1841 & n6332 ;
  assign n8236 = n8234 | n8235 ;
  assign n8237 = n5915 | n8236 ;
  assign n8238 = ( ~n4831 & n8236 ) | ( ~n4831 & n8237 ) | ( n8236 & n8237 ) ;
  assign n8239 = x14 & ~n8238 ;
  assign n8240 = ~x14 & n8238 ;
  assign n8241 = n8239 | n8240 ;
  assign n8242 = ( n7861 & ~n7871 ) | ( n7861 & n7873 ) | ( ~n7871 & n7873 ) ;
  assign n8243 = ( ~n7861 & n7874 ) | ( ~n7861 & n8242 ) | ( n7874 & n8242 ) ;
  assign n8244 = ( n8231 & n8241 ) | ( n8231 & ~n8243 ) | ( n8241 & ~n8243 ) ;
  assign n8245 = ~n1841 & n5909 ;
  assign n8246 = x14 & n8245 ;
  assign n8247 = n1687 & n5914 ;
  assign n8248 = n1792 & n6332 ;
  assign n8249 = n8247 | n8248 ;
  assign n8250 = n5915 | n8249 ;
  assign n8251 = ( n4331 & n8249 ) | ( n4331 & n8250 ) | ( n8249 & n8250 ) ;
  assign n8252 = x14 & ~n8251 ;
  assign n8253 = ( ~x14 & n8245 ) | ( ~x14 & n8251 ) | ( n8245 & n8251 ) ;
  assign n8254 = ( ~n8246 & n8252 ) | ( ~n8246 & n8253 ) | ( n8252 & n8253 ) ;
  assign n8255 = ( n7874 & ~n7884 ) | ( n7874 & n7886 ) | ( ~n7884 & n7886 ) ;
  assign n8256 = ( ~n7874 & n7887 ) | ( ~n7874 & n8255 ) | ( n7887 & n8255 ) ;
  assign n8257 = ( n8244 & n8254 ) | ( n8244 & ~n8256 ) | ( n8254 & ~n8256 ) ;
  assign n8258 = ( ~n7887 & n7897 ) | ( ~n7887 & n7899 ) | ( n7897 & n7899 ) ;
  assign n8259 = ( n7887 & ~n7900 ) | ( n7887 & n8258 ) | ( ~n7900 & n8258 ) ;
  assign n8260 = n1687 & n6332 ;
  assign n8261 = n1792 & n5909 ;
  assign n8262 = n1600 & n5914 ;
  assign n8263 = n8261 | n8262 ;
  assign n8264 = n8260 | n8263 ;
  assign n8265 = n5915 | n8264 ;
  assign n8266 = ( n4674 & n8264 ) | ( n4674 & n8265 ) | ( n8264 & n8265 ) ;
  assign n8267 = x14 & ~n8266 ;
  assign n8268 = ~x14 & n8266 ;
  assign n8269 = n8267 | n8268 ;
  assign n8270 = ( n8257 & n8259 ) | ( n8257 & n8269 ) | ( n8259 & n8269 ) ;
  assign n8271 = ~n1529 & n5914 ;
  assign n8272 = n1687 & n5909 ;
  assign n8273 = n8271 | n8272 ;
  assign n8274 = n1600 & n6332 ;
  assign n8275 = n8273 | n8274 ;
  assign n8276 = n5915 | n8275 ;
  assign n8277 = ( ~n4531 & n8275 ) | ( ~n4531 & n8276 ) | ( n8275 & n8276 ) ;
  assign n8278 = x14 & ~n8277 ;
  assign n8279 = ~x14 & n8277 ;
  assign n8280 = n8278 | n8279 ;
  assign n8281 = ( ~n7900 & n7910 ) | ( ~n7900 & n7912 ) | ( n7910 & n7912 ) ;
  assign n8282 = ( ~n7910 & n7913 ) | ( ~n7910 & n8281 ) | ( n7913 & n8281 ) ;
  assign n8283 = ( n8270 & n8280 ) | ( n8270 & ~n8282 ) | ( n8280 & ~n8282 ) ;
  assign n8284 = ( ~n7913 & n7923 ) | ( ~n7913 & n7925 ) | ( n7923 & n7925 ) ;
  assign n8285 = ( n7913 & ~n7926 ) | ( n7913 & n8284 ) | ( ~n7926 & n8284 ) ;
  assign n8286 = ~n1529 & n6332 ;
  assign n8287 = n1600 & n5909 ;
  assign n8288 = n1398 & n5914 ;
  assign n8289 = n8287 | n8288 ;
  assign n8290 = n8286 | n8289 ;
  assign n8291 = n5915 | n8290 ;
  assign n8292 = ( ~n4324 & n8290 ) | ( ~n4324 & n8291 ) | ( n8290 & n8291 ) ;
  assign n8293 = x14 & ~n8292 ;
  assign n8294 = ~x14 & n8292 ;
  assign n8295 = n8293 | n8294 ;
  assign n8296 = ( n8283 & n8285 ) | ( n8283 & n8295 ) | ( n8285 & n8295 ) ;
  assign n8297 = ( ~n7926 & n7928 ) | ( ~n7926 & n7938 ) | ( n7928 & n7938 ) ;
  assign n8298 = ( n7926 & ~n7939 ) | ( n7926 & n8297 ) | ( ~n7939 & n8297 ) ;
  assign n8299 = ~n1529 & n5909 ;
  assign n8300 = n1398 & n6332 ;
  assign n8301 = ( ~x14 & n8299 ) | ( ~x14 & n8300 ) | ( n8299 & n8300 ) ;
  assign n8302 = n1316 & n5914 ;
  assign n8303 = n5915 | n8302 ;
  assign n8304 = ( n4084 & n8302 ) | ( n4084 & n8303 ) | ( n8302 & n8303 ) ;
  assign n8305 = x14 & ~n8299 ;
  assign n8306 = n8304 | n8305 ;
  assign n8307 = ( n8300 & n8304 ) | ( n8300 & n8305 ) | ( n8304 & n8305 ) ;
  assign n8308 = ( n8301 & n8306 ) | ( n8301 & ~n8307 ) | ( n8306 & ~n8307 ) ;
  assign n8309 = ( n8296 & n8298 ) | ( n8296 & n8308 ) | ( n8298 & n8308 ) ;
  assign n8310 = ( ~n7939 & n7941 ) | ( ~n7939 & n7951 ) | ( n7941 & n7951 ) ;
  assign n8311 = ( n7939 & ~n7952 ) | ( n7939 & n8310 ) | ( ~n7952 & n8310 ) ;
  assign n8312 = n859 & n6570 ;
  assign n8313 = n995 & n6796 ;
  assign n8314 = n8312 | n8313 ;
  assign n8315 = ~n1118 & n6567 ;
  assign n8316 = n8314 | n8315 ;
  assign n8317 = n6571 | n8316 ;
  assign n8318 = ( ~n4034 & n8316 ) | ( ~n4034 & n8317 ) | ( n8316 & n8317 ) ;
  assign n8319 = x11 & ~n8318 ;
  assign n8320 = ~x11 & n8318 ;
  assign n8321 = n8319 | n8320 ;
  assign n8322 = ( n8309 & n8311 ) | ( n8309 & n8321 ) | ( n8311 & n8321 ) ;
  assign n8323 = ( ~n7952 & n7962 ) | ( ~n7952 & n7964 ) | ( n7962 & n7964 ) ;
  assign n8324 = ( n7952 & ~n7965 ) | ( n7952 & n8323 ) | ( ~n7965 & n8323 ) ;
  assign n8325 = n564 & n7341 ;
  assign n8326 = n7346 | n8325 ;
  assign n8327 = ( n3674 & n8325 ) | ( n3674 & n8326 ) | ( n8325 & n8326 ) ;
  assign n8328 = ~n3601 & n7345 ;
  assign n8329 = ( ~x8 & n8327 ) | ( ~x8 & n8328 ) | ( n8327 & n8328 ) ;
  assign n8330 = ~n3487 & n7644 ;
  assign n8331 = x8 & ~n8328 ;
  assign n8332 = n8330 | n8331 ;
  assign n8333 = ( n8327 & n8330 ) | ( n8327 & n8331 ) | ( n8330 & n8331 ) ;
  assign n8334 = ( n8329 & n8332 ) | ( n8329 & ~n8333 ) | ( n8332 & ~n8333 ) ;
  assign n8335 = ( n8322 & n8324 ) | ( n8322 & n8334 ) | ( n8324 & n8334 ) ;
  assign n8336 = x4 & n34 ;
  assign n8337 = x4 | n34 ;
  assign n8338 = n36 | n8337 ;
  assign n8339 = ~n8336 & n8338 ;
  assign n8340 = n39 & ~n8339 ;
  assign n8341 = n36 & n39 ;
  assign n8342 = ( ~n3516 & n3608 ) | ( ~n3516 & n8341 ) | ( n3608 & n8341 ) ;
  assign n8343 = ( ~n3607 & n8340 ) | ( ~n3607 & n8342 ) | ( n8340 & n8342 ) ;
  assign n8344 = x5 & ~n8343 ;
  assign n8345 = ~x5 & n8343 ;
  assign n8346 = n8344 | n8345 ;
  assign n8347 = ( ~n7965 & n7975 ) | ( ~n7965 & n7977 ) | ( n7975 & n7977 ) ;
  assign n8348 = ( ~n7975 & n7978 ) | ( ~n7975 & n8347 ) | ( n7978 & n8347 ) ;
  assign n8349 = ( n8335 & n8346 ) | ( n8335 & ~n8348 ) | ( n8346 & ~n8348 ) ;
  assign n8350 = ~n1529 & n6570 ;
  assign n8351 = n1687 & n6567 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = n1600 & n6796 ;
  assign n8354 = n8352 | n8353 ;
  assign n8355 = n6571 | n8354 ;
  assign n8356 = ( ~n4531 & n8354 ) | ( ~n4531 & n8355 ) | ( n8354 & n8355 ) ;
  assign n8357 = x11 & ~n8356 ;
  assign n8358 = ~x11 & n8356 ;
  assign n8359 = n8357 | n8358 ;
  assign n8360 = ( ~n8179 & n8189 ) | ( ~n8179 & n8191 ) | ( n8189 & n8191 ) ;
  assign n8361 = ( n8179 & ~n8192 ) | ( n8179 & n8360 ) | ( ~n8192 & n8360 ) ;
  assign n8362 = n1943 & n6796 ;
  assign n8363 = ~n2041 & n6567 ;
  assign n8364 = n8362 | n8363 ;
  assign n8365 = ~n1841 & n6570 ;
  assign n8366 = n8364 | n8365 ;
  assign n8367 = n6571 | n8366 ;
  assign n8368 = ( ~n4753 & n8366 ) | ( ~n4753 & n8367 ) | ( n8366 & n8367 ) ;
  assign n8369 = x11 & ~n8368 ;
  assign n8370 = ~x11 & n8368 ;
  assign n8371 = n8369 | n8370 ;
  assign n8372 = n3123 & n6567 ;
  assign n8373 = ~n2977 & n6796 ;
  assign n8374 = n8372 | n8373 ;
  assign n8375 = ~n2944 & n6570 ;
  assign n8376 = n8374 | n8375 ;
  assign n8377 = x11 & n8376 ;
  assign n8378 = ~n5926 & n6571 ;
  assign n8379 = x11 & ~n8378 ;
  assign n8380 = ( ~x11 & n8376 ) | ( ~x11 & n8378 ) | ( n8376 & n8378 ) ;
  assign n8381 = ( ~n8377 & n8379 ) | ( ~n8377 & n8380 ) | ( n8379 & n8380 ) ;
  assign n8382 = n3123 & n6796 ;
  assign n8383 = ~n2977 & n6570 ;
  assign n8384 = n8382 | n8383 ;
  assign n8385 = ~n3049 & n6567 ;
  assign n8386 = n8384 | n8385 ;
  assign n8387 = x11 & n8386 ;
  assign n8388 = n6000 & n6571 ;
  assign n8389 = ( ~x11 & n8386 ) | ( ~x11 & n8388 ) | ( n8386 & n8388 ) ;
  assign n8390 = x11 & ~n8388 ;
  assign n8391 = ( ~n8387 & n8389 ) | ( ~n8387 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8392 = n6571 | n6796 ;
  assign n8393 = ( n3049 & n6796 ) | ( n3049 & n8392 ) | ( n6796 & n8392 ) ;
  assign n8394 = ~n3232 & n8393 ;
  assign n8395 = ~n3232 & n6568 ;
  assign n8396 = ( n6568 & n6570 ) | ( n6568 & ~n8395 ) | ( n6570 & ~n8395 ) ;
  assign n8397 = ~n3049 & n8396 ;
  assign n8398 = n8394 | n8397 ;
  assign n8399 = x11 & ~n8395 ;
  assign n8400 = ~n8398 & n8399 ;
  assign n8401 = n5965 & n6571 ;
  assign n8402 = n3123 & n6570 ;
  assign n8403 = ~n3049 & n6796 ;
  assign n8404 = n8402 | n8403 ;
  assign n8405 = ~n3232 & n6567 ;
  assign n8406 = n8404 | n8405 ;
  assign n8407 = n8401 | n8406 ;
  assign n8408 = n8400 & ~n8407 ;
  assign n8409 = n7999 & n8391 ;
  assign n8410 = ( n8391 & n8408 ) | ( n8391 & n8409 ) | ( n8408 & n8409 ) ;
  assign n8411 = ( x14 & n8005 ) | ( x14 & n8007 ) | ( n8005 & n8007 ) ;
  assign n8412 = x14 & n5911 ;
  assign n8413 = n8005 & n8412 ;
  assign n8414 = ( n8000 & n8411 ) | ( n8000 & ~n8413 ) | ( n8411 & ~n8413 ) ;
  assign n8415 = ( n8381 & n8410 ) | ( n8381 & n8414 ) | ( n8410 & n8414 ) ;
  assign n8416 = ~n2888 & n6570 ;
  assign n8417 = ~n2977 & n6567 ;
  assign n8418 = ~n2944 & n6796 ;
  assign n8419 = n8417 | n8418 ;
  assign n8420 = n8416 | n8419 ;
  assign n8421 = x11 & n8420 ;
  assign n8422 = ~n6055 & n6571 ;
  assign n8423 = x11 & ~n8422 ;
  assign n8424 = ( ~x11 & n8420 ) | ( ~x11 & n8422 ) | ( n8420 & n8422 ) ;
  assign n8425 = ( ~n8421 & n8423 ) | ( ~n8421 & n8424 ) | ( n8423 & n8424 ) ;
  assign n8426 = x14 & n8007 ;
  assign n8427 = ~n7998 & n8426 ;
  assign n8428 = n7998 & ~n8426 ;
  assign n8429 = n8427 | n8428 ;
  assign n8430 = ( n8415 & n8425 ) | ( n8415 & n8429 ) | ( n8425 & n8429 ) ;
  assign n8431 = ~n2888 & n6796 ;
  assign n8432 = n2820 & n6570 ;
  assign n8433 = ~n2944 & n6567 ;
  assign n8434 = n8432 | n8433 ;
  assign n8435 = n8431 | n8434 ;
  assign n8436 = x11 & n8435 ;
  assign n8437 = n6106 & n6571 ;
  assign n8438 = ( ~x11 & n8435 ) | ( ~x11 & n8437 ) | ( n8435 & n8437 ) ;
  assign n8439 = x11 & ~n8437 ;
  assign n8440 = ( ~n8436 & n8438 ) | ( ~n8436 & n8439 ) | ( n8438 & n8439 ) ;
  assign n8441 = ( n8020 & n8430 ) | ( n8020 & n8440 ) | ( n8430 & n8440 ) ;
  assign n8442 = ~n2888 & n6567 ;
  assign n8443 = n2735 & n6570 ;
  assign n8444 = n2820 & n6796 ;
  assign n8445 = n8443 | n8444 ;
  assign n8446 = n8442 | n8445 ;
  assign n8447 = x11 & n8446 ;
  assign n8448 = ~n6157 & n6571 ;
  assign n8449 = x11 & ~n8448 ;
  assign n8450 = ( ~x11 & n8446 ) | ( ~x11 & n8448 ) | ( n8446 & n8448 ) ;
  assign n8451 = ( ~n8447 & n8449 ) | ( ~n8447 & n8450 ) | ( n8449 & n8450 ) ;
  assign n8452 = ( ~n8021 & n8031 ) | ( ~n8021 & n8035 ) | ( n8031 & n8035 ) ;
  assign n8453 = ( n8021 & ~n8036 ) | ( n8021 & n8452 ) | ( ~n8036 & n8452 ) ;
  assign n8454 = ( n8441 & n8451 ) | ( n8441 & n8453 ) | ( n8451 & n8453 ) ;
  assign n8455 = ( ~n8036 & n8046 ) | ( ~n8036 & n8050 ) | ( n8046 & n8050 ) ;
  assign n8456 = ( n8036 & ~n8051 ) | ( n8036 & n8455 ) | ( ~n8051 & n8455 ) ;
  assign n8457 = n2735 & n6796 ;
  assign n8458 = n2642 & n6570 ;
  assign n8459 = n8457 | n8458 ;
  assign n8460 = n2820 & n6567 ;
  assign n8461 = n8459 | n8460 ;
  assign n8462 = x11 & n8461 ;
  assign n8463 = n5598 & n6571 ;
  assign n8464 = ( ~x11 & n8461 ) | ( ~x11 & n8463 ) | ( n8461 & n8463 ) ;
  assign n8465 = x11 & ~n8463 ;
  assign n8466 = ( ~n8462 & n8464 ) | ( ~n8462 & n8465 ) | ( n8464 & n8465 ) ;
  assign n8467 = ( n8454 & n8456 ) | ( n8454 & n8466 ) | ( n8456 & n8466 ) ;
  assign n8468 = n2642 & n6796 ;
  assign n8469 = ~n2608 & n6570 ;
  assign n8470 = n8468 | n8469 ;
  assign n8471 = n2735 & n6567 ;
  assign n8472 = n8470 | n8471 ;
  assign n8473 = x11 & n8472 ;
  assign n8474 = ~n6216 & n6571 ;
  assign n8475 = ( ~x11 & n8472 ) | ( ~x11 & n8474 ) | ( n8472 & n8474 ) ;
  assign n8476 = x11 & ~n8474 ;
  assign n8477 = ( ~n8473 & n8475 ) | ( ~n8473 & n8476 ) | ( n8475 & n8476 ) ;
  assign n8478 = ( n7701 & ~n8051 ) | ( n7701 & n8061 ) | ( ~n8051 & n8061 ) ;
  assign n8479 = ( n8051 & ~n8062 ) | ( n8051 & n8478 ) | ( ~n8062 & n8478 ) ;
  assign n8480 = ( n8467 & n8477 ) | ( n8467 & n8479 ) | ( n8477 & n8479 ) ;
  assign n8481 = ( ~n8062 & n8072 ) | ( ~n8062 & n8074 ) | ( n8072 & n8074 ) ;
  assign n8482 = ( n8062 & ~n8075 ) | ( n8062 & n8481 ) | ( ~n8075 & n8481 ) ;
  assign n8483 = n2642 & n6567 ;
  assign n8484 = ~n2608 & n6796 ;
  assign n8485 = n8483 | n8484 ;
  assign n8486 = ~n2521 & n6570 ;
  assign n8487 = n8485 | n8486 ;
  assign n8488 = n6571 | n8487 ;
  assign n8489 = ( n6221 & n8487 ) | ( n6221 & n8488 ) | ( n8487 & n8488 ) ;
  assign n8490 = x11 & ~n8489 ;
  assign n8491 = ~x11 & n8489 ;
  assign n8492 = n8490 | n8491 ;
  assign n8493 = ( n8480 & n8482 ) | ( n8480 & n8492 ) | ( n8482 & n8492 ) ;
  assign n8494 = ( ~n8075 & n8077 ) | ( ~n8075 & n8087 ) | ( n8077 & n8087 ) ;
  assign n8495 = ( n8075 & ~n8088 ) | ( n8075 & n8494 ) | ( ~n8088 & n8494 ) ;
  assign n8496 = ~n2608 & n6567 ;
  assign n8497 = x11 & n8496 ;
  assign n8498 = ~n2467 & n6570 ;
  assign n8499 = ~n2521 & n6796 ;
  assign n8500 = n8498 | n8499 ;
  assign n8501 = n6571 | n8500 ;
  assign n8502 = ( ~n5693 & n8500 ) | ( ~n5693 & n8501 ) | ( n8500 & n8501 ) ;
  assign n8503 = x11 & ~n8502 ;
  assign n8504 = ( ~x11 & n8496 ) | ( ~x11 & n8502 ) | ( n8496 & n8502 ) ;
  assign n8505 = ( ~n8497 & n8503 ) | ( ~n8497 & n8504 ) | ( n8503 & n8504 ) ;
  assign n8506 = ( n8493 & n8495 ) | ( n8493 & n8505 ) | ( n8495 & n8505 ) ;
  assign n8507 = ( ~n8088 & n8098 ) | ( ~n8088 & n8100 ) | ( n8098 & n8100 ) ;
  assign n8508 = ( n8088 & ~n8101 ) | ( n8088 & n8507 ) | ( ~n8101 & n8507 ) ;
  assign n8509 = ~n2467 & n6796 ;
  assign n8510 = ~n2521 & n6567 ;
  assign n8511 = n2398 & n6570 ;
  assign n8512 = n8510 | n8511 ;
  assign n8513 = n8509 | n8512 ;
  assign n8514 = n6571 | n8513 ;
  assign n8515 = ( n5452 & n8513 ) | ( n5452 & n8514 ) | ( n8513 & n8514 ) ;
  assign n8516 = x11 & ~n8515 ;
  assign n8517 = ~x11 & n8515 ;
  assign n8518 = n8516 | n8517 ;
  assign n8519 = ( n8506 & n8508 ) | ( n8506 & n8518 ) | ( n8508 & n8518 ) ;
  assign n8520 = ( ~n8101 & n8111 ) | ( ~n8101 & n8113 ) | ( n8111 & n8113 ) ;
  assign n8521 = ( n8101 & ~n8114 ) | ( n8101 & n8520 ) | ( ~n8114 & n8520 ) ;
  assign n8522 = n2398 & n6796 ;
  assign n8523 = x11 & n8522 ;
  assign n8524 = ~n2467 & n6567 ;
  assign n8525 = ~n2364 & n6570 ;
  assign n8526 = n8524 | n8525 ;
  assign n8527 = n6571 | n8526 ;
  assign n8528 = ( n5713 & n8526 ) | ( n5713 & n8527 ) | ( n8526 & n8527 ) ;
  assign n8529 = x11 & ~n8528 ;
  assign n8530 = ( ~x11 & n8522 ) | ( ~x11 & n8528 ) | ( n8522 & n8528 ) ;
  assign n8531 = ( ~n8523 & n8529 ) | ( ~n8523 & n8530 ) | ( n8529 & n8530 ) ;
  assign n8532 = ( n8519 & n8521 ) | ( n8519 & n8531 ) | ( n8521 & n8531 ) ;
  assign n8533 = ( ~n8114 & n8124 ) | ( ~n8114 & n8126 ) | ( n8124 & n8126 ) ;
  assign n8534 = ( n8114 & ~n8127 ) | ( n8114 & n8533 ) | ( ~n8127 & n8533 ) ;
  assign n8535 = ~n2364 & n6796 ;
  assign n8536 = n2398 & n6567 ;
  assign n8537 = n8535 | n8536 ;
  assign n8538 = ~n2282 & n6570 ;
  assign n8539 = n8537 | n8538 ;
  assign n8540 = n6571 | n8539 ;
  assign n8541 = ( ~n5494 & n8539 ) | ( ~n5494 & n8540 ) | ( n8539 & n8540 ) ;
  assign n8542 = x11 & ~n8541 ;
  assign n8543 = ~x11 & n8541 ;
  assign n8544 = n8542 | n8543 ;
  assign n8545 = ( n8532 & n8534 ) | ( n8532 & n8544 ) | ( n8534 & n8544 ) ;
  assign n8546 = ~n2364 & n6567 ;
  assign n8547 = n2187 & n6570 ;
  assign n8548 = n8546 | n8547 ;
  assign n8549 = ~n2282 & n6796 ;
  assign n8550 = n8548 | n8549 ;
  assign n8551 = n6571 | n8550 ;
  assign n8552 = ( n5137 & n8550 ) | ( n5137 & n8551 ) | ( n8550 & n8551 ) ;
  assign n8553 = x11 & ~n8552 ;
  assign n8554 = ~x11 & n8552 ;
  assign n8555 = n8553 | n8554 ;
  assign n8556 = ( ~n8127 & n8129 ) | ( ~n8127 & n8139 ) | ( n8129 & n8139 ) ;
  assign n8557 = ( n8127 & ~n8140 ) | ( n8127 & n8556 ) | ( ~n8140 & n8556 ) ;
  assign n8558 = ( n8545 & n8555 ) | ( n8545 & n8557 ) | ( n8555 & n8557 ) ;
  assign n8559 = ( ~n8140 & n8142 ) | ( ~n8140 & n8152 ) | ( n8142 & n8152 ) ;
  assign n8560 = ( n8140 & ~n8153 ) | ( n8140 & n8559 ) | ( ~n8153 & n8559 ) ;
  assign n8561 = n2102 & n6570 ;
  assign n8562 = ~n2282 & n6567 ;
  assign n8563 = n8561 | n8562 ;
  assign n8564 = n2187 & n6796 ;
  assign n8565 = n8563 | n8564 ;
  assign n8566 = n6571 | n8565 ;
  assign n8567 = ( ~n5331 & n8565 ) | ( ~n5331 & n8566 ) | ( n8565 & n8566 ) ;
  assign n8568 = x11 & ~n8567 ;
  assign n8569 = ~x11 & n8567 ;
  assign n8570 = n8568 | n8569 ;
  assign n8571 = ( n8558 & n8560 ) | ( n8558 & n8570 ) | ( n8560 & n8570 ) ;
  assign n8572 = ( ~n8153 & n8163 ) | ( ~n8153 & n8165 ) | ( n8163 & n8165 ) ;
  assign n8573 = ( n8153 & ~n8166 ) | ( n8153 & n8572 ) | ( ~n8166 & n8572 ) ;
  assign n8574 = ~n2041 & n6570 ;
  assign n8575 = n2187 & n6567 ;
  assign n8576 = n8574 | n8575 ;
  assign n8577 = n2102 & n6796 ;
  assign n8578 = n8576 | n8577 ;
  assign n8579 = n6571 | n8578 ;
  assign n8580 = ( ~n4997 & n8578 ) | ( ~n4997 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = x11 & ~n8580 ;
  assign n8582 = ~x11 & n8580 ;
  assign n8583 = n8581 | n8582 ;
  assign n8584 = ( n8571 & n8573 ) | ( n8571 & n8583 ) | ( n8573 & n8583 ) ;
  assign n8585 = ( ~n8166 & n8168 ) | ( ~n8166 & n8178 ) | ( n8168 & n8178 ) ;
  assign n8586 = ( n8166 & ~n8179 ) | ( n8166 & n8585 ) | ( ~n8179 & n8585 ) ;
  assign n8587 = n1943 & n6570 ;
  assign n8588 = x11 & n8587 ;
  assign n8589 = n2102 & n6567 ;
  assign n8590 = ~n2041 & n6796 ;
  assign n8591 = n8589 | n8590 ;
  assign n8592 = n6571 | n8591 ;
  assign n8593 = ( ~n4985 & n8591 ) | ( ~n4985 & n8592 ) | ( n8591 & n8592 ) ;
  assign n8594 = x11 & ~n8593 ;
  assign n8595 = ( ~x11 & n8587 ) | ( ~x11 & n8593 ) | ( n8587 & n8593 ) ;
  assign n8596 = ( ~n8588 & n8594 ) | ( ~n8588 & n8595 ) | ( n8594 & n8595 ) ;
  assign n8597 = ( n8584 & n8586 ) | ( n8584 & n8596 ) | ( n8586 & n8596 ) ;
  assign n8598 = ( n8361 & n8371 ) | ( n8361 & n8597 ) | ( n8371 & n8597 ) ;
  assign n8599 = n1943 & n6567 ;
  assign n8600 = n1792 & n6570 ;
  assign n8601 = n8599 | n8600 ;
  assign n8602 = ~n1841 & n6796 ;
  assign n8603 = n8601 | n8602 ;
  assign n8604 = n6571 | n8603 ;
  assign n8605 = ( ~n4831 & n8603 ) | ( ~n4831 & n8604 ) | ( n8603 & n8604 ) ;
  assign n8606 = x11 & ~n8605 ;
  assign n8607 = ~x11 & n8605 ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = ( ~n8192 & n8194 ) | ( ~n8192 & n8204 ) | ( n8194 & n8204 ) ;
  assign n8610 = ( n8192 & ~n8205 ) | ( n8192 & n8609 ) | ( ~n8205 & n8609 ) ;
  assign n8611 = ( n8598 & n8608 ) | ( n8598 & n8610 ) | ( n8608 & n8610 ) ;
  assign n8612 = ( ~n8205 & n8207 ) | ( ~n8205 & n8217 ) | ( n8207 & n8217 ) ;
  assign n8613 = ( n8205 & ~n8218 ) | ( n8205 & n8612 ) | ( ~n8218 & n8612 ) ;
  assign n8614 = ~n1841 & n6567 ;
  assign n8615 = x11 & n8614 ;
  assign n8616 = n1687 & n6570 ;
  assign n8617 = n1792 & n6796 ;
  assign n8618 = n8616 | n8617 ;
  assign n8619 = n6571 | n8618 ;
  assign n8620 = ( n4331 & n8618 ) | ( n4331 & n8619 ) | ( n8618 & n8619 ) ;
  assign n8621 = x11 & ~n8620 ;
  assign n8622 = ( ~x11 & n8614 ) | ( ~x11 & n8620 ) | ( n8614 & n8620 ) ;
  assign n8623 = ( ~n8615 & n8621 ) | ( ~n8615 & n8622 ) | ( n8621 & n8622 ) ;
  assign n8624 = ( n8611 & n8613 ) | ( n8611 & n8623 ) | ( n8613 & n8623 ) ;
  assign n8625 = ( ~n8218 & n8228 ) | ( ~n8218 & n8230 ) | ( n8228 & n8230 ) ;
  assign n8626 = ( n8218 & ~n8231 ) | ( n8218 & n8625 ) | ( ~n8231 & n8625 ) ;
  assign n8627 = n1687 & n6796 ;
  assign n8628 = n1792 & n6567 ;
  assign n8629 = n1600 & n6570 ;
  assign n8630 = n8628 | n8629 ;
  assign n8631 = n8627 | n8630 ;
  assign n8632 = n6571 | n8631 ;
  assign n8633 = ( n4674 & n8631 ) | ( n4674 & n8632 ) | ( n8631 & n8632 ) ;
  assign n8634 = x11 & ~n8633 ;
  assign n8635 = ~x11 & n8633 ;
  assign n8636 = n8634 | n8635 ;
  assign n8637 = ( n8624 & n8626 ) | ( n8624 & n8636 ) | ( n8626 & n8636 ) ;
  assign n8638 = ( n8231 & n8241 ) | ( n8231 & n8243 ) | ( n8241 & n8243 ) ;
  assign n8639 = ( n8243 & n8244 ) | ( n8243 & ~n8638 ) | ( n8244 & ~n8638 ) ;
  assign n8640 = ( n8359 & n8637 ) | ( n8359 & ~n8639 ) | ( n8637 & ~n8639 ) ;
  assign n8641 = ~n1529 & n6796 ;
  assign n8642 = n1600 & n6567 ;
  assign n8643 = n1398 & n6570 ;
  assign n8644 = n8642 | n8643 ;
  assign n8645 = n8641 | n8644 ;
  assign n8646 = n6571 | n8645 ;
  assign n8647 = ( ~n4324 & n8645 ) | ( ~n4324 & n8646 ) | ( n8645 & n8646 ) ;
  assign n8648 = x11 & ~n8647 ;
  assign n8649 = ~x11 & n8647 ;
  assign n8650 = n8648 | n8649 ;
  assign n8651 = ( n8244 & ~n8254 ) | ( n8244 & n8256 ) | ( ~n8254 & n8256 ) ;
  assign n8652 = ( ~n8244 & n8257 ) | ( ~n8244 & n8651 ) | ( n8257 & n8651 ) ;
  assign n8653 = ( n8640 & n8650 ) | ( n8640 & ~n8652 ) | ( n8650 & ~n8652 ) ;
  assign n8654 = ( ~n8257 & n8259 ) | ( ~n8257 & n8269 ) | ( n8259 & n8269 ) ;
  assign n8655 = ( n8257 & ~n8270 ) | ( n8257 & n8654 ) | ( ~n8270 & n8654 ) ;
  assign n8656 = n1398 & n6796 ;
  assign n8657 = x11 & n8656 ;
  assign n8658 = ~n1529 & n6567 ;
  assign n8659 = n1316 & n6570 ;
  assign n8660 = n8658 | n8659 ;
  assign n8661 = n6571 | n8660 ;
  assign n8662 = ( n4084 & n8660 ) | ( n4084 & n8661 ) | ( n8660 & n8661 ) ;
  assign n8663 = x11 & ~n8662 ;
  assign n8664 = ( ~x11 & n8656 ) | ( ~x11 & n8662 ) | ( n8656 & n8662 ) ;
  assign n8665 = ( ~n8657 & n8663 ) | ( ~n8657 & n8664 ) | ( n8663 & n8664 ) ;
  assign n8666 = ( n8653 & n8655 ) | ( n8653 & n8665 ) | ( n8655 & n8665 ) ;
  assign n8667 = n1316 & n6796 ;
  assign n8668 = ~n1207 & n6570 ;
  assign n8669 = n1398 & n6567 ;
  assign n8670 = n8668 | n8669 ;
  assign n8671 = n8667 | n8670 ;
  assign n8672 = n6571 | n8671 ;
  assign n8673 = ( ~n4157 & n8671 ) | ( ~n4157 & n8672 ) | ( n8671 & n8672 ) ;
  assign n8674 = x11 & ~n8673 ;
  assign n8675 = ~x11 & n8673 ;
  assign n8676 = n8674 | n8675 ;
  assign n8677 = ( n8270 & n8280 ) | ( n8270 & n8282 ) | ( n8280 & n8282 ) ;
  assign n8678 = ( n8282 & n8283 ) | ( n8282 & ~n8677 ) | ( n8283 & ~n8677 ) ;
  assign n8679 = ( n8666 & n8676 ) | ( n8666 & ~n8678 ) | ( n8676 & ~n8678 ) ;
  assign n8680 = ( ~n8283 & n8285 ) | ( ~n8283 & n8295 ) | ( n8285 & n8295 ) ;
  assign n8681 = ( n8283 & ~n8296 ) | ( n8283 & n8680 ) | ( ~n8296 & n8680 ) ;
  assign n8682 = n1316 & n6567 ;
  assign n8683 = ~n1207 & n6796 ;
  assign n8684 = n8682 | n8683 ;
  assign n8685 = ~n1118 & n6570 ;
  assign n8686 = n8684 | n8685 ;
  assign n8687 = n6571 | n8686 ;
  assign n8688 = ( n3841 & n8686 ) | ( n3841 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8689 = x11 & ~n8688 ;
  assign n8690 = ~x11 & n8688 ;
  assign n8691 = n8689 | n8690 ;
  assign n8692 = ( n8679 & n8681 ) | ( n8679 & n8691 ) | ( n8681 & n8691 ) ;
  assign n8693 = n995 & n6570 ;
  assign n8694 = ~n1207 & n6567 ;
  assign n8695 = n8693 | n8694 ;
  assign n8696 = ~n1118 & n6796 ;
  assign n8697 = n8695 | n8696 ;
  assign n8698 = n6571 | n8697 ;
  assign n8699 = ( n4173 & n8697 ) | ( n4173 & n8698 ) | ( n8697 & n8698 ) ;
  assign n8700 = x11 & ~n8699 ;
  assign n8701 = ~x11 & n8699 ;
  assign n8702 = n8700 | n8701 ;
  assign n8703 = ( ~n8296 & n8298 ) | ( ~n8296 & n8308 ) | ( n8298 & n8308 ) ;
  assign n8704 = ( n8296 & ~n8309 ) | ( n8296 & n8703 ) | ( ~n8309 & n8703 ) ;
  assign n8705 = ( n8692 & n8702 ) | ( n8692 & n8704 ) | ( n8702 & n8704 ) ;
  assign n8706 = ~n3487 & n7345 ;
  assign n8707 = ~n721 & n7341 ;
  assign n8708 = n564 & n7644 ;
  assign n8709 = n8707 | n8708 ;
  assign n8710 = n8706 | n8709 ;
  assign n8711 = n7346 | n8710 ;
  assign n8712 = ( ~n3492 & n8710 ) | ( ~n3492 & n8711 ) | ( n8710 & n8711 ) ;
  assign n8713 = x8 & ~n8712 ;
  assign n8714 = ~x8 & n8712 ;
  assign n8715 = n8713 | n8714 ;
  assign n8716 = ( ~n8309 & n8311 ) | ( ~n8309 & n8321 ) | ( n8311 & n8321 ) ;
  assign n8717 = ( n8309 & ~n8322 ) | ( n8309 & n8716 ) | ( ~n8322 & n8716 ) ;
  assign n8718 = ( n8705 & n8715 ) | ( n8705 & n8717 ) | ( n8715 & n8717 ) ;
  assign n8719 = ~n3533 & n8340 ;
  assign n8720 = x5 & n8719 ;
  assign n8721 = ~n36 & n8339 ;
  assign n8722 = ~n3516 & n8721 ;
  assign n8723 = n8341 | n8722 ;
  assign n8724 = ( n3609 & n8722 ) | ( n3609 & n8723 ) | ( n8722 & n8723 ) ;
  assign n8725 = x5 & ~n8724 ;
  assign n8726 = ( ~x5 & n8719 ) | ( ~x5 & n8724 ) | ( n8719 & n8724 ) ;
  assign n8727 = ( ~n8720 & n8725 ) | ( ~n8720 & n8726 ) | ( n8725 & n8726 ) ;
  assign n8728 = ( ~n8322 & n8324 ) | ( ~n8322 & n8334 ) | ( n8324 & n8334 ) ;
  assign n8729 = ( n8322 & ~n8335 ) | ( n8322 & n8728 ) | ( ~n8335 & n8728 ) ;
  assign n8730 = ( n8718 & n8727 ) | ( n8718 & n8729 ) | ( n8727 & n8729 ) ;
  assign n8731 = ( ~n8705 & n8715 ) | ( ~n8705 & n8717 ) | ( n8715 & n8717 ) ;
  assign n8732 = ( n8705 & ~n8718 ) | ( n8705 & n8731 ) | ( ~n8718 & n8731 ) ;
  assign n8733 = n40 & ~n3516 ;
  assign n8734 = n8340 | n8733 ;
  assign n8735 = ( ~n3601 & n8733 ) | ( ~n3601 & n8734 ) | ( n8733 & n8734 ) ;
  assign n8736 = ~n3533 & n8721 ;
  assign n8737 = n8735 | n8736 ;
  assign n8738 = n8341 | n8737 ;
  assign n8739 = ( ~n4058 & n8737 ) | ( ~n4058 & n8738 ) | ( n8737 & n8738 ) ;
  assign n8740 = x5 & ~n8739 ;
  assign n8741 = ~x5 & n8739 ;
  assign n8742 = n8740 | n8741 ;
  assign n8743 = n3123 & n7341 ;
  assign n8744 = ~n2977 & n7644 ;
  assign n8745 = n8743 | n8744 ;
  assign n8746 = ~n2944 & n7345 ;
  assign n8747 = n8745 | n8746 ;
  assign n8748 = x8 & n8747 ;
  assign n8749 = ~n5926 & n7346 ;
  assign n8750 = x8 & ~n8749 ;
  assign n8751 = ( ~x8 & n8747 ) | ( ~x8 & n8749 ) | ( n8747 & n8749 ) ;
  assign n8752 = ( ~n8748 & n8750 ) | ( ~n8748 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8753 = x11 & n8395 ;
  assign n8754 = ~n8398 & n8753 ;
  assign n8755 = n8398 & ~n8753 ;
  assign n8756 = n8754 | n8755 ;
  assign n8757 = n3123 & n7644 ;
  assign n8758 = ~n2977 & n7345 ;
  assign n8759 = n8757 | n8758 ;
  assign n8760 = ~n3049 & n7341 ;
  assign n8761 = n8759 | n8760 ;
  assign n8762 = x8 & n8761 ;
  assign n8763 = n6000 & n7346 ;
  assign n8764 = ( ~x8 & n8761 ) | ( ~x8 & n8763 ) | ( n8761 & n8763 ) ;
  assign n8765 = x8 & ~n8763 ;
  assign n8766 = ( ~n8762 & n8764 ) | ( ~n8762 & n8765 ) | ( n8764 & n8765 ) ;
  assign n8767 = n3233 & n7342 ;
  assign n8768 = n7346 | n7644 ;
  assign n8769 = ( n3049 & n7644 ) | ( n3049 & n8768 ) | ( n7644 & n8768 ) ;
  assign n8770 = ~n3232 & n8769 ;
  assign n8771 = n3049 | n7345 ;
  assign n8772 = ( ~n3049 & n8770 ) | ( ~n3049 & n8771 ) | ( n8770 & n8771 ) ;
  assign n8773 = n8767 | n8772 ;
  assign n8774 = ~n3232 & n7342 ;
  assign n8775 = x8 & ~n8774 ;
  assign n8776 = ~n8773 & n8775 ;
  assign n8777 = n5965 & n7346 ;
  assign n8778 = n3123 & n7345 ;
  assign n8779 = ~n3049 & n7644 ;
  assign n8780 = n8778 | n8779 ;
  assign n8781 = ~n3232 & n7341 ;
  assign n8782 = n8780 | n8781 ;
  assign n8783 = n8777 | n8782 ;
  assign n8784 = n8776 & ~n8783 ;
  assign n8785 = n8395 & n8766 ;
  assign n8786 = ( n8766 & n8784 ) | ( n8766 & n8785 ) | ( n8784 & n8785 ) ;
  assign n8787 = ( n8752 & n8756 ) | ( n8752 & n8786 ) | ( n8756 & n8786 ) ;
  assign n8788 = ~n2888 & n7345 ;
  assign n8789 = ~n2977 & n7341 ;
  assign n8790 = ~n2944 & n7644 ;
  assign n8791 = n8789 | n8790 ;
  assign n8792 = n8788 | n8791 ;
  assign n8793 = x8 & n8792 ;
  assign n8794 = ~n6055 & n7346 ;
  assign n8795 = x8 & ~n8794 ;
  assign n8796 = ( ~x8 & n8792 ) | ( ~x8 & n8794 ) | ( n8792 & n8794 ) ;
  assign n8797 = ( ~n8793 & n8795 ) | ( ~n8793 & n8796 ) | ( n8795 & n8796 ) ;
  assign n8798 = x11 & ~n8400 ;
  assign n8799 = ~n8407 & n8798 ;
  assign n8800 = n8407 & ~n8798 ;
  assign n8801 = n8799 | n8800 ;
  assign n8802 = ( n8787 & n8797 ) | ( n8787 & n8801 ) | ( n8797 & n8801 ) ;
  assign n8803 = ~n2888 & n7644 ;
  assign n8804 = ~n2944 & n7341 ;
  assign n8805 = n2820 & n7345 ;
  assign n8806 = n8804 | n8805 ;
  assign n8807 = n8803 | n8806 ;
  assign n8808 = x8 & n8807 ;
  assign n8809 = n6106 & n7346 ;
  assign n8810 = x8 & ~n8809 ;
  assign n8811 = ( ~x8 & n8807 ) | ( ~x8 & n8809 ) | ( n8807 & n8809 ) ;
  assign n8812 = ( ~n8808 & n8810 ) | ( ~n8808 & n8811 ) | ( n8810 & n8811 ) ;
  assign n8813 = ( n7999 & ~n8391 ) | ( n7999 & n8408 ) | ( ~n8391 & n8408 ) ;
  assign n8814 = ( n8391 & ~n8410 ) | ( n8391 & n8813 ) | ( ~n8410 & n8813 ) ;
  assign n8815 = ( n8802 & n8812 ) | ( n8802 & n8814 ) | ( n8812 & n8814 ) ;
  assign n8816 = ~n2888 & n7341 ;
  assign n8817 = x8 & n8816 ;
  assign n8818 = n2735 & n7345 ;
  assign n8819 = n2820 & n7644 ;
  assign n8820 = n8818 | n8819 ;
  assign n8821 = n7346 | n8820 ;
  assign n8822 = ( ~n6157 & n8820 ) | ( ~n6157 & n8821 ) | ( n8820 & n8821 ) ;
  assign n8823 = x8 & ~n8822 ;
  assign n8824 = ( ~x8 & n8816 ) | ( ~x8 & n8822 ) | ( n8816 & n8822 ) ;
  assign n8825 = ( ~n8817 & n8823 ) | ( ~n8817 & n8824 ) | ( n8823 & n8824 ) ;
  assign n8826 = ( ~n8381 & n8410 ) | ( ~n8381 & n8414 ) | ( n8410 & n8414 ) ;
  assign n8827 = ( n8381 & ~n8415 ) | ( n8381 & n8826 ) | ( ~n8415 & n8826 ) ;
  assign n8828 = ( n8815 & n8825 ) | ( n8815 & n8827 ) | ( n8825 & n8827 ) ;
  assign n8829 = ( ~n8415 & n8425 ) | ( ~n8415 & n8429 ) | ( n8425 & n8429 ) ;
  assign n8830 = ( n8415 & ~n8430 ) | ( n8415 & n8829 ) | ( ~n8430 & n8829 ) ;
  assign n8831 = n2820 & n7341 ;
  assign n8832 = x8 & n8831 ;
  assign n8833 = n2735 & n7644 ;
  assign n8834 = n2642 & n7345 ;
  assign n8835 = n8833 | n8834 ;
  assign n8836 = n7346 | n8835 ;
  assign n8837 = ( n5598 & n8835 ) | ( n5598 & n8836 ) | ( n8835 & n8836 ) ;
  assign n8838 = x8 & ~n8837 ;
  assign n8839 = ( ~x8 & n8831 ) | ( ~x8 & n8837 ) | ( n8831 & n8837 ) ;
  assign n8840 = ( ~n8832 & n8838 ) | ( ~n8832 & n8839 ) | ( n8838 & n8839 ) ;
  assign n8841 = ( n8828 & n8830 ) | ( n8828 & n8840 ) | ( n8830 & n8840 ) ;
  assign n8842 = n2735 & n7341 ;
  assign n8843 = n2642 & n7644 ;
  assign n8844 = ~n2608 & n7345 ;
  assign n8845 = n8843 | n8844 ;
  assign n8846 = n8842 | n8845 ;
  assign n8847 = n7346 | n8846 ;
  assign n8848 = ( ~n6216 & n8846 ) | ( ~n6216 & n8847 ) | ( n8846 & n8847 ) ;
  assign n8849 = x8 & ~n8848 ;
  assign n8850 = ~x8 & n8848 ;
  assign n8851 = n8849 | n8850 ;
  assign n8852 = ( n8020 & ~n8430 ) | ( n8020 & n8440 ) | ( ~n8430 & n8440 ) ;
  assign n8853 = ( n8430 & ~n8441 ) | ( n8430 & n8852 ) | ( ~n8441 & n8852 ) ;
  assign n8854 = ( n8841 & n8851 ) | ( n8841 & n8853 ) | ( n8851 & n8853 ) ;
  assign n8855 = n2642 & n7341 ;
  assign n8856 = ~n2608 & n7644 ;
  assign n8857 = n8855 | n8856 ;
  assign n8858 = ~n2521 & n7345 ;
  assign n8859 = n8857 | n8858 ;
  assign n8860 = n7346 | n8859 ;
  assign n8861 = ( n6221 & n8859 ) | ( n6221 & n8860 ) | ( n8859 & n8860 ) ;
  assign n8862 = x8 & ~n8861 ;
  assign n8863 = ~x8 & n8861 ;
  assign n8864 = n8862 | n8863 ;
  assign n8865 = ( ~n8441 & n8451 ) | ( ~n8441 & n8453 ) | ( n8451 & n8453 ) ;
  assign n8866 = ( n8441 & ~n8454 ) | ( n8441 & n8865 ) | ( ~n8454 & n8865 ) ;
  assign n8867 = ( n8854 & n8864 ) | ( n8854 & n8866 ) | ( n8864 & n8866 ) ;
  assign n8868 = ( ~n8454 & n8456 ) | ( ~n8454 & n8466 ) | ( n8456 & n8466 ) ;
  assign n8869 = ( n8454 & ~n8467 ) | ( n8454 & n8868 ) | ( ~n8467 & n8868 ) ;
  assign n8870 = ~n2467 & n7345 ;
  assign n8871 = ~n2521 & n7644 ;
  assign n8872 = ~n2608 & n7341 ;
  assign n8873 = n8871 | n8872 ;
  assign n8874 = n8870 | n8873 ;
  assign n8875 = n7346 | n8874 ;
  assign n8876 = ( ~n5693 & n8874 ) | ( ~n5693 & n8875 ) | ( n8874 & n8875 ) ;
  assign n8877 = x8 & ~n8876 ;
  assign n8878 = ~x8 & n8876 ;
  assign n8879 = n8877 | n8878 ;
  assign n8880 = ( n8867 & n8869 ) | ( n8867 & n8879 ) | ( n8869 & n8879 ) ;
  assign n8881 = ( ~n8467 & n8477 ) | ( ~n8467 & n8479 ) | ( n8477 & n8479 ) ;
  assign n8882 = ( n8467 & ~n8480 ) | ( n8467 & n8881 ) | ( ~n8480 & n8881 ) ;
  assign n8883 = ~n2467 & n7644 ;
  assign n8884 = ~n2521 & n7341 ;
  assign n8885 = n2398 & n7345 ;
  assign n8886 = n8884 | n8885 ;
  assign n8887 = n8883 | n8886 ;
  assign n8888 = n7346 | n8887 ;
  assign n8889 = ( n5452 & n8887 ) | ( n5452 & n8888 ) | ( n8887 & n8888 ) ;
  assign n8890 = x8 & ~n8889 ;
  assign n8891 = ~x8 & n8889 ;
  assign n8892 = n8890 | n8891 ;
  assign n8893 = ( n8880 & n8882 ) | ( n8880 & n8892 ) | ( n8882 & n8892 ) ;
  assign n8894 = ( ~n8480 & n8482 ) | ( ~n8480 & n8492 ) | ( n8482 & n8492 ) ;
  assign n8895 = ( n8480 & ~n8493 ) | ( n8480 & n8894 ) | ( ~n8493 & n8894 ) ;
  assign n8896 = ~n2364 & n7345 ;
  assign n8897 = n2398 & n7644 ;
  assign n8898 = n8896 | n8897 ;
  assign n8899 = ~n2467 & n7341 ;
  assign n8900 = n8898 | n8899 ;
  assign n8901 = n7346 | n8900 ;
  assign n8902 = ( n5713 & n8900 ) | ( n5713 & n8901 ) | ( n8900 & n8901 ) ;
  assign n8903 = x8 & ~n8902 ;
  assign n8904 = ~x8 & n8902 ;
  assign n8905 = n8903 | n8904 ;
  assign n8906 = ( n8893 & n8895 ) | ( n8893 & n8905 ) | ( n8895 & n8905 ) ;
  assign n8907 = ( ~n8493 & n8495 ) | ( ~n8493 & n8505 ) | ( n8495 & n8505 ) ;
  assign n8908 = ( n8493 & ~n8506 ) | ( n8493 & n8907 ) | ( ~n8506 & n8907 ) ;
  assign n8909 = ~n2364 & n7644 ;
  assign n8910 = n2398 & n7341 ;
  assign n8911 = n8909 | n8910 ;
  assign n8912 = ~n2282 & n7345 ;
  assign n8913 = n8911 | n8912 ;
  assign n8914 = n7346 | n8913 ;
  assign n8915 = ( ~n5494 & n8913 ) | ( ~n5494 & n8914 ) | ( n8913 & n8914 ) ;
  assign n8916 = x8 & ~n8915 ;
  assign n8917 = ~x8 & n8915 ;
  assign n8918 = n8916 | n8917 ;
  assign n8919 = ( n8906 & n8908 ) | ( n8906 & n8918 ) | ( n8908 & n8918 ) ;
  assign n8920 = ( n8506 & ~n8508 ) | ( n8506 & n8518 ) | ( ~n8508 & n8518 ) ;
  assign n8921 = ( n8508 & ~n8519 ) | ( n8508 & n8920 ) | ( ~n8519 & n8920 ) ;
  assign n8922 = ~n2364 & n7341 ;
  assign n8923 = n2187 & n7345 ;
  assign n8924 = n8922 | n8923 ;
  assign n8925 = ~n2282 & n7644 ;
  assign n8926 = n8924 | n8925 ;
  assign n8927 = n7346 | n8926 ;
  assign n8928 = ( n5137 & n8926 ) | ( n5137 & n8927 ) | ( n8926 & n8927 ) ;
  assign n8929 = x8 & ~n8928 ;
  assign n8930 = ~x8 & n8928 ;
  assign n8931 = n8929 | n8930 ;
  assign n8932 = ( n8919 & n8921 ) | ( n8919 & n8931 ) | ( n8921 & n8931 ) ;
  assign n8933 = ( n8519 & ~n8521 ) | ( n8519 & n8531 ) | ( ~n8521 & n8531 ) ;
  assign n8934 = ( n8521 & ~n8532 ) | ( n8521 & n8933 ) | ( ~n8532 & n8933 ) ;
  assign n8935 = n2102 & n7345 ;
  assign n8936 = ~n2282 & n7341 ;
  assign n8937 = n8935 | n8936 ;
  assign n8938 = n2187 & n7644 ;
  assign n8939 = n8937 | n8938 ;
  assign n8940 = n7346 | n8939 ;
  assign n8941 = ( ~n5331 & n8939 ) | ( ~n5331 & n8940 ) | ( n8939 & n8940 ) ;
  assign n8942 = x8 & ~n8941 ;
  assign n8943 = ~x8 & n8941 ;
  assign n8944 = n8942 | n8943 ;
  assign n8945 = ( n8932 & n8934 ) | ( n8932 & n8944 ) | ( n8934 & n8944 ) ;
  assign n8946 = ( ~n8532 & n8534 ) | ( ~n8532 & n8544 ) | ( n8534 & n8544 ) ;
  assign n8947 = ( n8532 & ~n8545 ) | ( n8532 & n8946 ) | ( ~n8545 & n8946 ) ;
  assign n8948 = ~n2041 & n7345 ;
  assign n8949 = n2187 & n7341 ;
  assign n8950 = n8948 | n8949 ;
  assign n8951 = n2102 & n7644 ;
  assign n8952 = n8950 | n8951 ;
  assign n8953 = n7346 | n8952 ;
  assign n8954 = ( ~n4997 & n8952 ) | ( ~n4997 & n8953 ) | ( n8952 & n8953 ) ;
  assign n8955 = x8 & ~n8954 ;
  assign n8956 = ~x8 & n8954 ;
  assign n8957 = n8955 | n8956 ;
  assign n8958 = ( n8945 & n8947 ) | ( n8945 & n8957 ) | ( n8947 & n8957 ) ;
  assign n8959 = ( ~n8545 & n8555 ) | ( ~n8545 & n8557 ) | ( n8555 & n8557 ) ;
  assign n8960 = ( n8545 & ~n8558 ) | ( n8545 & n8959 ) | ( ~n8558 & n8959 ) ;
  assign n8961 = ~n2041 & n7644 ;
  assign n8962 = n1943 & n7345 ;
  assign n8963 = n8961 | n8962 ;
  assign n8964 = n2102 & n7341 ;
  assign n8965 = n8963 | n8964 ;
  assign n8966 = n7346 | n8965 ;
  assign n8967 = ( ~n4985 & n8965 ) | ( ~n4985 & n8966 ) | ( n8965 & n8966 ) ;
  assign n8968 = x8 & ~n8967 ;
  assign n8969 = ~x8 & n8967 ;
  assign n8970 = n8968 | n8969 ;
  assign n8971 = ( n8958 & n8960 ) | ( n8958 & n8970 ) | ( n8960 & n8970 ) ;
  assign n8972 = ( ~n8558 & n8560 ) | ( ~n8558 & n8570 ) | ( n8560 & n8570 ) ;
  assign n8973 = ( n8558 & ~n8571 ) | ( n8558 & n8972 ) | ( ~n8571 & n8972 ) ;
  assign n8974 = ~n2041 & n7341 ;
  assign n8975 = n1943 & n7644 ;
  assign n8976 = n8974 | n8975 ;
  assign n8977 = ~n1841 & n7345 ;
  assign n8978 = n8976 | n8977 ;
  assign n8979 = n7346 | n8978 ;
  assign n8980 = ( ~n4753 & n8978 ) | ( ~n4753 & n8979 ) | ( n8978 & n8979 ) ;
  assign n8981 = x8 & ~n8980 ;
  assign n8982 = ~x8 & n8980 ;
  assign n8983 = n8981 | n8982 ;
  assign n8984 = ( n8971 & n8973 ) | ( n8971 & n8983 ) | ( n8973 & n8983 ) ;
  assign n8985 = n1943 & n7341 ;
  assign n8986 = ~n1841 & n7644 ;
  assign n8987 = n8985 | n8986 ;
  assign n8988 = n1792 & n7345 ;
  assign n8989 = n8987 | n8988 ;
  assign n8990 = n7346 | n8989 ;
  assign n8991 = ( ~n4831 & n8989 ) | ( ~n4831 & n8990 ) | ( n8989 & n8990 ) ;
  assign n8992 = x8 & ~n8991 ;
  assign n8993 = ~x8 & n8991 ;
  assign n8994 = n8992 | n8993 ;
  assign n8995 = ( n8571 & ~n8573 ) | ( n8571 & n8583 ) | ( ~n8573 & n8583 ) ;
  assign n8996 = ( n8573 & ~n8584 ) | ( n8573 & n8995 ) | ( ~n8584 & n8995 ) ;
  assign n8997 = ( n8984 & n8994 ) | ( n8984 & n8996 ) | ( n8994 & n8996 ) ;
  assign n8998 = ( ~n8584 & n8586 ) | ( ~n8584 & n8596 ) | ( n8586 & n8596 ) ;
  assign n8999 = ( n8584 & ~n8597 ) | ( n8584 & n8998 ) | ( ~n8597 & n8998 ) ;
  assign n9000 = ~n1841 & n7341 ;
  assign n9001 = n1792 & n7644 ;
  assign n9002 = n9000 | n9001 ;
  assign n9003 = n1687 & n7345 ;
  assign n9004 = n9002 | n9003 ;
  assign n9005 = n7346 | n9004 ;
  assign n9006 = ( n4331 & n9004 ) | ( n4331 & n9005 ) | ( n9004 & n9005 ) ;
  assign n9007 = x8 & ~n9006 ;
  assign n9008 = ~x8 & n9006 ;
  assign n9009 = n9007 | n9008 ;
  assign n9010 = ( n8997 & n8999 ) | ( n8997 & n9009 ) | ( n8999 & n9009 ) ;
  assign n9011 = n1687 & n7644 ;
  assign n9012 = n1792 & n7341 ;
  assign n9013 = n1600 & n7345 ;
  assign n9014 = n9012 | n9013 ;
  assign n9015 = n9011 | n9014 ;
  assign n9016 = n7346 | n9015 ;
  assign n9017 = ( n4674 & n9015 ) | ( n4674 & n9016 ) | ( n9015 & n9016 ) ;
  assign n9018 = x8 & ~n9017 ;
  assign n9019 = ~x8 & n9017 ;
  assign n9020 = n9018 | n9019 ;
  assign n9021 = ( ~n8361 & n8371 ) | ( ~n8361 & n8597 ) | ( n8371 & n8597 ) ;
  assign n9022 = ( n8361 & ~n8598 ) | ( n8361 & n9021 ) | ( ~n8598 & n9021 ) ;
  assign n9023 = ( n9010 & n9020 ) | ( n9010 & n9022 ) | ( n9020 & n9022 ) ;
  assign n9024 = ( ~n8598 & n8608 ) | ( ~n8598 & n8610 ) | ( n8608 & n8610 ) ;
  assign n9025 = ( n8598 & ~n8611 ) | ( n8598 & n9024 ) | ( ~n8611 & n9024 ) ;
  assign n9026 = ~n1529 & n7345 ;
  assign n9027 = n1687 & n7341 ;
  assign n9028 = n9026 | n9027 ;
  assign n9029 = n1600 & n7644 ;
  assign n9030 = n9028 | n9029 ;
  assign n9031 = n7346 | n9030 ;
  assign n9032 = ( ~n4531 & n9030 ) | ( ~n4531 & n9031 ) | ( n9030 & n9031 ) ;
  assign n9033 = x8 & ~n9032 ;
  assign n9034 = ~x8 & n9032 ;
  assign n9035 = n9033 | n9034 ;
  assign n9036 = ( n9023 & n9025 ) | ( n9023 & n9035 ) | ( n9025 & n9035 ) ;
  assign n9037 = ( ~n8611 & n8613 ) | ( ~n8611 & n8623 ) | ( n8613 & n8623 ) ;
  assign n9038 = ( n8611 & ~n8624 ) | ( n8611 & n9037 ) | ( ~n8624 & n9037 ) ;
  assign n9039 = ~n1529 & n7644 ;
  assign n9040 = n1600 & n7341 ;
  assign n9041 = n1398 & n7345 ;
  assign n9042 = n9040 | n9041 ;
  assign n9043 = n9039 | n9042 ;
  assign n9044 = n7346 | n9043 ;
  assign n9045 = ( ~n4324 & n9043 ) | ( ~n4324 & n9044 ) | ( n9043 & n9044 ) ;
  assign n9046 = x8 & ~n9045 ;
  assign n9047 = ~x8 & n9045 ;
  assign n9048 = n9046 | n9047 ;
  assign n9049 = ( n9036 & n9038 ) | ( n9036 & n9048 ) | ( n9038 & n9048 ) ;
  assign n9050 = ( ~n8624 & n8626 ) | ( ~n8624 & n8636 ) | ( n8626 & n8636 ) ;
  assign n9051 = ( n8624 & ~n8637 ) | ( n8624 & n9050 ) | ( ~n8637 & n9050 ) ;
  assign n9052 = n1398 & n7644 ;
  assign n9053 = n7345 | n9052 ;
  assign n9054 = ( n1316 & n9052 ) | ( n1316 & n9053 ) | ( n9052 & n9053 ) ;
  assign n9055 = ~n1529 & n7341 ;
  assign n9056 = n9054 | n9055 ;
  assign n9057 = n7346 | n9056 ;
  assign n9058 = ( n4084 & n9056 ) | ( n4084 & n9057 ) | ( n9056 & n9057 ) ;
  assign n9059 = x8 & ~n9058 ;
  assign n9060 = ~x8 & n9058 ;
  assign n9061 = n9059 | n9060 ;
  assign n9062 = ( n9049 & n9051 ) | ( n9049 & n9061 ) | ( n9051 & n9061 ) ;
  assign n9063 = n1316 & n7644 ;
  assign n9064 = ~n1207 & n7345 ;
  assign n9065 = n1398 & n7341 ;
  assign n9066 = n9064 | n9065 ;
  assign n9067 = n9063 | n9066 ;
  assign n9068 = n7346 | n9067 ;
  assign n9069 = ( ~n4157 & n9067 ) | ( ~n4157 & n9068 ) | ( n9067 & n9068 ) ;
  assign n9070 = x8 & ~n9069 ;
  assign n9071 = ~x8 & n9069 ;
  assign n9072 = n9070 | n9071 ;
  assign n9073 = ( n8359 & n8637 ) | ( n8359 & n8639 ) | ( n8637 & n8639 ) ;
  assign n9074 = ( n8639 & n8640 ) | ( n8639 & ~n9073 ) | ( n8640 & ~n9073 ) ;
  assign n9075 = ( n9062 & n9072 ) | ( n9062 & ~n9074 ) | ( n9072 & ~n9074 ) ;
  assign n9076 = ~n1118 & n7345 ;
  assign n9077 = n1316 & n7341 ;
  assign n9078 = n9076 | n9077 ;
  assign n9079 = ~n1207 & n7644 ;
  assign n9080 = n9078 | n9079 ;
  assign n9081 = n7346 | n9080 ;
  assign n9082 = ( n3841 & n9080 ) | ( n3841 & n9081 ) | ( n9080 & n9081 ) ;
  assign n9083 = x8 & ~n9082 ;
  assign n9084 = ~x8 & n9082 ;
  assign n9085 = n9083 | n9084 ;
  assign n9086 = ( n8640 & n8650 ) | ( n8640 & n8652 ) | ( n8650 & n8652 ) ;
  assign n9087 = ( n8652 & n8653 ) | ( n8652 & ~n9086 ) | ( n8653 & ~n9086 ) ;
  assign n9088 = ( n9075 & n9085 ) | ( n9075 & ~n9087 ) | ( n9085 & ~n9087 ) ;
  assign n9089 = ( ~n8653 & n8655 ) | ( ~n8653 & n8665 ) | ( n8655 & n8665 ) ;
  assign n9090 = ( n8653 & ~n8666 ) | ( n8653 & n9089 ) | ( ~n8666 & n9089 ) ;
  assign n9091 = n995 & n7345 ;
  assign n9092 = ~n1207 & n7341 ;
  assign n9093 = n9091 | n9092 ;
  assign n9094 = ~n1118 & n7644 ;
  assign n9095 = n9093 | n9094 ;
  assign n9096 = n7346 | n9095 ;
  assign n9097 = ( n4173 & n9095 ) | ( n4173 & n9096 ) | ( n9095 & n9096 ) ;
  assign n9098 = x8 & ~n9097 ;
  assign n9099 = ~x8 & n9097 ;
  assign n9100 = n9098 | n9099 ;
  assign n9101 = ( n9088 & n9090 ) | ( n9088 & n9100 ) | ( n9090 & n9100 ) ;
  assign n9102 = ( n8666 & ~n8676 ) | ( n8666 & n8678 ) | ( ~n8676 & n8678 ) ;
  assign n9103 = ( ~n8666 & n8679 ) | ( ~n8666 & n9102 ) | ( n8679 & n9102 ) ;
  assign n9104 = n859 & n7345 ;
  assign n9105 = n995 & n7644 ;
  assign n9106 = n9104 | n9105 ;
  assign n9107 = ~n1118 & n7341 ;
  assign n9108 = n9106 | n9107 ;
  assign n9109 = n7346 | n9108 ;
  assign n9110 = ( ~n4034 & n9108 ) | ( ~n4034 & n9109 ) | ( n9108 & n9109 ) ;
  assign n9111 = x8 & ~n9110 ;
  assign n9112 = ~x8 & n9110 ;
  assign n9113 = n9111 | n9112 ;
  assign n9114 = ( n9101 & ~n9103 ) | ( n9101 & n9113 ) | ( ~n9103 & n9113 ) ;
  assign n9115 = ( ~n8679 & n8681 ) | ( ~n8679 & n8691 ) | ( n8681 & n8691 ) ;
  assign n9116 = ( n8679 & ~n8692 ) | ( n8679 & n9115 ) | ( ~n8692 & n9115 ) ;
  assign n9117 = n859 & n7644 ;
  assign n9118 = ~n721 & n7345 ;
  assign n9119 = n9117 | n9118 ;
  assign n9120 = n995 & n7341 ;
  assign n9121 = n9119 | n9120 ;
  assign n9122 = n7346 | n9121 ;
  assign n9123 = ( ~n3829 & n9121 ) | ( ~n3829 & n9122 ) | ( n9121 & n9122 ) ;
  assign n9124 = x8 & ~n9123 ;
  assign n9125 = ~x8 & n9123 ;
  assign n9126 = n9124 | n9125 ;
  assign n9127 = ( n9114 & n9116 ) | ( n9114 & n9126 ) | ( n9116 & n9126 ) ;
  assign n9128 = ( ~n8692 & n8702 ) | ( ~n8692 & n8704 ) | ( n8702 & n8704 ) ;
  assign n9129 = ( n8692 & ~n8705 ) | ( n8692 & n9128 ) | ( ~n8705 & n9128 ) ;
  assign n9130 = n564 & n7345 ;
  assign n9131 = n859 & n7341 ;
  assign n9132 = n9130 | n9131 ;
  assign n9133 = ~n721 & n7644 ;
  assign n9134 = n9132 | n9133 ;
  assign n9135 = n7346 | n9134 ;
  assign n9136 = ( ~n3268 & n9134 ) | ( ~n3268 & n9135 ) | ( n9134 & n9135 ) ;
  assign n9137 = x8 & ~n9136 ;
  assign n9138 = ~x8 & n9136 ;
  assign n9139 = n9137 | n9138 ;
  assign n9140 = ( n9127 & n9129 ) | ( n9127 & n9139 ) | ( n9129 & n9139 ) ;
  assign n9141 = ( n8732 & n8742 ) | ( n8732 & n9140 ) | ( n8742 & n9140 ) ;
  assign n9142 = ( ~n9127 & n9129 ) | ( ~n9127 & n9139 ) | ( n9129 & n9139 ) ;
  assign n9143 = ( n9127 & ~n9140 ) | ( n9127 & n9142 ) | ( ~n9140 & n9142 ) ;
  assign n9144 = ~n3487 & n8340 ;
  assign n9145 = x5 & n9144 ;
  assign n9146 = ~n3601 & n8721 ;
  assign n9147 = n40 & ~n3533 ;
  assign n9148 = n9146 | n9147 ;
  assign n9149 = n8341 | n9148 ;
  assign n9150 = ( ~n4223 & n9148 ) | ( ~n4223 & n9149 ) | ( n9148 & n9149 ) ;
  assign n9151 = x5 & ~n9150 ;
  assign n9152 = ( ~x5 & n9144 ) | ( ~x5 & n9150 ) | ( n9144 & n9150 ) ;
  assign n9153 = ( ~n9145 & n9151 ) | ( ~n9145 & n9152 ) | ( n9151 & n9152 ) ;
  assign n9154 = x0 | x1 ;
  assign n9155 = x2 & n9154 ;
  assign n9156 = ( x2 & n3516 ) | ( x2 & n9155 ) | ( n3516 & n9155 ) ;
  assign n9157 = n3607 & n9156 ;
  assign n9158 = x0 & x1 ;
  assign n9159 = x1 & x2 ;
  assign n9160 = n9158 | n9159 ;
  assign n9161 = ~n3607 & n9160 ;
  assign n9162 = n9157 | n9161 ;
  assign n9163 = ( n9143 & n9153 ) | ( n9143 & n9162 ) | ( n9153 & n9162 ) ;
  assign n9164 = n3123 & n8340 ;
  assign n9165 = x5 & n9164 ;
  assign n9166 = n40 & ~n2944 ;
  assign n9167 = ~n2977 & n8721 ;
  assign n9168 = n9166 | n9167 ;
  assign n9169 = n8341 | n9168 ;
  assign n9170 = ( ~n5926 & n9168 ) | ( ~n5926 & n9169 ) | ( n9168 & n9169 ) ;
  assign n9171 = x5 & ~n9170 ;
  assign n9172 = ( ~x5 & n9164 ) | ( ~x5 & n9170 ) | ( n9164 & n9170 ) ;
  assign n9173 = ( ~n9165 & n9171 ) | ( ~n9165 & n9172 ) | ( n9171 & n9172 ) ;
  assign n9174 = x8 & n8774 ;
  assign n9175 = ~n8773 & n9174 ;
  assign n9176 = n8773 & ~n9174 ;
  assign n9177 = n9175 | n9176 ;
  assign n9178 = n40 & ~n2977 ;
  assign n9179 = ~n3049 & n8340 ;
  assign n9180 = n9178 | n9179 ;
  assign n9181 = n3123 & n8721 ;
  assign n9182 = n9180 | n9181 ;
  assign n9183 = n8341 | n9182 ;
  assign n9184 = ( n6000 & n9182 ) | ( n6000 & n9183 ) | ( n9182 & n9183 ) ;
  assign n9185 = x5 & ~n9184 ;
  assign n9186 = ~x5 & n9184 ;
  assign n9187 = n9185 | n9186 ;
  assign n9188 = n40 & n3123 ;
  assign n9189 = ~n3049 & n8721 ;
  assign n9190 = n9188 | n9189 ;
  assign n9191 = n8341 | n9190 ;
  assign n9192 = ( n5965 & n9190 ) | ( n5965 & n9191 ) | ( n9190 & n9191 ) ;
  assign n9193 = ~n3232 & n8340 ;
  assign n9194 = n9192 | n9193 ;
  assign n9195 = n36 & ~n3049 ;
  assign n9196 = x5 & ~n8339 ;
  assign n9197 = ( x5 & n3232 ) | ( x5 & n9196 ) | ( n3232 & n9196 ) ;
  assign n9198 = ~n9195 & n9197 ;
  assign n9199 = ~n9194 & n9198 ;
  assign n9200 = ( n8774 & n9187 ) | ( n8774 & ~n9199 ) | ( n9187 & ~n9199 ) ;
  assign n9201 = n8774 & ~n9199 ;
  assign n9202 = ( n8774 & ~n9187 ) | ( n8774 & n9199 ) | ( ~n9187 & n9199 ) ;
  assign n9203 = ( n9200 & ~n9201 ) | ( n9200 & n9202 ) | ( ~n9201 & n9202 ) ;
  assign n9204 = ( n8774 & n9187 ) | ( n8774 & ~n9203 ) | ( n9187 & ~n9203 ) ;
  assign n9205 = ( n9173 & n9177 ) | ( n9173 & n9204 ) | ( n9177 & n9204 ) ;
  assign n9206 = n40 & ~n2888 ;
  assign n9207 = ~n2977 & n8340 ;
  assign n9208 = ~n2944 & n8721 ;
  assign n9209 = n9207 | n9208 ;
  assign n9210 = n9206 | n9209 ;
  assign n9211 = n8341 | n9210 ;
  assign n9212 = ( ~n6055 & n9210 ) | ( ~n6055 & n9211 ) | ( n9210 & n9211 ) ;
  assign n9213 = x5 & ~n9212 ;
  assign n9214 = ~x5 & n9212 ;
  assign n9215 = n9213 | n9214 ;
  assign n9216 = x8 & ~n8776 ;
  assign n9217 = ~n8783 & n9216 ;
  assign n9218 = n8783 & ~n9216 ;
  assign n9219 = n9217 | n9218 ;
  assign n9220 = ( n9205 & n9215 ) | ( n9205 & n9219 ) | ( n9215 & n9219 ) ;
  assign n9221 = ~n2888 & n8721 ;
  assign n9222 = ~n2944 & n8340 ;
  assign n9223 = n40 & n2820 ;
  assign n9224 = n9222 | n9223 ;
  assign n9225 = n9221 | n9224 ;
  assign n9226 = n8341 | n9225 ;
  assign n9227 = ( n6106 & n9225 ) | ( n6106 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9228 = x5 & ~n9227 ;
  assign n9229 = ~x5 & n9227 ;
  assign n9230 = n9228 | n9229 ;
  assign n9231 = ( n8395 & n8766 ) | ( n8395 & ~n8784 ) | ( n8766 & ~n8784 ) ;
  assign n9232 = ( n8395 & ~n8766 ) | ( n8395 & n8784 ) | ( ~n8766 & n8784 ) ;
  assign n9233 = ( ~n8785 & n9231 ) | ( ~n8785 & n9232 ) | ( n9231 & n9232 ) ;
  assign n9234 = ( n9220 & n9230 ) | ( n9220 & n9233 ) | ( n9230 & n9233 ) ;
  assign n9235 = ~n2888 & n8340 ;
  assign n9236 = x5 & n9235 ;
  assign n9237 = n40 & n2735 ;
  assign n9238 = n2820 & n8721 ;
  assign n9239 = n9237 | n9238 ;
  assign n9240 = n8341 | n9239 ;
  assign n9241 = ( ~n6157 & n9239 ) | ( ~n6157 & n9240 ) | ( n9239 & n9240 ) ;
  assign n9242 = x5 & ~n9241 ;
  assign n9243 = ( ~x5 & n9235 ) | ( ~x5 & n9241 ) | ( n9235 & n9241 ) ;
  assign n9244 = ( ~n9236 & n9242 ) | ( ~n9236 & n9243 ) | ( n9242 & n9243 ) ;
  assign n9245 = ( ~n8752 & n8756 ) | ( ~n8752 & n8786 ) | ( n8756 & n8786 ) ;
  assign n9246 = ( n8752 & ~n8787 ) | ( n8752 & n9245 ) | ( ~n8787 & n9245 ) ;
  assign n9247 = ( n9234 & n9244 ) | ( n9234 & n9246 ) | ( n9244 & n9246 ) ;
  assign n9248 = ( ~n8787 & n8797 ) | ( ~n8787 & n8801 ) | ( n8797 & n8801 ) ;
  assign n9249 = ( n8787 & ~n8802 ) | ( n8787 & n9248 ) | ( ~n8802 & n9248 ) ;
  assign n9250 = n2820 & n8340 ;
  assign n9251 = x5 & n9250 ;
  assign n9252 = n2735 & n8721 ;
  assign n9253 = n40 & n2642 ;
  assign n9254 = n9252 | n9253 ;
  assign n9255 = n8341 | n9254 ;
  assign n9256 = ( n5598 & n9254 ) | ( n5598 & n9255 ) | ( n9254 & n9255 ) ;
  assign n9257 = x5 & ~n9256 ;
  assign n9258 = ( ~x5 & n9250 ) | ( ~x5 & n9256 ) | ( n9250 & n9256 ) ;
  assign n9259 = ( ~n9251 & n9257 ) | ( ~n9251 & n9258 ) | ( n9257 & n9258 ) ;
  assign n9260 = ( n9247 & n9249 ) | ( n9247 & n9259 ) | ( n9249 & n9259 ) ;
  assign n9261 = ( ~n8802 & n8812 ) | ( ~n8802 & n8814 ) | ( n8812 & n8814 ) ;
  assign n9262 = ( n8802 & ~n8815 ) | ( n8802 & n9261 ) | ( ~n8815 & n9261 ) ;
  assign n9263 = n2735 & n8340 ;
  assign n9264 = n40 & ~n2608 ;
  assign n9265 = n2642 & n8721 ;
  assign n9266 = n9264 | n9265 ;
  assign n9267 = n9263 | n9266 ;
  assign n9268 = n8341 | n9267 ;
  assign n9269 = ( ~n6216 & n9267 ) | ( ~n6216 & n9268 ) | ( n9267 & n9268 ) ;
  assign n9270 = x5 & ~n9269 ;
  assign n9271 = ~x5 & n9269 ;
  assign n9272 = n9270 | n9271 ;
  assign n9273 = ( n9260 & n9262 ) | ( n9260 & n9272 ) | ( n9262 & n9272 ) ;
  assign n9274 = ( ~n8815 & n8825 ) | ( ~n8815 & n8827 ) | ( n8825 & n8827 ) ;
  assign n9275 = ( n8815 & ~n8828 ) | ( n8815 & n9274 ) | ( ~n8828 & n9274 ) ;
  assign n9276 = n2642 & n8340 ;
  assign n9277 = ~n2608 & n8721 ;
  assign n9278 = n9276 | n9277 ;
  assign n9279 = n40 & ~n2521 ;
  assign n9280 = n9278 | n9279 ;
  assign n9281 = n8341 | n9280 ;
  assign n9282 = ( n6221 & n9280 ) | ( n6221 & n9281 ) | ( n9280 & n9281 ) ;
  assign n9283 = x5 & ~n9282 ;
  assign n9284 = ~x5 & n9282 ;
  assign n9285 = n9283 | n9284 ;
  assign n9286 = ( n9273 & n9275 ) | ( n9273 & n9285 ) | ( n9275 & n9285 ) ;
  assign n9287 = ( ~n8828 & n8830 ) | ( ~n8828 & n8840 ) | ( n8830 & n8840 ) ;
  assign n9288 = ( n8828 & ~n8841 ) | ( n8828 & n9287 ) | ( ~n8841 & n9287 ) ;
  assign n9289 = ~n2608 & n8340 ;
  assign n9290 = x5 & n9289 ;
  assign n9291 = n40 & ~n2467 ;
  assign n9292 = ~n2521 & n8721 ;
  assign n9293 = n9291 | n9292 ;
  assign n9294 = n8341 | n9293 ;
  assign n9295 = ( ~n5693 & n9293 ) | ( ~n5693 & n9294 ) | ( n9293 & n9294 ) ;
  assign n9296 = x5 & ~n9295 ;
  assign n9297 = ( ~x5 & n9289 ) | ( ~x5 & n9295 ) | ( n9289 & n9295 ) ;
  assign n9298 = ( ~n9290 & n9296 ) | ( ~n9290 & n9297 ) | ( n9296 & n9297 ) ;
  assign n9299 = ( n9286 & n9288 ) | ( n9286 & n9298 ) | ( n9288 & n9298 ) ;
  assign n9300 = ( ~n8841 & n8851 ) | ( ~n8841 & n8853 ) | ( n8851 & n8853 ) ;
  assign n9301 = ( n8841 & ~n8854 ) | ( n8841 & n9300 ) | ( ~n8854 & n9300 ) ;
  assign n9302 = ~n2521 & n8340 ;
  assign n9303 = x5 & n9302 ;
  assign n9304 = ~n2467 & n8721 ;
  assign n9305 = n40 & n2398 ;
  assign n9306 = n9304 | n9305 ;
  assign n9307 = n8341 | n9306 ;
  assign n9308 = ( n5452 & n9306 ) | ( n5452 & n9307 ) | ( n9306 & n9307 ) ;
  assign n9309 = x5 & ~n9308 ;
  assign n9310 = ( ~x5 & n9302 ) | ( ~x5 & n9308 ) | ( n9302 & n9308 ) ;
  assign n9311 = ( ~n9303 & n9309 ) | ( ~n9303 & n9310 ) | ( n9309 & n9310 ) ;
  assign n9312 = ( n9299 & n9301 ) | ( n9299 & n9311 ) | ( n9301 & n9311 ) ;
  assign n9313 = ( ~n8854 & n8864 ) | ( ~n8854 & n8866 ) | ( n8864 & n8866 ) ;
  assign n9314 = ( n8854 & ~n8867 ) | ( n8854 & n9313 ) | ( ~n8867 & n9313 ) ;
  assign n9315 = n40 & ~n2364 ;
  assign n9316 = n2398 & n8721 ;
  assign n9317 = n9315 | n9316 ;
  assign n9318 = ~n2467 & n8340 ;
  assign n9319 = n9317 | n9318 ;
  assign n9320 = n8341 | n9319 ;
  assign n9321 = ( n5713 & n9319 ) | ( n5713 & n9320 ) | ( n9319 & n9320 ) ;
  assign n9322 = x5 & ~n9321 ;
  assign n9323 = ~x5 & n9321 ;
  assign n9324 = n9322 | n9323 ;
  assign n9325 = ( n9312 & n9314 ) | ( n9312 & n9324 ) | ( n9314 & n9324 ) ;
  assign n9326 = ( ~n8867 & n8869 ) | ( ~n8867 & n8879 ) | ( n8869 & n8879 ) ;
  assign n9327 = ( n8867 & ~n8880 ) | ( n8867 & n9326 ) | ( ~n8880 & n9326 ) ;
  assign n9328 = n2398 & n8340 ;
  assign n9329 = x5 & n9328 ;
  assign n9330 = ~n2364 & n8721 ;
  assign n9331 = n40 & ~n2282 ;
  assign n9332 = n9330 | n9331 ;
  assign n9333 = n8341 | n9332 ;
  assign n9334 = ( ~n5494 & n9332 ) | ( ~n5494 & n9333 ) | ( n9332 & n9333 ) ;
  assign n9335 = x5 & ~n9334 ;
  assign n9336 = ( ~x5 & n9328 ) | ( ~x5 & n9334 ) | ( n9328 & n9334 ) ;
  assign n9337 = ( ~n9329 & n9335 ) | ( ~n9329 & n9336 ) | ( n9335 & n9336 ) ;
  assign n9338 = ( n9325 & n9327 ) | ( n9325 & n9337 ) | ( n9327 & n9337 ) ;
  assign n9339 = ( ~n8880 & n8882 ) | ( ~n8880 & n8892 ) | ( n8882 & n8892 ) ;
  assign n9340 = ( n8880 & ~n8893 ) | ( n8880 & n9339 ) | ( ~n8893 & n9339 ) ;
  assign n9341 = ~n2364 & n8340 ;
  assign n9342 = n40 & n2187 ;
  assign n9343 = n9341 | n9342 ;
  assign n9344 = ~n2282 & n8721 ;
  assign n9345 = n9343 | n9344 ;
  assign n9346 = n8341 | n9345 ;
  assign n9347 = ( n5137 & n9345 ) | ( n5137 & n9346 ) | ( n9345 & n9346 ) ;
  assign n9348 = x5 & ~n9347 ;
  assign n9349 = ~x5 & n9347 ;
  assign n9350 = n9348 | n9349 ;
  assign n9351 = ( n9338 & n9340 ) | ( n9338 & n9350 ) | ( n9340 & n9350 ) ;
  assign n9352 = ( ~n8893 & n8895 ) | ( ~n8893 & n8905 ) | ( n8895 & n8905 ) ;
  assign n9353 = ( n8893 & ~n8906 ) | ( n8893 & n9352 ) | ( ~n8906 & n9352 ) ;
  assign n9354 = ~n2282 & n8340 ;
  assign n9355 = x5 & n9354 ;
  assign n9356 = n40 & n2102 ;
  assign n9357 = n2187 & n8721 ;
  assign n9358 = n9356 | n9357 ;
  assign n9359 = n8341 | n9358 ;
  assign n9360 = ( ~n5331 & n9358 ) | ( ~n5331 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9361 = x5 & ~n9360 ;
  assign n9362 = ( ~x5 & n9354 ) | ( ~x5 & n9360 ) | ( n9354 & n9360 ) ;
  assign n9363 = ( ~n9355 & n9361 ) | ( ~n9355 & n9362 ) | ( n9361 & n9362 ) ;
  assign n9364 = ( n9351 & n9353 ) | ( n9351 & n9363 ) | ( n9353 & n9363 ) ;
  assign n9365 = ( ~n8906 & n8908 ) | ( ~n8906 & n8918 ) | ( n8908 & n8918 ) ;
  assign n9366 = ( n8906 & ~n8919 ) | ( n8906 & n9365 ) | ( ~n8919 & n9365 ) ;
  assign n9367 = n40 & ~n2041 ;
  assign n9368 = n8341 | n9367 ;
  assign n9369 = ( ~n4997 & n9367 ) | ( ~n4997 & n9368 ) | ( n9367 & n9368 ) ;
  assign n9370 = n2187 & n8340 ;
  assign n9371 = ( ~x5 & n9369 ) | ( ~x5 & n9370 ) | ( n9369 & n9370 ) ;
  assign n9372 = n2102 & n8721 ;
  assign n9373 = x5 & ~n9370 ;
  assign n9374 = n9372 | n9373 ;
  assign n9375 = ( n9369 & n9372 ) | ( n9369 & n9373 ) | ( n9372 & n9373 ) ;
  assign n9376 = ( n9371 & n9374 ) | ( n9371 & ~n9375 ) | ( n9374 & ~n9375 ) ;
  assign n9377 = ( n9364 & n9366 ) | ( n9364 & n9376 ) | ( n9366 & n9376 ) ;
  assign n9378 = ( ~n8919 & n8921 ) | ( ~n8919 & n8931 ) | ( n8921 & n8931 ) ;
  assign n9379 = ( n8919 & ~n8932 ) | ( n8919 & n9378 ) | ( ~n8932 & n9378 ) ;
  assign n9380 = n40 & n1943 ;
  assign n9381 = n2102 & n8340 ;
  assign n9382 = n9380 | n9381 ;
  assign n9383 = ~n2041 & n8721 ;
  assign n9384 = n9382 | n9383 ;
  assign n9385 = n8341 | n9384 ;
  assign n9386 = ( ~n4985 & n9384 ) | ( ~n4985 & n9385 ) | ( n9384 & n9385 ) ;
  assign n9387 = x5 & ~n9386 ;
  assign n9388 = ~x5 & n9386 ;
  assign n9389 = n9387 | n9388 ;
  assign n9390 = ( n9377 & n9379 ) | ( n9377 & n9389 ) | ( n9379 & n9389 ) ;
  assign n9391 = ( ~n8932 & n8934 ) | ( ~n8932 & n8944 ) | ( n8934 & n8944 ) ;
  assign n9392 = ( n8932 & ~n8945 ) | ( n8932 & n9391 ) | ( ~n8945 & n9391 ) ;
  assign n9393 = n40 & ~n1841 ;
  assign n9394 = n8341 | n9393 ;
  assign n9395 = ( ~n4753 & n9393 ) | ( ~n4753 & n9394 ) | ( n9393 & n9394 ) ;
  assign n9396 = ~n2041 & n8340 ;
  assign n9397 = ( ~x5 & n9395 ) | ( ~x5 & n9396 ) | ( n9395 & n9396 ) ;
  assign n9398 = n1943 & n8721 ;
  assign n9399 = x5 & ~n9396 ;
  assign n9400 = n9398 | n9399 ;
  assign n9401 = ( n9395 & n9398 ) | ( n9395 & n9399 ) | ( n9398 & n9399 ) ;
  assign n9402 = ( n9397 & n9400 ) | ( n9397 & ~n9401 ) | ( n9400 & ~n9401 ) ;
  assign n9403 = ( n9390 & n9392 ) | ( n9390 & n9402 ) | ( n9392 & n9402 ) ;
  assign n9404 = ( ~n8945 & n8947 ) | ( ~n8945 & n8957 ) | ( n8947 & n8957 ) ;
  assign n9405 = ( n8945 & ~n8958 ) | ( n8945 & n9404 ) | ( ~n8958 & n9404 ) ;
  assign n9406 = n1943 & n8340 ;
  assign n9407 = n40 & n1792 ;
  assign n9408 = n9406 | n9407 ;
  assign n9409 = ~n1841 & n8721 ;
  assign n9410 = n9408 | n9409 ;
  assign n9411 = n8341 | n9410 ;
  assign n9412 = ( ~n4831 & n9410 ) | ( ~n4831 & n9411 ) | ( n9410 & n9411 ) ;
  assign n9413 = x5 & ~n9412 ;
  assign n9414 = ~x5 & n9412 ;
  assign n9415 = n9413 | n9414 ;
  assign n9416 = ( n9403 & n9405 ) | ( n9403 & n9415 ) | ( n9405 & n9415 ) ;
  assign n9417 = ( ~n8958 & n8960 ) | ( ~n8958 & n8970 ) | ( n8960 & n8970 ) ;
  assign n9418 = ( n8958 & ~n8971 ) | ( n8958 & n9417 ) | ( ~n8971 & n9417 ) ;
  assign n9419 = ~n1841 & n8340 ;
  assign n9420 = n40 & n1687 ;
  assign n9421 = n9419 | n9420 ;
  assign n9422 = n1792 & n8721 ;
  assign n9423 = n9421 | n9422 ;
  assign n9424 = n8341 | n9423 ;
  assign n9425 = ( n4331 & n9423 ) | ( n4331 & n9424 ) | ( n9423 & n9424 ) ;
  assign n9426 = x5 & ~n9425 ;
  assign n9427 = ~x5 & n9425 ;
  assign n9428 = n9426 | n9427 ;
  assign n9429 = ( n9416 & n9418 ) | ( n9416 & n9428 ) | ( n9418 & n9428 ) ;
  assign n9430 = ( ~n8971 & n8973 ) | ( ~n8971 & n8983 ) | ( n8973 & n8983 ) ;
  assign n9431 = ( n8971 & ~n8984 ) | ( n8971 & n9430 ) | ( ~n8984 & n9430 ) ;
  assign n9432 = n1687 & n8721 ;
  assign n9433 = n1792 & n8340 ;
  assign n9434 = n40 & n1600 ;
  assign n9435 = n9433 | n9434 ;
  assign n9436 = n9432 | n9435 ;
  assign n9437 = n8341 | n9436 ;
  assign n9438 = ( n4674 & n9436 ) | ( n4674 & n9437 ) | ( n9436 & n9437 ) ;
  assign n9439 = x5 & ~n9438 ;
  assign n9440 = ~x5 & n9438 ;
  assign n9441 = n9439 | n9440 ;
  assign n9442 = ( n9429 & n9431 ) | ( n9429 & n9441 ) | ( n9431 & n9441 ) ;
  assign n9443 = n40 & ~n1529 ;
  assign n9444 = n1687 & n8340 ;
  assign n9445 = n9443 | n9444 ;
  assign n9446 = n1600 & n8721 ;
  assign n9447 = n9445 | n9446 ;
  assign n9448 = n8341 | n9447 ;
  assign n9449 = ( ~n4531 & n9447 ) | ( ~n4531 & n9448 ) | ( n9447 & n9448 ) ;
  assign n9450 = x5 & ~n9449 ;
  assign n9451 = ~x5 & n9449 ;
  assign n9452 = n9450 | n9451 ;
  assign n9453 = ( ~n8984 & n8994 ) | ( ~n8984 & n8996 ) | ( n8994 & n8996 ) ;
  assign n9454 = ( n8984 & ~n8997 ) | ( n8984 & n9453 ) | ( ~n8997 & n9453 ) ;
  assign n9455 = ( n9442 & n9452 ) | ( n9442 & n9454 ) | ( n9452 & n9454 ) ;
  assign n9456 = ( ~n8997 & n8999 ) | ( ~n8997 & n9009 ) | ( n8999 & n9009 ) ;
  assign n9457 = ( n8997 & ~n9010 ) | ( n8997 & n9456 ) | ( ~n9010 & n9456 ) ;
  assign n9458 = ~n1529 & n8721 ;
  assign n9459 = n1600 & n8340 ;
  assign n9460 = n40 & n1398 ;
  assign n9461 = n9459 | n9460 ;
  assign n9462 = n9458 | n9461 ;
  assign n9463 = n8341 | n9462 ;
  assign n9464 = ( ~n4324 & n9462 ) | ( ~n4324 & n9463 ) | ( n9462 & n9463 ) ;
  assign n9465 = x5 & ~n9464 ;
  assign n9466 = ~x5 & n9464 ;
  assign n9467 = n9465 | n9466 ;
  assign n9468 = ( n9455 & n9457 ) | ( n9455 & n9467 ) | ( n9457 & n9467 ) ;
  assign n9469 = ( ~n9010 & n9020 ) | ( ~n9010 & n9022 ) | ( n9020 & n9022 ) ;
  assign n9470 = ( n9010 & ~n9023 ) | ( n9010 & n9469 ) | ( ~n9023 & n9469 ) ;
  assign n9471 = ~n1529 & n8340 ;
  assign n9472 = n40 & n1316 ;
  assign n9473 = n9471 | n9472 ;
  assign n9474 = n1398 & n8721 ;
  assign n9475 = n9473 | n9474 ;
  assign n9476 = n8341 | n9475 ;
  assign n9477 = ( n4084 & n9475 ) | ( n4084 & n9476 ) | ( n9475 & n9476 ) ;
  assign n9478 = x5 & ~n9477 ;
  assign n9479 = ~x5 & n9477 ;
  assign n9480 = n9478 | n9479 ;
  assign n9481 = ( n9468 & n9470 ) | ( n9468 & n9480 ) | ( n9470 & n9480 ) ;
  assign n9482 = ( ~n9023 & n9025 ) | ( ~n9023 & n9035 ) | ( n9025 & n9035 ) ;
  assign n9483 = ( n9023 & ~n9036 ) | ( n9023 & n9482 ) | ( ~n9036 & n9482 ) ;
  assign n9484 = n1398 & n8340 ;
  assign n9485 = x5 & n9484 ;
  assign n9486 = n1316 & n8721 ;
  assign n9487 = n40 & ~n1207 ;
  assign n9488 = n9486 | n9487 ;
  assign n9489 = n8341 | n9488 ;
  assign n9490 = ( ~n4157 & n9488 ) | ( ~n4157 & n9489 ) | ( n9488 & n9489 ) ;
  assign n9491 = x5 & ~n9490 ;
  assign n9492 = ( ~x5 & n9484 ) | ( ~x5 & n9490 ) | ( n9484 & n9490 ) ;
  assign n9493 = ( ~n9485 & n9491 ) | ( ~n9485 & n9492 ) | ( n9491 & n9492 ) ;
  assign n9494 = ( n9481 & n9483 ) | ( n9481 & n9493 ) | ( n9483 & n9493 ) ;
  assign n9495 = ( ~n9036 & n9038 ) | ( ~n9036 & n9048 ) | ( n9038 & n9048 ) ;
  assign n9496 = ( n9036 & ~n9049 ) | ( n9036 & n9495 ) | ( ~n9049 & n9495 ) ;
  assign n9497 = n1316 & n8340 ;
  assign n9498 = x5 & n9497 ;
  assign n9499 = n40 & ~n1118 ;
  assign n9500 = ~n1207 & n8721 ;
  assign n9501 = n9499 | n9500 ;
  assign n9502 = n8341 | n9501 ;
  assign n9503 = ( n3841 & n9501 ) | ( n3841 & n9502 ) | ( n9501 & n9502 ) ;
  assign n9504 = x5 & ~n9503 ;
  assign n9505 = ( ~x5 & n9497 ) | ( ~x5 & n9503 ) | ( n9497 & n9503 ) ;
  assign n9506 = ( ~n9498 & n9504 ) | ( ~n9498 & n9505 ) | ( n9504 & n9505 ) ;
  assign n9507 = ( n9494 & n9496 ) | ( n9494 & n9506 ) | ( n9496 & n9506 ) ;
  assign n9508 = ( ~n9049 & n9051 ) | ( ~n9049 & n9061 ) | ( n9051 & n9061 ) ;
  assign n9509 = ( n9049 & ~n9062 ) | ( n9049 & n9508 ) | ( ~n9062 & n9508 ) ;
  assign n9510 = n40 & n995 ;
  assign n9511 = ~n1207 & n8340 ;
  assign n9512 = n9510 | n9511 ;
  assign n9513 = ~n1118 & n8721 ;
  assign n9514 = n9512 | n9513 ;
  assign n9515 = n8341 | n9514 ;
  assign n9516 = ( n4173 & n9514 ) | ( n4173 & n9515 ) | ( n9514 & n9515 ) ;
  assign n9517 = x5 & ~n9516 ;
  assign n9518 = ~x5 & n9516 ;
  assign n9519 = n9517 | n9518 ;
  assign n9520 = ( n9507 & n9509 ) | ( n9507 & n9519 ) | ( n9509 & n9519 ) ;
  assign n9521 = ( n9062 & ~n9072 ) | ( n9062 & n9074 ) | ( ~n9072 & n9074 ) ;
  assign n9522 = ( ~n9062 & n9075 ) | ( ~n9062 & n9521 ) | ( n9075 & n9521 ) ;
  assign n9523 = n40 & n859 ;
  assign n9524 = n995 & n8721 ;
  assign n9525 = n9523 | n9524 ;
  assign n9526 = ~n1118 & n8340 ;
  assign n9527 = n9525 | n9526 ;
  assign n9528 = n8341 | n9527 ;
  assign n9529 = ( ~n4034 & n9527 ) | ( ~n4034 & n9528 ) | ( n9527 & n9528 ) ;
  assign n9530 = x5 & ~n9529 ;
  assign n9531 = ~x5 & n9529 ;
  assign n9532 = n9530 | n9531 ;
  assign n9533 = ( n9520 & ~n9522 ) | ( n9520 & n9532 ) | ( ~n9522 & n9532 ) ;
  assign n9534 = ( n9075 & ~n9085 ) | ( n9075 & n9087 ) | ( ~n9085 & n9087 ) ;
  assign n9535 = ( ~n9075 & n9088 ) | ( ~n9075 & n9534 ) | ( n9088 & n9534 ) ;
  assign n9536 = n859 & n8721 ;
  assign n9537 = n40 & ~n721 ;
  assign n9538 = n9536 | n9537 ;
  assign n9539 = n995 & n8340 ;
  assign n9540 = n9538 | n9539 ;
  assign n9541 = n8341 | n9540 ;
  assign n9542 = ( ~n3829 & n9540 ) | ( ~n3829 & n9541 ) | ( n9540 & n9541 ) ;
  assign n9543 = x5 & ~n9542 ;
  assign n9544 = ~x5 & n9542 ;
  assign n9545 = n9543 | n9544 ;
  assign n9546 = ( n9533 & ~n9535 ) | ( n9533 & n9545 ) | ( ~n9535 & n9545 ) ;
  assign n9547 = ( ~n9088 & n9090 ) | ( ~n9088 & n9100 ) | ( n9090 & n9100 ) ;
  assign n9548 = ( n9088 & ~n9101 ) | ( n9088 & n9547 ) | ( ~n9101 & n9547 ) ;
  assign n9549 = n859 & n8340 ;
  assign n9550 = x5 & n9549 ;
  assign n9551 = n40 & n564 ;
  assign n9552 = ~n721 & n8721 ;
  assign n9553 = n9551 | n9552 ;
  assign n9554 = n8341 | n9553 ;
  assign n9555 = ( ~n3268 & n9553 ) | ( ~n3268 & n9554 ) | ( n9553 & n9554 ) ;
  assign n9556 = x5 & ~n9555 ;
  assign n9557 = ( ~x5 & n9549 ) | ( ~x5 & n9555 ) | ( n9549 & n9555 ) ;
  assign n9558 = ( ~n9550 & n9556 ) | ( ~n9550 & n9557 ) | ( n9556 & n9557 ) ;
  assign n9559 = ( n9546 & n9548 ) | ( n9546 & n9558 ) | ( n9548 & n9558 ) ;
  assign n9560 = ( n9101 & n9103 ) | ( n9101 & ~n9113 ) | ( n9103 & ~n9113 ) ;
  assign n9561 = ( ~n9101 & n9114 ) | ( ~n9101 & n9560 ) | ( n9114 & n9560 ) ;
  assign n9562 = n40 & ~n3487 ;
  assign n9563 = ~n721 & n8340 ;
  assign n9564 = n564 & n8721 ;
  assign n9565 = n9563 | n9564 ;
  assign n9566 = n9562 | n9565 ;
  assign n9567 = n8341 | n9566 ;
  assign n9568 = ( ~n3492 & n9566 ) | ( ~n3492 & n9567 ) | ( n9566 & n9567 ) ;
  assign n9569 = x5 & ~n9568 ;
  assign n9570 = ~x5 & n9568 ;
  assign n9571 = n9569 | n9570 ;
  assign n9572 = ( n9559 & ~n9561 ) | ( n9559 & n9571 ) | ( ~n9561 & n9571 ) ;
  assign n9573 = ~n3487 & n8721 ;
  assign n9574 = n40 & ~n3601 ;
  assign n9575 = n564 & n8340 ;
  assign n9576 = n9574 | n9575 ;
  assign n9577 = n9573 | n9576 ;
  assign n9578 = n8341 | n9577 ;
  assign n9579 = ( n3674 & n9577 ) | ( n3674 & n9578 ) | ( n9577 & n9578 ) ;
  assign n9580 = x5 & ~n9579 ;
  assign n9581 = ~x5 & n9579 ;
  assign n9582 = n9580 | n9581 ;
  assign n9583 = ( ~n9114 & n9116 ) | ( ~n9114 & n9126 ) | ( n9116 & n9126 ) ;
  assign n9584 = ( n9114 & ~n9127 ) | ( n9114 & n9583 ) | ( ~n9127 & n9583 ) ;
  assign n9585 = ( n9572 & n9582 ) | ( n9572 & n9584 ) | ( n9582 & n9584 ) ;
  assign n9586 = ( ~n9364 & n9366 ) | ( ~n9364 & n9376 ) | ( n9366 & n9376 ) ;
  assign n9587 = ( n9364 & ~n9377 ) | ( n9364 & n9586 ) | ( ~n9377 & n9586 ) ;
  assign n9588 = x0 & ~x1 ;
  assign n9589 = x2 & n9588 ;
  assign n9590 = x2 & ~n9588 ;
  assign n9591 = n9158 & ~n9590 ;
  assign n9592 = n9589 | n9591 ;
  assign n9593 = x0 & ~n9592 ;
  assign n9594 = n1792 & n9593 ;
  assign n9595 = n9592 | n9594 ;
  assign n9596 = ( ~n4831 & n9594 ) | ( ~n4831 & n9595 ) | ( n9594 & n9595 ) ;
  assign n9597 = n41 & ~n1841 ;
  assign n9598 = ( x2 & ~n9596 ) | ( x2 & n9597 ) | ( ~n9596 & n9597 ) ;
  assign n9599 = ~x2 & n9596 ;
  assign n9600 = x2 & ~n9154 ;
  assign n9601 = n1943 & n9600 ;
  assign n9602 = ( x2 & n9597 ) | ( x2 & n9601 ) | ( n9597 & n9601 ) ;
  assign n9603 = ( n9598 & n9599 ) | ( n9598 & ~n9602 ) | ( n9599 & ~n9602 ) ;
  assign n9604 = ( ~n9338 & n9340 ) | ( ~n9338 & n9350 ) | ( n9340 & n9350 ) ;
  assign n9605 = ( n9338 & ~n9351 ) | ( n9338 & n9604 ) | ( ~n9351 & n9604 ) ;
  assign n9606 = n1943 & n9593 ;
  assign n9607 = n41 & ~n2041 ;
  assign n9608 = n9606 | n9607 ;
  assign n9609 = x2 & n9608 ;
  assign n9610 = ~x2 & n9608 ;
  assign n9611 = n2102 & n9600 ;
  assign n9612 = ( x2 & n4985 ) | ( x2 & n9590 ) | ( n4985 & n9590 ) ;
  assign n9613 = ~n4985 & n9591 ;
  assign n9614 = ( ~n9611 & n9612 ) | ( ~n9611 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9615 = ( ~n9609 & n9610 ) | ( ~n9609 & n9614 ) | ( n9610 & n9614 ) ;
  assign n9616 = ~n2944 & n9593 ;
  assign n9617 = n41 & ~n2977 ;
  assign n9618 = n9616 | n9617 ;
  assign n9619 = n9592 | n9618 ;
  assign n9620 = ( ~n5926 & n9618 ) | ( ~n5926 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9621 = x2 & n9620 ;
  assign n9622 = x2 & ~n3123 ;
  assign n9623 = n9155 | n9622 ;
  assign n9624 = n9620 | n9623 ;
  assign n9625 = ~n9621 & n9624 ;
  assign n9626 = ( x4 & n34 ) | ( x4 & n3232 ) | ( n34 & n3232 ) ;
  assign n9627 = ( n8337 & n9195 ) | ( n8337 & n9626 ) | ( n9195 & n9626 ) ;
  assign n9628 = ( n8337 & ~n9195 ) | ( n8337 & n9626 ) | ( ~n9195 & n9626 ) ;
  assign n9629 = ( n9195 & ~n9627 ) | ( n9195 & n9628 ) | ( ~n9627 & n9628 ) ;
  assign n9630 = ~n2977 & n9593 ;
  assign n9631 = ~n3049 & n9600 ;
  assign n9632 = n9630 | n9631 ;
  assign n9633 = n9592 | n9632 ;
  assign n9634 = ( n6000 & n9632 ) | ( n6000 & n9633 ) | ( n9632 & n9633 ) ;
  assign n9635 = n35 & ~n3232 ;
  assign n9636 = n9634 & ~n9635 ;
  assign n9637 = n41 & n3123 ;
  assign n9638 = ( n9634 & n9635 ) | ( n9634 & n9637 ) | ( n9635 & n9637 ) ;
  assign n9639 = ~x0 & x2 ;
  assign n9640 = n9622 | n9639 ;
  assign n9641 = n33 & ~n3232 ;
  assign n9642 = ~n3049 & n9154 ;
  assign n9643 = n3232 & ~n9642 ;
  assign n9644 = n9641 | n9643 ;
  assign n9645 = ( n9640 & n9641 ) | ( n9640 & n9644 ) | ( n9641 & n9644 ) ;
  assign n9646 = ~n9637 & n9645 ;
  assign n9647 = ( ~n9636 & n9638 ) | ( ~n9636 & n9646 ) | ( n9638 & n9646 ) ;
  assign n9648 = ( n9625 & n9629 ) | ( n9625 & n9647 ) | ( n9629 & n9647 ) ;
  assign n9649 = ~n2888 & n9593 ;
  assign n9650 = n41 & ~n2944 ;
  assign n9651 = n9649 | n9650 ;
  assign n9652 = n9592 | n9651 ;
  assign n9653 = ( ~n6055 & n9651 ) | ( ~n6055 & n9652 ) | ( n9651 & n9652 ) ;
  assign n9654 = ~x2 & n9653 ;
  assign n9655 = ( x2 & n2977 ) | ( x2 & n9155 ) | ( n2977 & n9155 ) ;
  assign n9656 = ~n9653 & n9655 ;
  assign n9657 = n9654 | n9656 ;
  assign n9658 = x5 & ~n9198 ;
  assign n9659 = ~n9194 & n9658 ;
  assign n9660 = n9194 & ~n9658 ;
  assign n9661 = n9659 | n9660 ;
  assign n9662 = ( n9648 & n9657 ) | ( n9648 & n9661 ) | ( n9657 & n9661 ) ;
  assign n9663 = n41 & ~n2888 ;
  assign n9664 = n2820 & n9593 ;
  assign n9665 = n9663 | n9664 ;
  assign n9666 = n9592 | n9665 ;
  assign n9667 = ( n6106 & n9665 ) | ( n6106 & n9666 ) | ( n9665 & n9666 ) ;
  assign n9668 = ~x2 & n9667 ;
  assign n9669 = ( x2 & n2944 ) | ( x2 & n9155 ) | ( n2944 & n9155 ) ;
  assign n9670 = ~n9667 & n9669 ;
  assign n9671 = n9668 | n9670 ;
  assign n9672 = ( n9203 & n9662 ) | ( n9203 & n9671 ) | ( n9662 & n9671 ) ;
  assign n9673 = n2735 & n9593 ;
  assign n9674 = n41 & n2820 ;
  assign n9675 = n9673 | n9674 ;
  assign n9676 = n9592 | n9675 ;
  assign n9677 = ( ~n6157 & n9675 ) | ( ~n6157 & n9676 ) | ( n9675 & n9676 ) ;
  assign n9678 = x2 & n9677 ;
  assign n9679 = ( x2 & n2888 ) | ( x2 & n9155 ) | ( n2888 & n9155 ) ;
  assign n9680 = n9677 | n9679 ;
  assign n9681 = ~n9678 & n9680 ;
  assign n9682 = ( ~n9173 & n9177 ) | ( ~n9173 & n9204 ) | ( n9177 & n9204 ) ;
  assign n9683 = ( n9173 & ~n9205 ) | ( n9173 & n9682 ) | ( ~n9205 & n9682 ) ;
  assign n9684 = ( n9672 & n9681 ) | ( n9672 & n9683 ) | ( n9681 & n9683 ) ;
  assign n9685 = ( ~n9205 & n9215 ) | ( ~n9205 & n9219 ) | ( n9215 & n9219 ) ;
  assign n9686 = ( n9205 & ~n9220 ) | ( n9205 & n9685 ) | ( ~n9220 & n9685 ) ;
  assign n9687 = n5598 & n9591 ;
  assign n9688 = ( x2 & ~n5598 ) | ( x2 & n9590 ) | ( ~n5598 & n9590 ) ;
  assign n9689 = n41 & n2735 ;
  assign n9690 = n2642 & n9593 ;
  assign n9691 = n9689 | n9690 ;
  assign n9692 = n2820 & n9600 ;
  assign n9693 = n9691 | n9692 ;
  assign n9694 = n9688 & n9693 ;
  assign n9695 = n9688 | n9691 ;
  assign n9696 = ( n9687 & ~n9694 ) | ( n9687 & n9695 ) | ( ~n9694 & n9695 ) ;
  assign n9697 = ( n9684 & n9686 ) | ( n9684 & n9696 ) | ( n9686 & n9696 ) ;
  assign n9698 = ( ~n9220 & n9230 ) | ( ~n9220 & n9233 ) | ( n9230 & n9233 ) ;
  assign n9699 = ( n9220 & ~n9234 ) | ( n9220 & n9698 ) | ( ~n9234 & n9698 ) ;
  assign n9700 = n2735 & n9600 ;
  assign n9701 = n41 & n2642 ;
  assign n9702 = ~n2608 & n9593 ;
  assign n9703 = n9701 | n9702 ;
  assign n9704 = n9700 | n9703 ;
  assign n9705 = n9592 | n9704 ;
  assign n9706 = ( ~n6216 & n9704 ) | ( ~n6216 & n9705 ) | ( n9704 & n9705 ) ;
  assign n9707 = x2 & ~n9706 ;
  assign n9708 = ~x2 & n9706 ;
  assign n9709 = n9707 | n9708 ;
  assign n9710 = ( n9697 & n9699 ) | ( n9697 & n9709 ) | ( n9699 & n9709 ) ;
  assign n9711 = ( ~n9234 & n9244 ) | ( ~n9234 & n9246 ) | ( n9244 & n9246 ) ;
  assign n9712 = ( n9234 & ~n9247 ) | ( n9234 & n9711 ) | ( ~n9247 & n9711 ) ;
  assign n9713 = ~n2521 & n9593 ;
  assign n9714 = n9592 | n9713 ;
  assign n9715 = ( n6221 & n9713 ) | ( n6221 & n9714 ) | ( n9713 & n9714 ) ;
  assign n9716 = n41 & ~n2608 ;
  assign n9717 = ( x2 & ~n9715 ) | ( x2 & n9716 ) | ( ~n9715 & n9716 ) ;
  assign n9718 = ~x2 & n9715 ;
  assign n9719 = n2642 & n9600 ;
  assign n9720 = ( x2 & n9716 ) | ( x2 & n9719 ) | ( n9716 & n9719 ) ;
  assign n9721 = ( n9717 & n9718 ) | ( n9717 & ~n9720 ) | ( n9718 & ~n9720 ) ;
  assign n9722 = ( n9710 & n9712 ) | ( n9710 & n9721 ) | ( n9712 & n9721 ) ;
  assign n9723 = ( ~n9247 & n9249 ) | ( ~n9247 & n9259 ) | ( n9249 & n9259 ) ;
  assign n9724 = ( n9247 & ~n9260 ) | ( n9247 & n9723 ) | ( ~n9260 & n9723 ) ;
  assign n9725 = ~n2467 & n9593 ;
  assign n9726 = n41 & ~n2521 ;
  assign n9727 = n9725 | n9726 ;
  assign n9728 = n9592 | n9727 ;
  assign n9729 = ( ~n5693 & n9727 ) | ( ~n5693 & n9728 ) | ( n9727 & n9728 ) ;
  assign n9730 = x2 & n9729 ;
  assign n9731 = ( x2 & n2608 ) | ( x2 & n9155 ) | ( n2608 & n9155 ) ;
  assign n9732 = n9729 | n9731 ;
  assign n9733 = ~n9730 & n9732 ;
  assign n9734 = ( n9722 & n9724 ) | ( n9722 & n9733 ) | ( n9724 & n9733 ) ;
  assign n9735 = n2398 & n9593 ;
  assign n9736 = x2 & n9735 ;
  assign n9737 = n41 & ~n2467 ;
  assign n9738 = ~n2521 & n9600 ;
  assign n9739 = n9737 | n9738 ;
  assign n9740 = n9592 | n9739 ;
  assign n9741 = ( n5452 & n9739 ) | ( n5452 & n9740 ) | ( n9739 & n9740 ) ;
  assign n9742 = x2 & ~n9741 ;
  assign n9743 = ( ~x2 & n9735 ) | ( ~x2 & n9741 ) | ( n9735 & n9741 ) ;
  assign n9744 = ( ~n9736 & n9742 ) | ( ~n9736 & n9743 ) | ( n9742 & n9743 ) ;
  assign n9745 = ( ~n9260 & n9262 ) | ( ~n9260 & n9272 ) | ( n9262 & n9272 ) ;
  assign n9746 = ( n9260 & ~n9273 ) | ( n9260 & n9745 ) | ( ~n9273 & n9745 ) ;
  assign n9747 = ( n9734 & n9744 ) | ( n9734 & n9746 ) | ( n9744 & n9746 ) ;
  assign n9748 = ( ~n9273 & n9275 ) | ( ~n9273 & n9285 ) | ( n9275 & n9285 ) ;
  assign n9749 = ( n9273 & ~n9286 ) | ( n9273 & n9748 ) | ( ~n9286 & n9748 ) ;
  assign n9750 = ~n2364 & n9593 ;
  assign n9751 = n41 & n2398 ;
  assign n9752 = n9750 | n9751 ;
  assign n9753 = ~x2 & n9752 ;
  assign n9754 = ~n2467 & n9600 ;
  assign n9755 = n9752 | n9754 ;
  assign n9756 = ( x2 & ~n5713 ) | ( x2 & n9590 ) | ( ~n5713 & n9590 ) ;
  assign n9757 = n5713 & n9591 ;
  assign n9758 = ( ~n9755 & n9756 ) | ( ~n9755 & n9757 ) | ( n9756 & n9757 ) ;
  assign n9759 = n9753 | n9758 ;
  assign n9760 = ( n9747 & n9749 ) | ( n9747 & n9759 ) | ( n9749 & n9759 ) ;
  assign n9761 = ( ~n9286 & n9288 ) | ( ~n9286 & n9298 ) | ( n9288 & n9298 ) ;
  assign n9762 = ( n9286 & ~n9299 ) | ( n9286 & n9761 ) | ( ~n9299 & n9761 ) ;
  assign n9763 = n41 & ~n2364 ;
  assign n9764 = x2 & n9763 ;
  assign n9765 = ~n2282 & n9593 ;
  assign n9766 = n2398 & n9600 ;
  assign n9767 = n9765 | n9766 ;
  assign n9768 = n9592 | n9767 ;
  assign n9769 = ( ~n5494 & n9767 ) | ( ~n5494 & n9768 ) | ( n9767 & n9768 ) ;
  assign n9770 = x2 & ~n9769 ;
  assign n9771 = ( ~x2 & n9763 ) | ( ~x2 & n9769 ) | ( n9763 & n9769 ) ;
  assign n9772 = ( ~n9764 & n9770 ) | ( ~n9764 & n9771 ) | ( n9770 & n9771 ) ;
  assign n9773 = ( n9760 & n9762 ) | ( n9760 & n9772 ) | ( n9762 & n9772 ) ;
  assign n9774 = ( ~n9299 & n9301 ) | ( ~n9299 & n9311 ) | ( n9301 & n9311 ) ;
  assign n9775 = ( n9299 & ~n9312 ) | ( n9299 & n9774 ) | ( ~n9312 & n9774 ) ;
  assign n9776 = n41 & ~n2282 ;
  assign n9777 = n2187 & n9593 ;
  assign n9778 = n9776 | n9777 ;
  assign n9779 = n9592 | n9778 ;
  assign n9780 = ( n5137 & n9778 ) | ( n5137 & n9779 ) | ( n9778 & n9779 ) ;
  assign n9781 = x2 & n9780 ;
  assign n9782 = ( x2 & n2364 ) | ( x2 & n9155 ) | ( n2364 & n9155 ) ;
  assign n9783 = n9780 | n9782 ;
  assign n9784 = ~n9781 & n9783 ;
  assign n9785 = ( n9773 & n9775 ) | ( n9773 & n9784 ) | ( n9775 & n9784 ) ;
  assign n9786 = n2102 & n9593 ;
  assign n9787 = n41 & n2187 ;
  assign n9788 = n9786 | n9787 ;
  assign n9789 = n9592 | n9788 ;
  assign n9790 = ( ~n5331 & n9788 ) | ( ~n5331 & n9789 ) | ( n9788 & n9789 ) ;
  assign n9791 = x2 & n9790 ;
  assign n9792 = ( x2 & n2282 ) | ( x2 & n9155 ) | ( n2282 & n9155 ) ;
  assign n9793 = n9790 | n9792 ;
  assign n9794 = ~n9791 & n9793 ;
  assign n9795 = ( ~n9312 & n9314 ) | ( ~n9312 & n9324 ) | ( n9314 & n9324 ) ;
  assign n9796 = ( n9312 & ~n9325 ) | ( n9312 & n9795 ) | ( ~n9325 & n9795 ) ;
  assign n9797 = ( n9785 & n9794 ) | ( n9785 & n9796 ) | ( n9794 & n9796 ) ;
  assign n9798 = ( ~n9325 & n9327 ) | ( ~n9325 & n9337 ) | ( n9327 & n9337 ) ;
  assign n9799 = ( n9325 & ~n9338 ) | ( n9325 & n9798 ) | ( ~n9338 & n9798 ) ;
  assign n9800 = ~n2041 & n9593 ;
  assign n9801 = n41 & n2102 ;
  assign n9802 = n9800 | n9801 ;
  assign n9803 = n2187 & n9600 ;
  assign n9804 = n9802 | n9803 ;
  assign n9805 = n9592 | n9804 ;
  assign n9806 = ( ~n4997 & n9804 ) | ( ~n4997 & n9805 ) | ( n9804 & n9805 ) ;
  assign n9807 = x2 & ~n9806 ;
  assign n9808 = ~x2 & n9806 ;
  assign n9809 = n9807 | n9808 ;
  assign n9810 = ( n9797 & n9799 ) | ( n9797 & n9809 ) | ( n9799 & n9809 ) ;
  assign n9811 = ( n9605 & n9615 ) | ( n9605 & n9810 ) | ( n9615 & n9810 ) ;
  assign n9812 = ( ~n9351 & n9353 ) | ( ~n9351 & n9363 ) | ( n9353 & n9363 ) ;
  assign n9813 = ( n9351 & ~n9364 ) | ( n9351 & n9812 ) | ( ~n9364 & n9812 ) ;
  assign n9814 = n41 & n1943 ;
  assign n9815 = ~n1841 & n9593 ;
  assign n9816 = n9814 | n9815 ;
  assign n9817 = n9592 | n9816 ;
  assign n9818 = ( ~n4753 & n9816 ) | ( ~n4753 & n9817 ) | ( n9816 & n9817 ) ;
  assign n9819 = x2 & n9818 ;
  assign n9820 = ( x2 & n2041 ) | ( x2 & n9155 ) | ( n2041 & n9155 ) ;
  assign n9821 = n9818 | n9820 ;
  assign n9822 = ~n9819 & n9821 ;
  assign n9823 = ( n9811 & n9813 ) | ( n9811 & n9822 ) | ( n9813 & n9822 ) ;
  assign n9824 = ( n9587 & n9603 ) | ( n9587 & n9823 ) | ( n9603 & n9823 ) ;
  assign n9825 = ( ~n9377 & n9379 ) | ( ~n9377 & n9389 ) | ( n9379 & n9389 ) ;
  assign n9826 = ( n9377 & ~n9390 ) | ( n9377 & n9825 ) | ( ~n9390 & n9825 ) ;
  assign n9827 = n1687 & n9593 ;
  assign n9828 = n9592 | n9827 ;
  assign n9829 = ( n4331 & n9827 ) | ( n4331 & n9828 ) | ( n9827 & n9828 ) ;
  assign n9830 = n41 & n1792 ;
  assign n9831 = ( x2 & ~n9829 ) | ( x2 & n9830 ) | ( ~n9829 & n9830 ) ;
  assign n9832 = ~x2 & n9829 ;
  assign n9833 = ~n1841 & n9600 ;
  assign n9834 = ( x2 & n9830 ) | ( x2 & n9833 ) | ( n9830 & n9833 ) ;
  assign n9835 = ( n9831 & n9832 ) | ( n9831 & ~n9834 ) | ( n9832 & ~n9834 ) ;
  assign n9836 = ( n9824 & n9826 ) | ( n9824 & n9835 ) | ( n9826 & n9835 ) ;
  assign n9837 = ( ~n9390 & n9392 ) | ( ~n9390 & n9402 ) | ( n9392 & n9402 ) ;
  assign n9838 = ( n9390 & ~n9403 ) | ( n9390 & n9837 ) | ( ~n9403 & n9837 ) ;
  assign n9839 = n41 & n1687 ;
  assign n9840 = n1600 & n9593 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = n9592 | n9841 ;
  assign n9843 = ( n4674 & n9841 ) | ( n4674 & n9842 ) | ( n9841 & n9842 ) ;
  assign n9844 = x2 & n9843 ;
  assign n9845 = ( x2 & ~n1792 ) | ( x2 & n9155 ) | ( ~n1792 & n9155 ) ;
  assign n9846 = n9843 | n9845 ;
  assign n9847 = ~n9844 & n9846 ;
  assign n9848 = ( n9836 & n9838 ) | ( n9836 & n9847 ) | ( n9838 & n9847 ) ;
  assign n9849 = ( ~n9403 & n9405 ) | ( ~n9403 & n9415 ) | ( n9405 & n9415 ) ;
  assign n9850 = ( n9403 & ~n9416 ) | ( n9403 & n9849 ) | ( ~n9416 & n9849 ) ;
  assign n9851 = ~n1529 & n9593 ;
  assign n9852 = n41 & n1600 ;
  assign n9853 = n9851 | n9852 ;
  assign n9854 = n9592 | n9853 ;
  assign n9855 = ( ~n4531 & n9853 ) | ( ~n4531 & n9854 ) | ( n9853 & n9854 ) ;
  assign n9856 = x2 & n9855 ;
  assign n9857 = ( x2 & ~n1687 ) | ( x2 & n9155 ) | ( ~n1687 & n9155 ) ;
  assign n9858 = n9855 | n9857 ;
  assign n9859 = ~n9856 & n9858 ;
  assign n9860 = ( n9848 & n9850 ) | ( n9848 & n9859 ) | ( n9850 & n9859 ) ;
  assign n9861 = n41 & ~n1529 ;
  assign n9862 = n1600 & n9600 ;
  assign n9863 = n1398 & n9593 ;
  assign n9864 = n9862 | n9863 ;
  assign n9865 = n9861 | n9864 ;
  assign n9866 = n9592 | n9865 ;
  assign n9867 = ( ~n4324 & n9865 ) | ( ~n4324 & n9866 ) | ( n9865 & n9866 ) ;
  assign n9868 = x2 & ~n9867 ;
  assign n9869 = ~x2 & n9867 ;
  assign n9870 = n9868 | n9869 ;
  assign n9871 = ( ~n9416 & n9418 ) | ( ~n9416 & n9428 ) | ( n9418 & n9428 ) ;
  assign n9872 = ( n9416 & ~n9429 ) | ( n9416 & n9871 ) | ( ~n9429 & n9871 ) ;
  assign n9873 = ( n9860 & n9870 ) | ( n9860 & n9872 ) | ( n9870 & n9872 ) ;
  assign n9874 = n1316 & n9593 ;
  assign n9875 = n9592 | n9874 ;
  assign n9876 = ( n4084 & n9874 ) | ( n4084 & n9875 ) | ( n9874 & n9875 ) ;
  assign n9877 = n41 & n1398 ;
  assign n9878 = ( x2 & ~n9876 ) | ( x2 & n9877 ) | ( ~n9876 & n9877 ) ;
  assign n9879 = ~x2 & n9876 ;
  assign n9880 = n1529 | n9154 ;
  assign n9881 = n9877 & n9880 ;
  assign n9882 = ( x2 & ~n9880 ) | ( x2 & n9881 ) | ( ~n9880 & n9881 ) ;
  assign n9883 = ( n9878 & n9879 ) | ( n9878 & ~n9882 ) | ( n9879 & ~n9882 ) ;
  assign n9884 = ( ~n9429 & n9431 ) | ( ~n9429 & n9441 ) | ( n9431 & n9441 ) ;
  assign n9885 = ( n9429 & ~n9442 ) | ( n9429 & n9884 ) | ( ~n9442 & n9884 ) ;
  assign n9886 = ( n9873 & n9883 ) | ( n9873 & n9885 ) | ( n9883 & n9885 ) ;
  assign n9887 = ( ~n9442 & n9452 ) | ( ~n9442 & n9454 ) | ( n9452 & n9454 ) ;
  assign n9888 = ( n9442 & ~n9455 ) | ( n9442 & n9887 ) | ( ~n9455 & n9887 ) ;
  assign n9889 = n41 & n1316 ;
  assign n9890 = x2 & n9889 ;
  assign n9891 = ~n1207 & n9593 ;
  assign n9892 = n1398 & n9600 ;
  assign n9893 = n9891 | n9892 ;
  assign n9894 = n9592 | n9893 ;
  assign n9895 = ( ~n4157 & n9893 ) | ( ~n4157 & n9894 ) | ( n9893 & n9894 ) ;
  assign n9896 = x2 & ~n9895 ;
  assign n9897 = ( ~x2 & n9889 ) | ( ~x2 & n9895 ) | ( n9889 & n9895 ) ;
  assign n9898 = ( ~n9890 & n9896 ) | ( ~n9890 & n9897 ) | ( n9896 & n9897 ) ;
  assign n9899 = ( n9886 & n9888 ) | ( n9886 & n9898 ) | ( n9888 & n9898 ) ;
  assign n9900 = ( ~n9455 & n9457 ) | ( ~n9455 & n9467 ) | ( n9457 & n9467 ) ;
  assign n9901 = ( n9455 & ~n9468 ) | ( n9455 & n9900 ) | ( ~n9468 & n9900 ) ;
  assign n9902 = ~n1118 & n9593 ;
  assign n9903 = n9592 | n9902 ;
  assign n9904 = ( n3841 & n9902 ) | ( n3841 & n9903 ) | ( n9902 & n9903 ) ;
  assign n9905 = n41 & ~n1207 ;
  assign n9906 = ( x2 & ~n9904 ) | ( x2 & n9905 ) | ( ~n9904 & n9905 ) ;
  assign n9907 = ~x2 & n9904 ;
  assign n9908 = n1316 & ~n9154 ;
  assign n9909 = n9905 & ~n9908 ;
  assign n9910 = ( x2 & n9908 ) | ( x2 & n9909 ) | ( n9908 & n9909 ) ;
  assign n9911 = ( n9906 & n9907 ) | ( n9906 & ~n9910 ) | ( n9907 & ~n9910 ) ;
  assign n9912 = ( n9899 & n9901 ) | ( n9899 & n9911 ) | ( n9901 & n9911 ) ;
  assign n9913 = ( ~n9468 & n9470 ) | ( ~n9468 & n9480 ) | ( n9470 & n9480 ) ;
  assign n9914 = ( n9468 & ~n9481 ) | ( n9468 & n9913 ) | ( ~n9481 & n9913 ) ;
  assign n9915 = n995 & n9593 ;
  assign n9916 = n41 & ~n1118 ;
  assign n9917 = n9915 | n9916 ;
  assign n9918 = n9592 | n9917 ;
  assign n9919 = ( n4173 & n9917 ) | ( n4173 & n9918 ) | ( n9917 & n9918 ) ;
  assign n9920 = x2 & n9919 ;
  assign n9921 = ( x2 & n1207 ) | ( x2 & n9155 ) | ( n1207 & n9155 ) ;
  assign n9922 = n9919 | n9921 ;
  assign n9923 = ~n9920 & n9922 ;
  assign n9924 = ( n9912 & n9914 ) | ( n9912 & n9923 ) | ( n9914 & n9923 ) ;
  assign n9925 = ( ~n9481 & n9483 ) | ( ~n9481 & n9493 ) | ( n9483 & n9493 ) ;
  assign n9926 = ( n9481 & ~n9494 ) | ( n9481 & n9925 ) | ( ~n9494 & n9925 ) ;
  assign n9927 = n859 & n9593 ;
  assign n9928 = n9592 | n9927 ;
  assign n9929 = ( ~n4034 & n9927 ) | ( ~n4034 & n9928 ) | ( n9927 & n9928 ) ;
  assign n9930 = n41 & n995 ;
  assign n9931 = ( x2 & ~n9929 ) | ( x2 & n9930 ) | ( ~n9929 & n9930 ) ;
  assign n9932 = ~x2 & n9929 ;
  assign n9933 = n1118 | n9154 ;
  assign n9934 = n9930 & n9933 ;
  assign n9935 = ( x2 & ~n9933 ) | ( x2 & n9934 ) | ( ~n9933 & n9934 ) ;
  assign n9936 = ( n9931 & n9932 ) | ( n9931 & ~n9935 ) | ( n9932 & ~n9935 ) ;
  assign n9937 = ( n9924 & n9926 ) | ( n9924 & n9936 ) | ( n9926 & n9936 ) ;
  assign n9938 = ~n3829 & n9591 ;
  assign n9939 = ( x2 & n3829 ) | ( x2 & n9590 ) | ( n3829 & n9590 ) ;
  assign n9940 = ~n721 & n9593 ;
  assign n9941 = n41 & n859 ;
  assign n9942 = n9940 | n9941 ;
  assign n9943 = n995 & n9600 ;
  assign n9944 = n9942 | n9943 ;
  assign n9945 = n9939 & n9944 ;
  assign n9946 = n9939 | n9942 ;
  assign n9947 = ( n9938 & ~n9945 ) | ( n9938 & n9946 ) | ( ~n9945 & n9946 ) ;
  assign n9948 = ( ~n9494 & n9496 ) | ( ~n9494 & n9506 ) | ( n9496 & n9506 ) ;
  assign n9949 = ( n9494 & ~n9507 ) | ( n9494 & n9948 ) | ( ~n9507 & n9948 ) ;
  assign n9950 = ( n9937 & n9947 ) | ( n9937 & n9949 ) | ( n9947 & n9949 ) ;
  assign n9951 = ( ~n9507 & n9509 ) | ( ~n9507 & n9519 ) | ( n9509 & n9519 ) ;
  assign n9952 = ( n9507 & ~n9520 ) | ( n9507 & n9951 ) | ( ~n9520 & n9951 ) ;
  assign n9953 = n859 & n9600 ;
  assign n9954 = n41 & ~n721 ;
  assign n9955 = n9953 | n9954 ;
  assign n9956 = n564 & n9593 ;
  assign n9957 = n9955 | n9956 ;
  assign n9958 = n9592 | n9957 ;
  assign n9959 = ( ~n3268 & n9957 ) | ( ~n3268 & n9958 ) | ( n9957 & n9958 ) ;
  assign n9960 = x2 & ~n9959 ;
  assign n9961 = ~x2 & n9959 ;
  assign n9962 = n9960 | n9961 ;
  assign n9963 = ( n9950 & n9952 ) | ( n9950 & n9962 ) | ( n9952 & n9962 ) ;
  assign n9964 = ~n3492 & n9592 ;
  assign n9965 = ~n3487 & n9593 ;
  assign n9966 = ~n721 & n9600 ;
  assign n9967 = n41 & n564 ;
  assign n9968 = n9966 | n9967 ;
  assign n9969 = n9965 | n9968 ;
  assign n9970 = ( x2 & ~n9964 ) | ( x2 & n9969 ) | ( ~n9964 & n9969 ) ;
  assign n9971 = ( x2 & n9964 ) | ( x2 & ~n9969 ) | ( n9964 & ~n9969 ) ;
  assign n9972 = ( ~x2 & n9970 ) | ( ~x2 & n9971 ) | ( n9970 & n9971 ) ;
  assign n9973 = ( n9520 & n9522 ) | ( n9520 & n9532 ) | ( n9522 & n9532 ) ;
  assign n9974 = ( n9522 & n9533 ) | ( n9522 & ~n9973 ) | ( n9533 & ~n9973 ) ;
  assign n9975 = ( n9963 & n9972 ) | ( n9963 & ~n9974 ) | ( n9972 & ~n9974 ) ;
  assign n9976 = ~n3601 & n9593 ;
  assign n9977 = n41 & ~n3487 ;
  assign n9978 = n9976 | n9977 ;
  assign n9979 = n9592 | n9978 ;
  assign n9980 = ( n3674 & n9978 ) | ( n3674 & n9979 ) | ( n9978 & n9979 ) ;
  assign n9981 = x2 & n9980 ;
  assign n9982 = ( x2 & ~n564 ) | ( x2 & n9155 ) | ( ~n564 & n9155 ) ;
  assign n9983 = n9980 | n9982 ;
  assign n9984 = ~n9981 & n9983 ;
  assign n9985 = ( n9533 & n9535 ) | ( n9533 & n9545 ) | ( n9535 & n9545 ) ;
  assign n9986 = ( n9535 & n9546 ) | ( n9535 & ~n9985 ) | ( n9546 & ~n9985 ) ;
  assign n9987 = ( n9975 & n9984 ) | ( n9975 & ~n9986 ) | ( n9984 & ~n9986 ) ;
  assign n9988 = ( ~n9546 & n9548 ) | ( ~n9546 & n9558 ) | ( n9548 & n9558 ) ;
  assign n9989 = ( n9546 & ~n9559 ) | ( n9546 & n9988 ) | ( ~n9559 & n9988 ) ;
  assign n9990 = n41 & ~n3601 ;
  assign n9991 = ~n3533 & n9593 ;
  assign n9992 = n9990 | n9991 ;
  assign n9993 = n9592 | n9992 ;
  assign n9994 = ( ~n4223 & n9992 ) | ( ~n4223 & n9993 ) | ( n9992 & n9993 ) ;
  assign n9995 = x2 & n9994 ;
  assign n9996 = ( x2 & n3487 ) | ( x2 & n9155 ) | ( n3487 & n9155 ) ;
  assign n9997 = n9994 | n9996 ;
  assign n9998 = ~n9995 & n9997 ;
  assign n9999 = ( n9987 & n9989 ) | ( n9987 & n9998 ) | ( n9989 & n9998 ) ;
  assign n10000 = ~n4058 & n9592 ;
  assign n10001 = ~n3601 & n9600 ;
  assign n10002 = n41 & ~n3533 ;
  assign n10003 = n10001 | n10002 ;
  assign n10004 = ~n3516 & n9593 ;
  assign n10005 = n10003 | n10004 ;
  assign n10006 = ( x2 & ~n10000 ) | ( x2 & n10005 ) | ( ~n10000 & n10005 ) ;
  assign n10007 = ( x2 & n10000 ) | ( x2 & ~n10005 ) | ( n10000 & ~n10005 ) ;
  assign n10008 = ( ~x2 & n10006 ) | ( ~x2 & n10007 ) | ( n10006 & n10007 ) ;
  assign n10009 = ( n9559 & n9561 ) | ( n9559 & ~n9571 ) | ( n9561 & ~n9571 ) ;
  assign n10010 = ( ~n9559 & n9572 ) | ( ~n9559 & n10009 ) | ( n9572 & n10009 ) ;
  assign n10011 = ( n9999 & n10008 ) | ( n9999 & ~n10010 ) | ( n10008 & ~n10010 ) ;
  assign n10012 = ( ~n9572 & n9582 ) | ( ~n9572 & n9584 ) | ( n9582 & n9584 ) ;
  assign n10013 = ( n9572 & ~n9585 ) | ( n9572 & n10012 ) | ( ~n9585 & n10012 ) ;
  assign n10014 = n41 & ~n3516 ;
  assign n10015 = n9592 | n10014 ;
  assign n10016 = ( n3609 & n10014 ) | ( n3609 & n10015 ) | ( n10014 & n10015 ) ;
  assign n10017 = ~n3533 & n9600 ;
  assign n10018 = ( x2 & n10016 ) | ( x2 & ~n10017 ) | ( n10016 & ~n10017 ) ;
  assign n10019 = ( x2 & n10016 ) | ( x2 & n10017 ) | ( n10016 & n10017 ) ;
  assign n10020 = n10018 & ~n10019 ;
  assign n10021 = ( n10011 & n10013 ) | ( n10011 & n10020 ) | ( n10013 & n10020 ) ;
  assign n10022 = ( ~n9143 & n9153 ) | ( ~n9143 & n9162 ) | ( n9153 & n9162 ) ;
  assign n10023 = ( n9143 & ~n9163 ) | ( n9143 & n10022 ) | ( ~n9163 & n10022 ) ;
  assign n10024 = ( n9585 & n10021 ) | ( n9585 & n10023 ) | ( n10021 & n10023 ) ;
  assign n10025 = ( ~n8732 & n8742 ) | ( ~n8732 & n9140 ) | ( n8742 & n9140 ) ;
  assign n10026 = ( n8732 & ~n9141 ) | ( n8732 & n10025 ) | ( ~n9141 & n10025 ) ;
  assign n10027 = ( n9163 & n10024 ) | ( n9163 & n10026 ) | ( n10024 & n10026 ) ;
  assign n10028 = ( ~n8718 & n8727 ) | ( ~n8718 & n8729 ) | ( n8727 & n8729 ) ;
  assign n10029 = ( n8718 & ~n8730 ) | ( n8718 & n10028 ) | ( ~n8730 & n10028 ) ;
  assign n10030 = ( n9141 & n10027 ) | ( n9141 & n10029 ) | ( n10027 & n10029 ) ;
  assign n10031 = ( n8335 & ~n8346 ) | ( n8335 & n8348 ) | ( ~n8346 & n8348 ) ;
  assign n10032 = ( ~n8335 & n8349 ) | ( ~n8335 & n10031 ) | ( n8349 & n10031 ) ;
  assign n10033 = ( n8730 & n10030 ) | ( n8730 & ~n10032 ) | ( n10030 & ~n10032 ) ;
  assign n10034 = ( ~n7978 & n7988 ) | ( ~n7978 & n7990 ) | ( n7988 & n7990 ) ;
  assign n10035 = ( n7978 & ~n7991 ) | ( n7978 & n10034 ) | ( ~n7991 & n10034 ) ;
  assign n10036 = ( n8349 & n10033 ) | ( n8349 & n10035 ) | ( n10033 & n10035 ) ;
  assign n10037 = ( ~n7642 & n7652 ) | ( ~n7642 & n7654 ) | ( n7652 & n7654 ) ;
  assign n10038 = ( ~n7652 & n7655 ) | ( ~n7652 & n10037 ) | ( n7655 & n10037 ) ;
  assign n10039 = ( n7991 & n10036 ) | ( n7991 & ~n10038 ) | ( n10036 & ~n10038 ) ;
  assign n10040 = ( ~n7332 & n7334 ) | ( ~n7332 & n7351 ) | ( n7334 & n7351 ) ;
  assign n10041 = ( n7332 & ~n7352 ) | ( n7332 & n10040 ) | ( ~n7352 & n10040 ) ;
  assign n10042 = ( n7655 & n10039 ) | ( n7655 & n10041 ) | ( n10039 & n10041 ) ;
  assign n10043 = ( ~n7050 & n7060 ) | ( ~n7050 & n7062 ) | ( n7060 & n7062 ) ;
  assign n10044 = ( n7050 & ~n7063 ) | ( n7050 & n10043 ) | ( ~n7063 & n10043 ) ;
  assign n10045 = ( n7352 & n10042 ) | ( n7352 & n10044 ) | ( n10042 & n10044 ) ;
  assign n10046 = ( ~n6794 & n6804 ) | ( ~n6794 & n6806 ) | ( n6804 & n6806 ) ;
  assign n10047 = ( n6794 & ~n6807 ) | ( n6794 & n10046 ) | ( ~n6807 & n10046 ) ;
  assign n10048 = ( n7063 & n10045 ) | ( n7063 & n10047 ) | ( n10045 & n10047 ) ;
  assign n10049 = ( ~n6560 & n6576 ) | ( ~n6560 & n6578 ) | ( n6576 & n6578 ) ;
  assign n10050 = ( n6560 & ~n6579 ) | ( n6560 & n10049 ) | ( ~n6579 & n10049 ) ;
  assign n10051 = ( n6807 & n10048 ) | ( n6807 & n10050 ) | ( n10048 & n10050 ) ;
  assign n10052 = ( ~n6442 & n6452 ) | ( ~n6442 & n6454 ) | ( n6452 & n6454 ) ;
  assign n10053 = ( n6442 & ~n6455 ) | ( n6442 & n10052 ) | ( ~n6455 & n10052 ) ;
  assign n10054 = ( n6579 & n10051 ) | ( n6579 & n10053 ) | ( n10051 & n10053 ) ;
  assign n10055 = ( ~n6328 & n6330 ) | ( ~n6328 & n6340 ) | ( n6330 & n6340 ) ;
  assign n10056 = ( n6328 & ~n6341 ) | ( n6328 & n10055 ) | ( ~n6341 & n10055 ) ;
  assign n10057 = ( n6455 & n10054 ) | ( n6455 & n10056 ) | ( n10054 & n10056 ) ;
  assign n10058 = ( ~n5902 & n5920 ) | ( ~n5902 & n5922 ) | ( n5920 & n5922 ) ;
  assign n10059 = ( n5902 & ~n5923 ) | ( n5902 & n10058 ) | ( ~n5923 & n10058 ) ;
  assign n10060 = ( n6341 & n10057 ) | ( n6341 & n10059 ) | ( n10057 & n10059 ) ;
  assign n10061 = ( n5801 & ~n5811 ) | ( n5801 & n5813 ) | ( ~n5811 & n5813 ) ;
  assign n10062 = ( ~n5801 & n5814 ) | ( ~n5801 & n10061 ) | ( n5814 & n10061 ) ;
  assign n10063 = ( n5923 & n10060 ) | ( n5923 & ~n10062 ) | ( n10060 & ~n10062 ) ;
  assign n10064 = ( ~n5582 & n5592 ) | ( ~n5582 & n5594 ) | ( n5592 & n5594 ) ;
  assign n10065 = ( n5582 & ~n5595 ) | ( n5582 & n10064 ) | ( ~n5595 & n10064 ) ;
  assign n10066 = ( n5814 & n10063 ) | ( n5814 & n10065 ) | ( n10063 & n10065 ) ;
  assign n10067 = ( n5406 & ~n5423 ) | ( n5406 & n5425 ) | ( ~n5423 & n5425 ) ;
  assign n10068 = ( ~n5406 & n5426 ) | ( ~n5406 & n10067 ) | ( n5426 & n10067 ) ;
  assign n10069 = ( n5595 & n10066 ) | ( n5595 & ~n10068 ) | ( n10066 & ~n10068 ) ;
  assign n10070 = ( ~n5245 & n5307 ) | ( ~n5245 & n5317 ) | ( n5307 & n5317 ) ;
  assign n10071 = ( n5245 & ~n5318 ) | ( n5245 & n10070 ) | ( ~n5318 & n10070 ) ;
  assign n10072 = ( n5426 & n10069 ) | ( n5426 & n10071 ) | ( n10069 & n10071 ) ;
  assign n10073 = ( ~n5230 & n5240 ) | ( ~n5230 & n5242 ) | ( n5240 & n5242 ) ;
  assign n10074 = ( n5230 & ~n5243 ) | ( n5230 & n10073 ) | ( ~n5243 & n10073 ) ;
  assign n10075 = ( n5318 & n10072 ) | ( n5318 & n10074 ) | ( n10072 & n10074 ) ;
  assign n10076 = ( n4867 & n4884 ) | ( n4867 & n4886 ) | ( n4884 & n4886 ) ;
  assign n10077 = ( n4886 & n4887 ) | ( n4886 & ~n10076 ) | ( n4887 & ~n10076 ) ;
  assign n10078 = ( n5243 & n10075 ) | ( n5243 & ~n10077 ) | ( n10075 & ~n10077 ) ;
  assign n10079 = ( ~n4711 & n4713 ) | ( ~n4711 & n4723 ) | ( n4713 & n4723 ) ;
  assign n10080 = ( n4711 & ~n4724 ) | ( n4711 & n10079 ) | ( ~n4724 & n10079 ) ;
  assign n10081 = ( n4887 & n10078 ) | ( n4887 & n10080 ) | ( n10078 & n10080 ) ;
  assign n10082 = ( ~n4635 & n4645 ) | ( ~n4635 & n4647 ) | ( n4645 & n4647 ) ;
  assign n10083 = ( ~n4645 & n4648 ) | ( ~n4645 & n10082 ) | ( n4648 & n10082 ) ;
  assign n10084 = ( n4724 & n10081 ) | ( n4724 & ~n10083 ) | ( n10081 & ~n10083 ) ;
  assign n10085 = ( ~n4577 & n4596 ) | ( ~n4577 & n4598 ) | ( n4596 & n4598 ) ;
  assign n10086 = ( n4577 & ~n4599 ) | ( n4577 & n10085 ) | ( ~n4599 & n10085 ) ;
  assign n10087 = ( n4648 & n10084 ) | ( n4648 & n10086 ) | ( n10084 & n10086 ) ;
  assign n10088 = ( ~n4238 & n4240 ) | ( ~n4238 & n4250 ) | ( n4240 & n4250 ) ;
  assign n10089 = ( n4238 & ~n4251 ) | ( n4238 & n10088 ) | ( ~n4251 & n10088 ) ;
  assign n10090 = ( n4599 & n10087 ) | ( n4599 & n10089 ) | ( n10087 & n10089 ) ;
  assign n10091 = ( ~n4196 & n4208 ) | ( ~n4196 & n4210 ) | ( n4208 & n4210 ) ;
  assign n10092 = ( n4196 & ~n4211 ) | ( n4196 & n10091 ) | ( ~n4211 & n10091 ) ;
  assign n10093 = ( n4251 & n10090 ) | ( n4251 & n10092 ) | ( n10090 & n10092 ) ;
  assign n10094 = ( n3837 & n4052 ) | ( n3837 & n4054 ) | ( n4052 & n4054 ) ;
  assign n10095 = ( n3837 & n4055 ) | ( n3837 & ~n10094 ) | ( n4055 & ~n10094 ) ;
  assign n10096 = n3501 & ~n3601 ;
  assign n10097 = ~n3533 & n4039 ;
  assign n10098 = n10096 | n10097 ;
  assign n10099 = n3541 | n10098 ;
  assign n10100 = ( ~n4223 & n10098 ) | ( ~n4223 & n10099 ) | ( n10098 & n10099 ) ;
  assign n10101 = ~n3487 & n3536 ;
  assign n10102 = n10100 | n10101 ;
  assign n10103 = ( ~n3516 & n3608 ) | ( ~n3516 & n4203 ) | ( n3608 & n4203 ) ;
  assign n10104 = ( n2083 & ~n3607 ) | ( n2083 & n10103 ) | ( ~n3607 & n10103 ) ;
  assign n10105 = ( n6269 & ~n10102 ) | ( n6269 & n10104 ) | ( ~n10102 & n10104 ) ;
  assign n10106 = ( n6269 & n10102 ) | ( n6269 & ~n10104 ) | ( n10102 & ~n10104 ) ;
  assign n10107 = ( ~n6269 & n10105 ) | ( ~n6269 & n10106 ) | ( n10105 & n10106 ) ;
  assign n10108 = n10095 | n10107 ;
  assign n10109 = n10095 & n10107 ;
  assign n10110 = n10108 & ~n10109 ;
  assign n10111 = ( n4211 & n10093 ) | ( n4211 & n10110 ) | ( n10093 & n10110 ) ;
  assign n10112 = x29 & n10102 ;
  assign n10113 = ~x26 & n10112 ;
  assign n10114 = ( ~n10095 & n10112 ) | ( ~n10095 & n10113 ) | ( n10112 & n10113 ) ;
  assign n10115 = ~x26 & n10104 ;
  assign n10116 = n3535 & ~n10104 ;
  assign n10117 = n10115 | n10116 ;
  assign n10118 = n6268 | n10095 ;
  assign n10119 = ( n10102 & n10117 ) | ( n10102 & n10118 ) | ( n10117 & n10118 ) ;
  assign n10120 = ~n10114 & n10119 ;
  assign n10121 = ( n4055 & n4067 ) | ( n4055 & ~n4069 ) | ( n4067 & ~n4069 ) ;
  assign n10122 = ( ~n4055 & n4070 ) | ( ~n4055 & n10121 ) | ( n4070 & n10121 ) ;
  assign n10123 = ( n10111 & n10120 ) | ( n10111 & n10122 ) | ( n10120 & n10122 ) ;
  assign n10124 = ( ~n3496 & n3613 ) | ( ~n3496 & n3684 ) | ( n3613 & n3684 ) ;
  assign n10125 = ( n3496 & ~n3685 ) | ( n3496 & n10124 ) | ( ~n3685 & n10124 ) ;
  assign n10126 = ( ~n4070 & n10123 ) | ( ~n4070 & n10125 ) | ( n10123 & n10125 ) ;
  assign n10127 = n1507 | n4953 ;
  assign n10128 = n964 | n1703 ;
  assign n10129 = n3623 | n3811 ;
  assign n10130 = n10128 | n10129 ;
  assign n10131 = n104 | n593 ;
  assign n10132 = n244 | n275 ;
  assign n10133 = n10131 | n10132 ;
  assign n10134 = n647 | n942 ;
  assign n10135 = n860 | n10134 ;
  assign n10136 = n10133 | n10135 ;
  assign n10137 = n10130 | n10136 ;
  assign n10138 = n10127 | n10137 ;
  assign n10139 = n440 | n661 ;
  assign n10140 = n711 | n10139 ;
  assign n10141 = n1722 | n10140 ;
  assign n10142 = n2257 | n10141 ;
  assign n10143 = n2434 | n2979 ;
  assign n10144 = n1106 | n10143 ;
  assign n10145 = n841 | n1843 ;
  assign n10146 = n789 | n10145 ;
  assign n10147 = n455 | n1044 ;
  assign n10148 = n494 | n10147 ;
  assign n10149 = n1998 | n10148 ;
  assign n10150 = n10146 | n10149 ;
  assign n10151 = n10144 | n10150 ;
  assign n10152 = n10142 | n10151 ;
  assign n10153 = n10138 | n10152 ;
  assign n10154 = n429 | n527 ;
  assign n10155 = n614 | n798 ;
  assign n10156 = n55 | n10155 ;
  assign n10157 = n10154 | n10156 ;
  assign n10158 = n417 | n10157 ;
  assign n10159 = n778 | n2092 ;
  assign n10160 = n2572 | n10159 ;
  assign n10161 = n10158 | n10160 ;
  assign n10162 = n153 | n176 ;
  assign n10163 = n318 | n10162 ;
  assign n10164 = n10161 | n10163 ;
  assign n10165 = n10153 | n10164 ;
  assign n10166 = n1812 & ~n10165 ;
  assign n10167 = ( n3402 & n3683 ) | ( n3402 & n10166 ) | ( n3683 & n10166 ) ;
  assign n10168 = ( ~n3402 & n3683 ) | ( ~n3402 & n10166 ) | ( n3683 & n10166 ) ;
  assign n10169 = ( n3402 & ~n10167 ) | ( n3402 & n10168 ) | ( ~n10167 & n10168 ) ;
  assign n10170 = n3273 & n3601 ;
  assign n10171 = n3270 & ~n3533 ;
  assign n10172 = n10170 | n10171 ;
  assign n10173 = n390 | n10172 ;
  assign n10174 = ( ~n4223 & n10172 ) | ( ~n4223 & n10173 ) | ( n10172 & n10173 ) ;
  assign n10175 = n3274 & ~n3601 ;
  assign n10176 = n10174 | n10175 ;
  assign n10177 = ( x29 & n65 ) | ( x29 & n3535 ) | ( n65 & n3535 ) ;
  assign n10178 = ( x29 & ~n3516 ) | ( x29 & n10177 ) | ( ~n3516 & n10177 ) ;
  assign n10179 = ( n10169 & n10176 ) | ( n10169 & n10178 ) | ( n10176 & n10178 ) ;
  assign n10180 = ( ~n10169 & n10176 ) | ( ~n10169 & n10178 ) | ( n10176 & n10178 ) ;
  assign n10181 = ( n10169 & ~n10179 ) | ( n10169 & n10180 ) | ( ~n10179 & n10180 ) ;
  assign n10182 = ( n3685 & n10126 ) | ( n3685 & ~n10181 ) | ( n10126 & ~n10181 ) ;
  assign n10183 = ( n3402 & ~n3683 ) | ( n3402 & n10166 ) | ( ~n3683 & n10166 ) ;
  assign n10184 = n3273 & ~n3601 ;
  assign n10185 = n390 | n10184 ;
  assign n10186 = ( ~n4058 & n10184 ) | ( ~n4058 & n10185 ) | ( n10184 & n10185 ) ;
  assign n10187 = n3274 & ~n3533 ;
  assign n10188 = n10186 | n10187 ;
  assign n10189 = n3480 | n3591 ;
  assign n10190 = n518 | n798 ;
  assign n10191 = n508 | n10190 ;
  assign n10192 = n1287 | n10191 ;
  assign n10193 = n3594 | n10192 ;
  assign n10194 = n2269 | n10193 ;
  assign n10195 = n252 | n419 ;
  assign n10196 = n517 | n10195 ;
  assign n10197 = n3384 | n10196 ;
  assign n10198 = n1967 | n10197 ;
  assign n10199 = n10194 | n10198 ;
  assign n10200 = n10189 | n10199 ;
  assign n10201 = n3419 | n3579 ;
  assign n10202 = n10200 | n10201 ;
  assign n10203 = n684 | n6013 ;
  assign n10204 = n3462 | n10203 ;
  assign n10205 = n10202 | n10204 ;
  assign n10206 = ( x29 & ~n10166 ) | ( x29 & n10205 ) | ( ~n10166 & n10205 ) ;
  assign n10207 = ( x29 & n10166 ) | ( x29 & ~n10205 ) | ( n10166 & ~n10205 ) ;
  assign n10208 = ( ~x29 & n10206 ) | ( ~x29 & n10207 ) | ( n10206 & n10207 ) ;
  assign n10209 = ( ~n10183 & n10188 ) | ( ~n10183 & n10208 ) | ( n10188 & n10208 ) ;
  assign n10210 = ( n10183 & n10188 ) | ( n10183 & n10208 ) | ( n10188 & n10208 ) ;
  assign n10211 = ( n10183 & n10209 ) | ( n10183 & ~n10210 ) | ( n10209 & ~n10210 ) ;
  assign n10212 = ( n10180 & n10182 ) | ( n10180 & n10211 ) | ( n10182 & n10211 ) ;
  assign n10213 = ( n10180 & ~n10182 ) | ( n10180 & n10211 ) | ( ~n10182 & n10211 ) ;
  assign n10214 = ( n10182 & ~n10212 ) | ( n10182 & n10213 ) | ( ~n10212 & n10213 ) ;
  assign n10215 = n41 & n10214 ;
  assign n10216 = x2 & n10215 ;
  assign n10217 = n3274 & ~n3516 ;
  assign n10218 = n390 | n10217 ;
  assign n10219 = ( n3609 & n10217 ) | ( n3609 & n10218 ) | ( n10217 & n10218 ) ;
  assign n10220 = n813 | n3525 ;
  assign n10221 = n1086 | n3463 ;
  assign n10222 = n3037 | n10221 ;
  assign n10223 = n3509 | n10222 ;
  assign n10224 = n2675 | n3424 ;
  assign n10225 = n10223 | n10224 ;
  assign n10226 = n5062 | n10225 ;
  assign n10227 = n10220 | n10226 ;
  assign n10228 = n3580 & ~n10189 ;
  assign n10229 = ~n10227 & n10228 ;
  assign n10230 = ( ~n10207 & n10219 ) | ( ~n10207 & n10229 ) | ( n10219 & n10229 ) ;
  assign n10231 = ( n10207 & n10219 ) | ( n10207 & ~n10229 ) | ( n10219 & ~n10229 ) ;
  assign n10232 = ( ~n10219 & n10230 ) | ( ~n10219 & n10231 ) | ( n10230 & n10231 ) ;
  assign n10233 = ( ~n10210 & n10212 ) | ( ~n10210 & n10232 ) | ( n10212 & n10232 ) ;
  assign n10234 = ( n10210 & n10212 ) | ( n10210 & ~n10232 ) | ( n10212 & ~n10232 ) ;
  assign n10235 = ( ~n10212 & n10233 ) | ( ~n10212 & n10234 ) | ( n10233 & n10234 ) ;
  assign n10236 = ( ~n3685 & n10126 ) | ( ~n3685 & n10181 ) | ( n10126 & n10181 ) ;
  assign n10237 = ( ~n10126 & n10182 ) | ( ~n10126 & n10236 ) | ( n10182 & n10236 ) ;
  assign n10238 = ( n4251 & ~n10090 ) | ( n4251 & n10092 ) | ( ~n10090 & n10092 ) ;
  assign n10239 = ( n10090 & ~n10093 ) | ( n10090 & n10238 ) | ( ~n10093 & n10238 ) ;
  assign n10240 = ( ~n4599 & n10087 ) | ( ~n4599 & n10089 ) | ( n10087 & n10089 ) ;
  assign n10241 = ( n4599 & ~n10090 ) | ( n4599 & n10240 ) | ( ~n10090 & n10240 ) ;
  assign n10242 = ( n4648 & ~n10084 ) | ( n4648 & n10086 ) | ( ~n10084 & n10086 ) ;
  assign n10243 = ( n10084 & ~n10087 ) | ( n10084 & n10242 ) | ( ~n10087 & n10242 ) ;
  assign n10244 = ( ~n4887 & n10078 ) | ( ~n4887 & n10080 ) | ( n10078 & n10080 ) ;
  assign n10245 = ( n4887 & ~n10081 ) | ( n4887 & n10244 ) | ( ~n10081 & n10244 ) ;
  assign n10246 = ( n5318 & ~n10072 ) | ( n5318 & n10074 ) | ( ~n10072 & n10074 ) ;
  assign n10247 = ( n10072 & ~n10075 ) | ( n10072 & n10246 ) | ( ~n10075 & n10246 ) ;
  assign n10248 = ( ~n5595 & n10066 ) | ( ~n5595 & n10068 ) | ( n10066 & n10068 ) ;
  assign n10249 = ( ~n10066 & n10069 ) | ( ~n10066 & n10248 ) | ( n10069 & n10248 ) ;
  assign n10250 = ( n5814 & ~n10063 ) | ( n5814 & n10065 ) | ( ~n10063 & n10065 ) ;
  assign n10251 = ( n10063 & ~n10066 ) | ( n10063 & n10250 ) | ( ~n10066 & n10250 ) ;
  assign n10252 = ( ~n5923 & n10060 ) | ( ~n5923 & n10062 ) | ( n10060 & n10062 ) ;
  assign n10253 = ( ~n10060 & n10063 ) | ( ~n10060 & n10252 ) | ( n10063 & n10252 ) ;
  assign n10254 = ( ~n6341 & n10057 ) | ( ~n6341 & n10059 ) | ( n10057 & n10059 ) ;
  assign n10255 = ( n6341 & ~n10060 ) | ( n6341 & n10254 ) | ( ~n10060 & n10254 ) ;
  assign n10256 = ( n6455 & ~n10054 ) | ( n6455 & n10056 ) | ( ~n10054 & n10056 ) ;
  assign n10257 = ( n10054 & ~n10057 ) | ( n10054 & n10256 ) | ( ~n10057 & n10256 ) ;
  assign n10258 = ( n6579 & ~n10051 ) | ( n6579 & n10053 ) | ( ~n10051 & n10053 ) ;
  assign n10259 = ( n10051 & ~n10054 ) | ( n10051 & n10258 ) | ( ~n10054 & n10258 ) ;
  assign n10260 = ( n6807 & ~n10048 ) | ( n6807 & n10050 ) | ( ~n10048 & n10050 ) ;
  assign n10261 = ( n10048 & ~n10051 ) | ( n10048 & n10260 ) | ( ~n10051 & n10260 ) ;
  assign n10262 = ( ~n7063 & n10045 ) | ( ~n7063 & n10047 ) | ( n10045 & n10047 ) ;
  assign n10263 = ( n7063 & ~n10048 ) | ( n7063 & n10262 ) | ( ~n10048 & n10262 ) ;
  assign n10264 = ( ~n7352 & n10042 ) | ( ~n7352 & n10044 ) | ( n10042 & n10044 ) ;
  assign n10265 = ( n7352 & ~n10045 ) | ( n7352 & n10264 ) | ( ~n10045 & n10264 ) ;
  assign n10266 = ( n7655 & ~n10039 ) | ( n7655 & n10041 ) | ( ~n10039 & n10041 ) ;
  assign n10267 = ( n10039 & ~n10042 ) | ( n10039 & n10266 ) | ( ~n10042 & n10266 ) ;
  assign n10268 = ( ~n7991 & n10036 ) | ( ~n7991 & n10038 ) | ( n10036 & n10038 ) ;
  assign n10269 = ( ~n10036 & n10039 ) | ( ~n10036 & n10268 ) | ( n10039 & n10268 ) ;
  assign n10270 = ( n8349 & ~n10033 ) | ( n8349 & n10035 ) | ( ~n10033 & n10035 ) ;
  assign n10271 = ( n10033 & ~n10036 ) | ( n10033 & n10270 ) | ( ~n10036 & n10270 ) ;
  assign n10272 = ( ~n9141 & n10027 ) | ( ~n9141 & n10029 ) | ( n10027 & n10029 ) ;
  assign n10273 = ( n9141 & ~n10030 ) | ( n9141 & n10272 ) | ( ~n10030 & n10272 ) ;
  assign n10274 = ( n9163 & ~n10024 ) | ( n9163 & n10026 ) | ( ~n10024 & n10026 ) ;
  assign n10275 = ( n10024 & ~n10027 ) | ( n10024 & n10274 ) | ( ~n10027 & n10274 ) ;
  assign n10276 = ( n9585 & ~n10021 ) | ( n9585 & n10023 ) | ( ~n10021 & n10023 ) ;
  assign n10277 = ( n10021 & ~n10024 ) | ( n10021 & n10276 ) | ( ~n10024 & n10276 ) ;
  assign n10278 = ( n9999 & ~n10008 ) | ( n9999 & n10010 ) | ( ~n10008 & n10010 ) ;
  assign n10279 = ( ~n9999 & n10011 ) | ( ~n9999 & n10278 ) | ( n10011 & n10278 ) ;
  assign n10280 = ( ~n9987 & n9989 ) | ( ~n9987 & n9998 ) | ( n9989 & n9998 ) ;
  assign n10281 = ( n9987 & ~n9999 ) | ( n9987 & n10280 ) | ( ~n9999 & n10280 ) ;
  assign n10282 = ( n9975 & ~n9984 ) | ( n9975 & n9986 ) | ( ~n9984 & n9986 ) ;
  assign n10283 = ( ~n9975 & n9987 ) | ( ~n9975 & n10282 ) | ( n9987 & n10282 ) ;
  assign n10284 = ( n9963 & ~n9972 ) | ( n9963 & n9974 ) | ( ~n9972 & n9974 ) ;
  assign n10285 = ( ~n9963 & n9975 ) | ( ~n9963 & n10284 ) | ( n9975 & n10284 ) ;
  assign n10286 = ~n10283 & n10285 ;
  assign n10287 = ~n10281 & n10286 ;
  assign n10288 = ( ~n10281 & n10283 ) | ( ~n10281 & n10287 ) | ( n10283 & n10287 ) ;
  assign n10289 = n10279 | n10288 ;
  assign n10290 = ( n10011 & ~n10013 ) | ( n10011 & n10020 ) | ( ~n10013 & n10020 ) ;
  assign n10291 = ( n10013 & ~n10021 ) | ( n10013 & n10290 ) | ( ~n10021 & n10290 ) ;
  assign n10292 = n10289 & ~n10291 ;
  assign n10293 = n10277 & ~n10292 ;
  assign n10294 = n10275 | n10293 ;
  assign n10295 = n10273 & n10294 ;
  assign n10296 = ( ~n8730 & n10030 ) | ( ~n8730 & n10032 ) | ( n10030 & n10032 ) ;
  assign n10297 = ( ~n10030 & n10033 ) | ( ~n10030 & n10296 ) | ( n10033 & n10296 ) ;
  assign n10298 = ~n10295 & n10297 ;
  assign n10299 = n10271 & ~n10298 ;
  assign n10300 = n10269 & ~n10299 ;
  assign n10301 = n10267 & ~n10300 ;
  assign n10302 = n10265 | n10301 ;
  assign n10303 = n10263 & n10302 ;
  assign n10304 = n10261 | n10303 ;
  assign n10305 = n10259 & n10304 ;
  assign n10306 = n10257 | n10305 ;
  assign n10307 = n10255 & n10306 ;
  assign n10308 = n10253 & ~n10307 ;
  assign n10309 = n10251 & ~n10308 ;
  assign n10310 = n10249 & ~n10309 ;
  assign n10311 = ( n5426 & ~n10069 ) | ( n5426 & n10071 ) | ( ~n10069 & n10071 ) ;
  assign n10312 = ( n10069 & ~n10072 ) | ( n10069 & n10311 ) | ( ~n10072 & n10311 ) ;
  assign n10313 = ~n10310 & n10312 ;
  assign n10314 = n10247 | n10313 ;
  assign n10315 = ( ~n5243 & n10075 ) | ( ~n5243 & n10077 ) | ( n10075 & n10077 ) ;
  assign n10316 = ( ~n10075 & n10078 ) | ( ~n10075 & n10315 ) | ( n10078 & n10315 ) ;
  assign n10317 = n10314 & ~n10316 ;
  assign n10318 = n10245 | n10317 ;
  assign n10319 = ( ~n4724 & n10081 ) | ( ~n4724 & n10083 ) | ( n10081 & n10083 ) ;
  assign n10320 = ( ~n10081 & n10084 ) | ( ~n10081 & n10319 ) | ( n10084 & n10319 ) ;
  assign n10321 = n10318 & ~n10320 ;
  assign n10322 = n10243 | n10321 ;
  assign n10323 = n10241 & n10322 ;
  assign n10324 = n10239 | n10323 ;
  assign n10325 = ( n4211 & ~n10093 ) | ( n4211 & n10110 ) | ( ~n10093 & n10110 ) ;
  assign n10326 = ( n10093 & ~n10111 ) | ( n10093 & n10325 ) | ( ~n10111 & n10325 ) ;
  assign n10327 = n10324 & n10326 ;
  assign n10328 = ( n10111 & n10120 ) | ( n10111 & ~n10122 ) | ( n10120 & ~n10122 ) ;
  assign n10329 = ( n10122 & ~n10123 ) | ( n10122 & n10328 ) | ( ~n10123 & n10328 ) ;
  assign n10330 = n10327 | n10329 ;
  assign n10331 = ( n4070 & n10123 ) | ( n4070 & ~n10125 ) | ( n10123 & ~n10125 ) ;
  assign n10332 = ( ~n10123 & n10126 ) | ( ~n10123 & n10331 ) | ( n10126 & n10331 ) ;
  assign n10333 = n10330 & ~n10332 ;
  assign n10334 = n10237 & ~n10333 ;
  assign n10335 = n10214 & ~n10334 ;
  assign n10336 = n10281 & ~n10283 ;
  assign n10337 = n10279 & ~n10336 ;
  assign n10338 = n10291 & ~n10337 ;
  assign n10339 = n10277 | n10338 ;
  assign n10340 = n10275 & n10339 ;
  assign n10341 = n10273 | n10340 ;
  assign n10342 = ~n10297 & n10341 ;
  assign n10343 = n10271 | n10342 ;
  assign n10344 = ~n10269 & n10343 ;
  assign n10345 = n10267 | n10344 ;
  assign n10346 = n10265 & n10345 ;
  assign n10347 = n10263 | n10346 ;
  assign n10348 = n10261 & n10347 ;
  assign n10349 = n10259 | n10348 ;
  assign n10350 = n10257 & n10349 ;
  assign n10351 = n10255 | n10350 ;
  assign n10352 = ~n10253 & n10351 ;
  assign n10353 = n10251 | n10352 ;
  assign n10354 = ~n10249 & n10353 ;
  assign n10355 = n10312 | n10354 ;
  assign n10356 = n10247 & n10355 ;
  assign n10357 = n10316 & ~n10356 ;
  assign n10358 = n10245 & ~n10357 ;
  assign n10359 = n10320 & ~n10358 ;
  assign n10360 = n10243 & ~n10359 ;
  assign n10361 = n10241 | n10360 ;
  assign n10362 = n10239 & n10361 ;
  assign n10363 = n10326 | n10362 ;
  assign n10364 = n10329 & n10363 ;
  assign n10365 = n10332 & ~n10364 ;
  assign n10366 = n10237 | n10365 ;
  assign n10367 = ~n10214 & n10366 ;
  assign n10368 = ( n10235 & n10335 ) | ( n10235 & n10367 ) | ( n10335 & n10367 ) ;
  assign n10369 = n10235 | n10335 ;
  assign n10370 = ( ~n10235 & n10335 ) | ( ~n10235 & n10367 ) | ( n10335 & n10367 ) ;
  assign n10371 = ( ~n10368 & n10369 ) | ( ~n10368 & n10370 ) | ( n10369 & n10370 ) ;
  assign n10372 = n9600 & ~n10237 ;
  assign n10373 = n9593 | n10372 ;
  assign n10374 = ( ~n10235 & n10372 ) | ( ~n10235 & n10373 ) | ( n10372 & n10373 ) ;
  assign n10375 = n9592 | n10374 ;
  assign n10376 = ( n10371 & n10374 ) | ( n10371 & n10375 ) | ( n10374 & n10375 ) ;
  assign n10377 = x2 & ~n10376 ;
  assign n10378 = ( ~x2 & n10215 ) | ( ~x2 & n10376 ) | ( n10215 & n10376 ) ;
  assign n10379 = ( ~n10216 & n10377 ) | ( ~n10216 & n10378 ) | ( n10377 & n10378 ) ;
  assign n10380 = n10330 & n10365 ;
  assign n10381 = n10329 & ~n10363 ;
  assign n10382 = ( ~n10329 & n10333 ) | ( ~n10329 & n10381 ) | ( n10333 & n10381 ) ;
  assign n10383 = ( n10332 & ~n10380 ) | ( n10332 & n10382 ) | ( ~n10380 & n10382 ) ;
  assign n10384 = n9592 & ~n10383 ;
  assign n10385 = n9593 & ~n10332 ;
  assign n10386 = n41 & n10329 ;
  assign n10387 = n10385 | n10386 ;
  assign n10388 = x2 | n10387 ;
  assign n10389 = ( ~n10384 & n10387 ) | ( ~n10384 & n10388 ) | ( n10387 & n10388 ) ;
  assign n10390 = n9591 & ~n10383 ;
  assign n10391 = n10389 | n10390 ;
  assign n10392 = n9600 & n10326 ;
  assign n10393 = ( x2 & n10387 ) | ( x2 & n10392 ) | ( n10387 & n10392 ) ;
  assign n10394 = n10391 & ~n10393 ;
  assign n10395 = ( ~n10327 & n10329 ) | ( ~n10327 & n10363 ) | ( n10329 & n10363 ) ;
  assign n10396 = ~n10327 & n10329 ;
  assign n10397 = ( n10381 & n10395 ) | ( n10381 & ~n10396 ) | ( n10395 & ~n10396 ) ;
  assign n10398 = n9592 & n10397 ;
  assign n10399 = n9593 & n10329 ;
  assign n10400 = n41 & n10326 ;
  assign n10401 = n10399 | n10400 ;
  assign n10402 = x2 | n10401 ;
  assign n10403 = ( ~n10398 & n10401 ) | ( ~n10398 & n10402 ) | ( n10401 & n10402 ) ;
  assign n10404 = n9591 & n10397 ;
  assign n10405 = n10403 | n10404 ;
  assign n10406 = n9600 & n10239 ;
  assign n10407 = ( x2 & n10401 ) | ( x2 & n10406 ) | ( n10401 & n10406 ) ;
  assign n10408 = n10405 & ~n10407 ;
  assign n10409 = n40 & ~n10320 ;
  assign n10410 = x5 & n10409 ;
  assign n10411 = ( n10318 & ~n10320 ) | ( n10318 & n10358 ) | ( ~n10320 & n10358 ) ;
  assign n10412 = ~n10318 & n10320 ;
  assign n10413 = ( n10318 & n10320 ) | ( n10318 & ~n10358 ) | ( n10320 & ~n10358 ) ;
  assign n10414 = ( n10411 & n10412 ) | ( n10411 & n10413 ) | ( n10412 & n10413 ) ;
  assign n10415 = n8721 & n10245 ;
  assign n10416 = n8340 & ~n10316 ;
  assign n10417 = n10415 | n10416 ;
  assign n10418 = n8341 | n10417 ;
  assign n10419 = ( ~n10414 & n10417 ) | ( ~n10414 & n10418 ) | ( n10417 & n10418 ) ;
  assign n10420 = x5 & ~n10419 ;
  assign n10421 = ( ~x5 & n10409 ) | ( ~x5 & n10419 ) | ( n10409 & n10419 ) ;
  assign n10422 = ( ~n10410 & n10420 ) | ( ~n10410 & n10421 ) | ( n10420 & n10421 ) ;
  assign n10423 = n7644 & n10312 ;
  assign n10424 = x8 & n10423 ;
  assign n10425 = n10247 & ~n10355 ;
  assign n10426 = ( n10247 & ~n10313 ) | ( n10247 & n10355 ) | ( ~n10313 & n10355 ) ;
  assign n10427 = n10247 & ~n10313 ;
  assign n10428 = ( n10425 & n10426 ) | ( n10425 & ~n10427 ) | ( n10426 & ~n10427 ) ;
  assign n10429 = n7341 & ~n10249 ;
  assign n10430 = n7345 | n10429 ;
  assign n10431 = ( n10247 & n10429 ) | ( n10247 & n10430 ) | ( n10429 & n10430 ) ;
  assign n10432 = n7346 | n10431 ;
  assign n10433 = ( n10428 & n10431 ) | ( n10428 & n10432 ) | ( n10431 & n10432 ) ;
  assign n10434 = x8 & ~n10433 ;
  assign n10435 = ( ~x8 & n10423 ) | ( ~x8 & n10433 ) | ( n10423 & n10433 ) ;
  assign n10436 = ( ~n10424 & n10434 ) | ( ~n10424 & n10435 ) | ( n10434 & n10435 ) ;
  assign n10437 = n7644 & n10251 ;
  assign n10438 = x8 & n10437 ;
  assign n10439 = n10249 & ~n10353 ;
  assign n10440 = ( n10249 & ~n10309 ) | ( n10249 & n10353 ) | ( ~n10309 & n10353 ) ;
  assign n10441 = ( ~n10310 & n10439 ) | ( ~n10310 & n10440 ) | ( n10439 & n10440 ) ;
  assign n10442 = n7341 & ~n10253 ;
  assign n10443 = n7345 | n10442 ;
  assign n10444 = ( ~n10249 & n10442 ) | ( ~n10249 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10445 = n7346 | n10444 ;
  assign n10446 = ( ~n10441 & n10444 ) | ( ~n10441 & n10445 ) | ( n10444 & n10445 ) ;
  assign n10447 = x8 & ~n10446 ;
  assign n10448 = ( ~x8 & n10437 ) | ( ~x8 & n10446 ) | ( n10437 & n10446 ) ;
  assign n10449 = ( ~n10438 & n10447 ) | ( ~n10438 & n10448 ) | ( n10447 & n10448 ) ;
  assign n10450 = n6570 & n10291 ;
  assign n10451 = x11 & n10450 ;
  assign n10452 = ~n10289 & n10291 ;
  assign n10453 = ( n10289 & n10291 ) | ( n10289 & ~n10337 ) | ( n10291 & ~n10337 ) ;
  assign n10454 = ( ~n10338 & n10452 ) | ( ~n10338 & n10453 ) | ( n10452 & n10453 ) ;
  assign n10455 = n6796 & ~n10279 ;
  assign n10456 = n6567 & n10281 ;
  assign n10457 = n10455 | n10456 ;
  assign n10458 = n6571 | n10457 ;
  assign n10459 = ( n10454 & n10457 ) | ( n10454 & n10458 ) | ( n10457 & n10458 ) ;
  assign n10460 = x11 & ~n10459 ;
  assign n10461 = ( ~x11 & n10450 ) | ( ~x11 & n10459 ) | ( n10450 & n10459 ) ;
  assign n10462 = ( ~n10451 & n10460 ) | ( ~n10451 & n10461 ) | ( n10460 & n10461 ) ;
  assign n10463 = n10281 & ~n10286 ;
  assign n10464 = n10287 | n10463 ;
  assign n10465 = n6571 & n10464 ;
  assign n10466 = n6570 & n10281 ;
  assign n10467 = n6796 & ~n10283 ;
  assign n10468 = n6567 & ~n10285 ;
  assign n10469 = n10467 | n10468 ;
  assign n10470 = n10466 | n10469 ;
  assign n10471 = n10465 | n10470 ;
  assign n10472 = n6571 & n10283 ;
  assign n10473 = n6796 & ~n10285 ;
  assign n10474 = ( ~n10285 & n10472 ) | ( ~n10285 & n10473 ) | ( n10472 & n10473 ) ;
  assign n10475 = ( n6568 & n6570 ) | ( n6568 & n10285 ) | ( n6570 & n10285 ) ;
  assign n10476 = ~n10283 & n10475 ;
  assign n10477 = n10474 | n10476 ;
  assign n10478 = n6568 & ~n10285 ;
  assign n10479 = x11 & ~n10478 ;
  assign n10480 = ~n10477 & n10479 ;
  assign n10481 = ~n10471 & n10480 ;
  assign n10482 = n5910 & ~n10285 ;
  assign n10483 = n10481 | n10482 ;
  assign n10484 = ( ~n10279 & n10288 ) | ( ~n10279 & n10336 ) | ( n10288 & n10336 ) ;
  assign n10485 = n10279 & ~n10288 ;
  assign n10486 = ( n10279 & n10288 ) | ( n10279 & n10336 ) | ( n10288 & n10336 ) ;
  assign n10487 = ( n10484 & n10485 ) | ( n10484 & ~n10486 ) | ( n10485 & ~n10486 ) ;
  assign n10488 = n6571 & n10487 ;
  assign n10489 = n6570 & ~n10279 ;
  assign n10490 = n6796 & n10281 ;
  assign n10491 = n6567 & ~n10283 ;
  assign n10492 = n10490 | n10491 ;
  assign n10493 = n10489 | n10492 ;
  assign n10494 = n10488 | n10493 ;
  assign n10495 = ~x11 & x12 ;
  assign n10496 = ~n10285 & n10495 ;
  assign n10497 = n10494 & n10496 ;
  assign n10498 = n10494 & ~n10496 ;
  assign n10499 = ( n10483 & n10497 ) | ( n10483 & ~n10498 ) | ( n10497 & ~n10498 ) ;
  assign n10500 = n5915 & n10283 ;
  assign n10501 = n6332 & ~n10285 ;
  assign n10502 = ( ~n10285 & n10500 ) | ( ~n10285 & n10501 ) | ( n10500 & n10501 ) ;
  assign n10503 = n5911 & n10286 ;
  assign n10504 = ( n5914 & ~n10283 ) | ( n5914 & n10503 ) | ( ~n10283 & n10503 ) ;
  assign n10505 = n10502 | n10504 ;
  assign n10506 = n5911 & ~n10285 ;
  assign n10507 = n10505 | n10506 ;
  assign n10508 = ( x14 & ~n10505 ) | ( x14 & n10506 ) | ( ~n10505 & n10506 ) ;
  assign n10509 = x14 & ~n10505 ;
  assign n10510 = ( n10507 & ~n10508 ) | ( n10507 & n10509 ) | ( ~n10508 & n10509 ) ;
  assign n10511 = ( n10462 & n10499 ) | ( n10462 & n10510 ) | ( n10499 & n10510 ) ;
  assign n10512 = n6796 & n10291 ;
  assign n10513 = x11 & n10512 ;
  assign n10514 = n10277 & n10338 ;
  assign n10515 = ( ~n10277 & n10292 ) | ( ~n10277 & n10338 ) | ( n10292 & n10338 ) ;
  assign n10516 = ( n10293 & ~n10514 ) | ( n10293 & n10515 ) | ( ~n10514 & n10515 ) ;
  assign n10517 = n6567 & ~n10279 ;
  assign n10518 = n6570 | n10517 ;
  assign n10519 = ( n10277 & n10517 ) | ( n10277 & n10518 ) | ( n10517 & n10518 ) ;
  assign n10520 = n6571 | n10519 ;
  assign n10521 = ( ~n10516 & n10519 ) | ( ~n10516 & n10520 ) | ( n10519 & n10520 ) ;
  assign n10522 = x11 & ~n10521 ;
  assign n10523 = ( ~x11 & n10512 ) | ( ~x11 & n10521 ) | ( n10512 & n10521 ) ;
  assign n10524 = ( ~n10513 & n10522 ) | ( ~n10513 & n10523 ) | ( n10522 & n10523 ) ;
  assign n10525 = x14 & n10507 ;
  assign n10526 = n5915 & n10464 ;
  assign n10527 = n5914 & n10281 ;
  assign n10528 = n6332 & ~n10283 ;
  assign n10529 = n5909 & ~n10285 ;
  assign n10530 = n10528 | n10529 ;
  assign n10531 = n10527 | n10530 ;
  assign n10532 = n10526 | n10531 ;
  assign n10533 = n10525 & ~n10532 ;
  assign n10534 = ~n10525 & n10532 ;
  assign n10535 = n10533 | n10534 ;
  assign n10536 = ( n10511 & n10524 ) | ( n10511 & n10535 ) | ( n10524 & n10535 ) ;
  assign n10537 = n5915 & n10487 ;
  assign n10538 = n5914 & ~n10279 ;
  assign n10539 = n6332 & n10281 ;
  assign n10540 = n5909 & ~n10283 ;
  assign n10541 = n10539 | n10540 ;
  assign n10542 = n10538 | n10541 ;
  assign n10543 = n10537 | n10542 ;
  assign n10544 = x14 & ~n10507 ;
  assign n10545 = ~n10532 & n10544 ;
  assign n10546 = n10285 | n10545 ;
  assign n10547 = n10543 & ~n10546 ;
  assign n10548 = ~n10543 & n10545 ;
  assign n10549 = ( x15 & n10547 ) | ( x15 & n10548 ) | ( n10547 & n10548 ) ;
  assign n10550 = x15 | n10285 ;
  assign n10551 = ~x14 & n10550 ;
  assign n10552 = ( n10545 & n10550 ) | ( n10545 & n10551 ) | ( n10550 & n10551 ) ;
  assign n10553 = n10546 & ~n10552 ;
  assign n10554 = ~n10543 & n10553 ;
  assign n10555 = ( ~n10285 & n10543 ) | ( ~n10285 & n10550 ) | ( n10543 & n10550 ) ;
  assign n10556 = ( n10547 & ~n10553 ) | ( n10547 & n10555 ) | ( ~n10553 & n10555 ) ;
  assign n10557 = ( ~n10549 & n10554 ) | ( ~n10549 & n10556 ) | ( n10554 & n10556 ) ;
  assign n10558 = n6796 & n10277 ;
  assign n10559 = x11 & n10558 ;
  assign n10560 = ( n10275 & ~n10293 ) | ( n10275 & n10339 ) | ( ~n10293 & n10339 ) ;
  assign n10561 = n10275 & ~n10293 ;
  assign n10562 = ( n10275 & n10293 ) | ( n10275 & ~n10339 ) | ( n10293 & ~n10339 ) ;
  assign n10563 = ( n10560 & ~n10561 ) | ( n10560 & n10562 ) | ( ~n10561 & n10562 ) ;
  assign n10564 = n6567 & n10291 ;
  assign n10565 = n6570 | n10564 ;
  assign n10566 = ( n10275 & n10564 ) | ( n10275 & n10565 ) | ( n10564 & n10565 ) ;
  assign n10567 = n6571 | n10566 ;
  assign n10568 = ( n10563 & n10566 ) | ( n10563 & n10567 ) | ( n10566 & n10567 ) ;
  assign n10569 = x11 & ~n10568 ;
  assign n10570 = ( ~x11 & n10558 ) | ( ~x11 & n10568 ) | ( n10558 & n10568 ) ;
  assign n10571 = ( ~n10559 & n10569 ) | ( ~n10559 & n10570 ) | ( n10569 & n10570 ) ;
  assign n10572 = ( n10536 & n10557 ) | ( n10536 & n10571 ) | ( n10557 & n10571 ) ;
  assign n10573 = n6796 & n10275 ;
  assign n10574 = x11 & n10573 ;
  assign n10575 = n10273 & n10340 ;
  assign n10576 = ( n10273 & n10294 ) | ( n10273 & ~n10340 ) | ( n10294 & ~n10340 ) ;
  assign n10577 = ( ~n10295 & n10575 ) | ( ~n10295 & n10576 ) | ( n10575 & n10576 ) ;
  assign n10578 = n6567 & n10277 ;
  assign n10579 = n6570 | n10578 ;
  assign n10580 = ( n10273 & n10578 ) | ( n10273 & n10579 ) | ( n10578 & n10579 ) ;
  assign n10581 = n6571 | n10580 ;
  assign n10582 = ( n10577 & n10580 ) | ( n10577 & n10581 ) | ( n10580 & n10581 ) ;
  assign n10583 = x11 & ~n10582 ;
  assign n10584 = ( ~x11 & n10573 ) | ( ~x11 & n10582 ) | ( n10573 & n10582 ) ;
  assign n10585 = ( ~n10574 & n10583 ) | ( ~n10574 & n10584 ) | ( n10583 & n10584 ) ;
  assign n10586 = ( n10543 & ~n10548 ) | ( n10543 & n10550 ) | ( ~n10548 & n10550 ) ;
  assign n10587 = ( n5414 & n10549 ) | ( n5414 & ~n10586 ) | ( n10549 & ~n10586 ) ;
  assign n10588 = n5914 & n10291 ;
  assign n10589 = x14 & n10588 ;
  assign n10590 = n6332 & ~n10279 ;
  assign n10591 = n5909 & n10281 ;
  assign n10592 = n10590 | n10591 ;
  assign n10593 = n5915 | n10592 ;
  assign n10594 = ( n10454 & n10592 ) | ( n10454 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10595 = x14 & ~n10594 ;
  assign n10596 = ( ~x14 & n10588 ) | ( ~x14 & n10594 ) | ( n10588 & n10594 ) ;
  assign n10597 = ( ~n10589 & n10595 ) | ( ~n10589 & n10596 ) | ( n10595 & n10596 ) ;
  assign n10598 = n5418 & n10283 ;
  assign n10599 = n5584 & ~n10285 ;
  assign n10600 = ( ~n10285 & n10598 ) | ( ~n10285 & n10599 ) | ( n10598 & n10599 ) ;
  assign n10601 = ( n5414 & n5417 ) | ( n5414 & n10285 ) | ( n5417 & n10285 ) ;
  assign n10602 = ~n10283 & n10601 ;
  assign n10603 = n10600 | n10602 ;
  assign n10604 = x17 & n5414 ;
  assign n10605 = ~n10285 & n10604 ;
  assign n10606 = ~n10603 & n10605 ;
  assign n10607 = n10603 & ~n10605 ;
  assign n10608 = n10606 | n10607 ;
  assign n10609 = ( ~n10587 & n10597 ) | ( ~n10587 & n10608 ) | ( n10597 & n10608 ) ;
  assign n10610 = ( n10587 & n10597 ) | ( n10587 & n10608 ) | ( n10597 & n10608 ) ;
  assign n10611 = ( n10587 & n10609 ) | ( n10587 & ~n10610 ) | ( n10609 & ~n10610 ) ;
  assign n10612 = ( n10572 & n10585 ) | ( n10572 & n10611 ) | ( n10585 & n10611 ) ;
  assign n10613 = n6796 & n10273 ;
  assign n10614 = x11 & n10613 ;
  assign n10615 = n10297 & ~n10341 ;
  assign n10616 = ( ~n10295 & n10297 ) | ( ~n10295 & n10341 ) | ( n10297 & n10341 ) ;
  assign n10617 = ( ~n10298 & n10615 ) | ( ~n10298 & n10616 ) | ( n10615 & n10616 ) ;
  assign n10618 = n6567 & n10275 ;
  assign n10619 = n6570 | n10618 ;
  assign n10620 = ( ~n10297 & n10618 ) | ( ~n10297 & n10619 ) | ( n10618 & n10619 ) ;
  assign n10621 = n6571 | n10620 ;
  assign n10622 = ( ~n10617 & n10620 ) | ( ~n10617 & n10621 ) | ( n10620 & n10621 ) ;
  assign n10623 = x11 & ~n10622 ;
  assign n10624 = ( ~x11 & n10613 ) | ( ~x11 & n10622 ) | ( n10613 & n10622 ) ;
  assign n10625 = ( ~n10614 & n10623 ) | ( ~n10614 & n10624 ) | ( n10623 & n10624 ) ;
  assign n10626 = n6332 & n10291 ;
  assign n10627 = x14 & n10626 ;
  assign n10628 = n5909 & ~n10279 ;
  assign n10629 = n5914 | n10628 ;
  assign n10630 = ( n10277 & n10628 ) | ( n10277 & n10629 ) | ( n10628 & n10629 ) ;
  assign n10631 = n5915 | n10630 ;
  assign n10632 = ( ~n10516 & n10630 ) | ( ~n10516 & n10631 ) | ( n10630 & n10631 ) ;
  assign n10633 = x14 & ~n10632 ;
  assign n10634 = ( ~x14 & n10626 ) | ( ~x14 & n10632 ) | ( n10626 & n10632 ) ;
  assign n10635 = ( ~n10627 & n10633 ) | ( ~n10627 & n10634 ) | ( n10633 & n10634 ) ;
  assign n10636 = n10603 | n10605 ;
  assign n10637 = x17 & ~n10636 ;
  assign n10638 = n5418 & n10464 ;
  assign n10639 = n5417 & n10281 ;
  assign n10640 = n5584 & ~n10283 ;
  assign n10641 = n5413 & ~n10285 ;
  assign n10642 = n10640 | n10641 ;
  assign n10643 = n10639 | n10642 ;
  assign n10644 = n10638 | n10643 ;
  assign n10645 = n10637 & ~n10644 ;
  assign n10646 = ( x17 & n10644 ) | ( x17 & ~n10645 ) | ( n10644 & ~n10645 ) ;
  assign n10647 = ( x17 & n10637 ) | ( x17 & n10644 ) | ( n10637 & n10644 ) ;
  assign n10648 = ( n10637 & n10646 ) | ( n10637 & ~n10647 ) | ( n10646 & ~n10647 ) ;
  assign n10649 = ( ~n10610 & n10635 ) | ( ~n10610 & n10648 ) | ( n10635 & n10648 ) ;
  assign n10650 = ( n10610 & n10635 ) | ( n10610 & n10648 ) | ( n10635 & n10648 ) ;
  assign n10651 = ( n10610 & n10649 ) | ( n10610 & ~n10650 ) | ( n10649 & ~n10650 ) ;
  assign n10652 = ( n10612 & n10625 ) | ( n10612 & n10651 ) | ( n10625 & n10651 ) ;
  assign n10653 = ( n10271 & n10298 ) | ( n10271 & n10342 ) | ( n10298 & n10342 ) ;
  assign n10654 = n10271 | n10298 ;
  assign n10655 = ( ~n10271 & n10298 ) | ( ~n10271 & n10342 ) | ( n10298 & n10342 ) ;
  assign n10656 = ( ~n10653 & n10654 ) | ( ~n10653 & n10655 ) | ( n10654 & n10655 ) ;
  assign n10657 = n6571 & ~n10656 ;
  assign n10658 = x11 & n10657 ;
  assign n10659 = n6567 & n10273 ;
  assign n10660 = n6570 | n10659 ;
  assign n10661 = ( n10271 & n10659 ) | ( n10271 & n10660 ) | ( n10659 & n10660 ) ;
  assign n10662 = n6796 & ~n10297 ;
  assign n10663 = n10661 | n10662 ;
  assign n10664 = x11 & ~n10663 ;
  assign n10665 = ( ~x11 & n10657 ) | ( ~x11 & n10663 ) | ( n10657 & n10663 ) ;
  assign n10666 = ( ~n10658 & n10664 ) | ( ~n10658 & n10665 ) | ( n10664 & n10665 ) ;
  assign n10667 = n6332 & n10277 ;
  assign n10668 = x14 & n10667 ;
  assign n10669 = n5909 & n10291 ;
  assign n10670 = n5914 | n10669 ;
  assign n10671 = ( n10275 & n10669 ) | ( n10275 & n10670 ) | ( n10669 & n10670 ) ;
  assign n10672 = n5915 | n10671 ;
  assign n10673 = ( n10563 & n10671 ) | ( n10563 & n10672 ) | ( n10671 & n10672 ) ;
  assign n10674 = x14 & ~n10673 ;
  assign n10675 = ( ~x14 & n10667 ) | ( ~x14 & n10673 ) | ( n10667 & n10673 ) ;
  assign n10676 = ( ~n10668 & n10674 ) | ( ~n10668 & n10675 ) | ( n10674 & n10675 ) ;
  assign n10677 = n5584 & n10281 ;
  assign n10678 = x17 & n10677 ;
  assign n10679 = n5413 & ~n10283 ;
  assign n10680 = n5417 | n10679 ;
  assign n10681 = ( ~n10279 & n10679 ) | ( ~n10279 & n10680 ) | ( n10679 & n10680 ) ;
  assign n10682 = n5418 | n10681 ;
  assign n10683 = ( n10487 & n10681 ) | ( n10487 & n10682 ) | ( n10681 & n10682 ) ;
  assign n10684 = x17 & ~n10683 ;
  assign n10685 = ( ~x17 & n10677 ) | ( ~x17 & n10683 ) | ( n10677 & n10683 ) ;
  assign n10686 = ( ~n10678 & n10684 ) | ( ~n10678 & n10685 ) | ( n10684 & n10685 ) ;
  assign n10687 = n4875 & ~n10285 ;
  assign n10688 = ( n10645 & ~n10686 ) | ( n10645 & n10687 ) | ( ~n10686 & n10687 ) ;
  assign n10689 = n10645 | n10687 ;
  assign n10690 = n10686 & n10689 ;
  assign n10691 = ( n10686 & n10688 ) | ( n10686 & ~n10690 ) | ( n10688 & ~n10690 ) ;
  assign n10692 = ( ~n10650 & n10676 ) | ( ~n10650 & n10691 ) | ( n10676 & n10691 ) ;
  assign n10693 = ( n10650 & n10676 ) | ( n10650 & n10691 ) | ( n10676 & n10691 ) ;
  assign n10694 = ( n10650 & n10692 ) | ( n10650 & ~n10693 ) | ( n10692 & ~n10693 ) ;
  assign n10695 = ( n10652 & n10666 ) | ( n10652 & n10694 ) | ( n10666 & n10694 ) ;
  assign n10696 = n10269 & ~n10343 ;
  assign n10697 = ( n10269 & ~n10299 ) | ( n10269 & n10343 ) | ( ~n10299 & n10343 ) ;
  assign n10698 = ( ~n10300 & n10696 ) | ( ~n10300 & n10697 ) | ( n10696 & n10697 ) ;
  assign n10699 = n6570 & ~n10269 ;
  assign n10700 = n6571 | n10699 ;
  assign n10701 = ( ~n10698 & n10699 ) | ( ~n10698 & n10700 ) | ( n10699 & n10700 ) ;
  assign n10702 = n6567 & ~n10297 ;
  assign n10703 = ( ~x11 & n10701 ) | ( ~x11 & n10702 ) | ( n10701 & n10702 ) ;
  assign n10704 = n6796 & n10271 ;
  assign n10705 = x11 & ~n10702 ;
  assign n10706 = n10704 | n10705 ;
  assign n10707 = ( n10701 & n10704 ) | ( n10701 & n10705 ) | ( n10704 & n10705 ) ;
  assign n10708 = ( n10703 & n10706 ) | ( n10703 & ~n10707 ) | ( n10706 & ~n10707 ) ;
  assign n10709 = n6332 & n10275 ;
  assign n10710 = x14 & n10709 ;
  assign n10711 = n5909 & n10277 ;
  assign n10712 = n5914 | n10711 ;
  assign n10713 = ( n10273 & n10711 ) | ( n10273 & n10712 ) | ( n10711 & n10712 ) ;
  assign n10714 = n5915 | n10713 ;
  assign n10715 = ( n10577 & n10713 ) | ( n10577 & n10714 ) | ( n10713 & n10714 ) ;
  assign n10716 = x14 & ~n10715 ;
  assign n10717 = ( ~x14 & n10709 ) | ( ~x14 & n10715 ) | ( n10709 & n10715 ) ;
  assign n10718 = ( ~n10710 & n10716 ) | ( ~n10710 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10719 = n5417 & n10291 ;
  assign n10720 = x17 & n10719 ;
  assign n10721 = n5584 & ~n10279 ;
  assign n10722 = n5413 & n10281 ;
  assign n10723 = n10721 | n10722 ;
  assign n10724 = n5418 | n10723 ;
  assign n10725 = ( n10454 & n10723 ) | ( n10454 & n10724 ) | ( n10723 & n10724 ) ;
  assign n10726 = x17 & ~n10725 ;
  assign n10727 = ( ~x17 & n10719 ) | ( ~x17 & n10725 ) | ( n10719 & n10725 ) ;
  assign n10728 = ( ~n10720 & n10726 ) | ( ~n10720 & n10727 ) | ( n10726 & n10727 ) ;
  assign n10729 = ( n5232 & n7364 ) | ( n5232 & n10283 ) | ( n7364 & n10283 ) ;
  assign n10730 = ~n10285 & n10729 ;
  assign n10731 = n4875 & n10286 ;
  assign n10732 = n10730 | n10731 ;
  assign n10733 = n4878 & ~n10283 ;
  assign n10734 = n10732 | n10733 ;
  assign n10735 = x20 & n10687 ;
  assign n10736 = ~n10734 & n10735 ;
  assign n10737 = n10734 & ~n10735 ;
  assign n10738 = n10736 | n10737 ;
  assign n10739 = ( n10690 & n10728 ) | ( n10690 & n10738 ) | ( n10728 & n10738 ) ;
  assign n10740 = ( n10690 & ~n10728 ) | ( n10690 & n10738 ) | ( ~n10728 & n10738 ) ;
  assign n10741 = ( n10728 & ~n10739 ) | ( n10728 & n10740 ) | ( ~n10739 & n10740 ) ;
  assign n10742 = ( ~n10693 & n10718 ) | ( ~n10693 & n10741 ) | ( n10718 & n10741 ) ;
  assign n10743 = ( n10693 & n10718 ) | ( n10693 & n10741 ) | ( n10718 & n10741 ) ;
  assign n10744 = ( n10693 & n10742 ) | ( n10693 & ~n10743 ) | ( n10742 & ~n10743 ) ;
  assign n10745 = ( n10695 & n10708 ) | ( n10695 & n10744 ) | ( n10708 & n10744 ) ;
  assign n10746 = n6332 & n10273 ;
  assign n10747 = x14 & n10746 ;
  assign n10748 = n5909 & n10275 ;
  assign n10749 = n5914 | n10748 ;
  assign n10750 = ( ~n10297 & n10748 ) | ( ~n10297 & n10749 ) | ( n10748 & n10749 ) ;
  assign n10751 = n5915 | n10750 ;
  assign n10752 = ( ~n10617 & n10750 ) | ( ~n10617 & n10751 ) | ( n10750 & n10751 ) ;
  assign n10753 = x14 & ~n10752 ;
  assign n10754 = ( ~x14 & n10746 ) | ( ~x14 & n10752 ) | ( n10746 & n10752 ) ;
  assign n10755 = ( ~n10747 & n10753 ) | ( ~n10747 & n10754 ) | ( n10753 & n10754 ) ;
  assign n10756 = n5584 & n10291 ;
  assign n10757 = x17 & n10756 ;
  assign n10758 = n5413 & ~n10279 ;
  assign n10759 = n5417 | n10758 ;
  assign n10760 = ( n10277 & n10758 ) | ( n10277 & n10759 ) | ( n10758 & n10759 ) ;
  assign n10761 = n5418 | n10760 ;
  assign n10762 = ( ~n10516 & n10760 ) | ( ~n10516 & n10761 ) | ( n10760 & n10761 ) ;
  assign n10763 = x17 & ~n10762 ;
  assign n10764 = ( ~x17 & n10756 ) | ( ~x17 & n10762 ) | ( n10756 & n10762 ) ;
  assign n10765 = ( ~n10757 & n10763 ) | ( ~n10757 & n10764 ) | ( n10763 & n10764 ) ;
  assign n10766 = n4879 & n10464 ;
  assign n10767 = n4878 & n10281 ;
  assign n10768 = n5232 & ~n10283 ;
  assign n10769 = n4874 & ~n10285 ;
  assign n10770 = n10768 | n10769 ;
  assign n10771 = n10767 | n10770 ;
  assign n10772 = n10766 | n10771 ;
  assign n10773 = ~x20 & n10772 ;
  assign n10774 = x20 & ~n10687 ;
  assign n10775 = ~n10734 & n10774 ;
  assign n10776 = ( x20 & n10772 ) | ( x20 & ~n10775 ) | ( n10772 & ~n10775 ) ;
  assign n10777 = n10772 & ~n10775 ;
  assign n10778 = ( n10773 & n10776 ) | ( n10773 & ~n10777 ) | ( n10776 & ~n10777 ) ;
  assign n10779 = ( ~n10739 & n10765 ) | ( ~n10739 & n10778 ) | ( n10765 & n10778 ) ;
  assign n10780 = ( n10739 & n10765 ) | ( n10739 & n10778 ) | ( n10765 & n10778 ) ;
  assign n10781 = ( n10739 & n10779 ) | ( n10739 & ~n10780 ) | ( n10779 & ~n10780 ) ;
  assign n10782 = ( ~n10743 & n10755 ) | ( ~n10743 & n10781 ) | ( n10755 & n10781 ) ;
  assign n10783 = ( n10743 & n10755 ) | ( n10743 & n10781 ) | ( n10755 & n10781 ) ;
  assign n10784 = ( n10743 & n10782 ) | ( n10743 & ~n10783 ) | ( n10782 & ~n10783 ) ;
  assign n10785 = n10267 & n10344 ;
  assign n10786 = ( ~n10267 & n10300 ) | ( ~n10267 & n10344 ) | ( n10300 & n10344 ) ;
  assign n10787 = ( n10301 & ~n10785 ) | ( n10301 & n10786 ) | ( ~n10785 & n10786 ) ;
  assign n10788 = n6571 & ~n10787 ;
  assign n10789 = x11 & n10788 ;
  assign n10790 = n6567 & n10271 ;
  assign n10791 = n6570 | n10790 ;
  assign n10792 = ( n10267 & n10790 ) | ( n10267 & n10791 ) | ( n10790 & n10791 ) ;
  assign n10793 = n6796 & ~n10269 ;
  assign n10794 = n10792 | n10793 ;
  assign n10795 = x11 & ~n10794 ;
  assign n10796 = ( ~x11 & n10788 ) | ( ~x11 & n10794 ) | ( n10788 & n10794 ) ;
  assign n10797 = ( ~n10789 & n10795 ) | ( ~n10789 & n10796 ) | ( n10795 & n10796 ) ;
  assign n10798 = ( n10745 & n10784 ) | ( n10745 & n10797 ) | ( n10784 & n10797 ) ;
  assign n10799 = n6796 & n10267 ;
  assign n10800 = x11 & n10799 ;
  assign n10801 = n10265 & ~n10345 ;
  assign n10802 = ( n10265 & ~n10301 ) | ( n10265 & n10345 ) | ( ~n10301 & n10345 ) ;
  assign n10803 = n10265 & ~n10301 ;
  assign n10804 = ( n10801 & n10802 ) | ( n10801 & ~n10803 ) | ( n10802 & ~n10803 ) ;
  assign n10805 = n6567 & ~n10269 ;
  assign n10806 = n6570 | n10805 ;
  assign n10807 = ( n10265 & n10805 ) | ( n10265 & n10806 ) | ( n10805 & n10806 ) ;
  assign n10808 = n6571 | n10807 ;
  assign n10809 = ( n10804 & n10807 ) | ( n10804 & n10808 ) | ( n10807 & n10808 ) ;
  assign n10810 = x11 & ~n10809 ;
  assign n10811 = ( ~x11 & n10799 ) | ( ~x11 & n10809 ) | ( n10799 & n10809 ) ;
  assign n10812 = ( ~n10800 & n10810 ) | ( ~n10800 & n10811 ) | ( n10810 & n10811 ) ;
  assign n10813 = n6332 & ~n10297 ;
  assign n10814 = x14 & n10813 ;
  assign n10815 = n5909 & n10273 ;
  assign n10816 = n5914 | n10815 ;
  assign n10817 = ( n10271 & n10815 ) | ( n10271 & n10816 ) | ( n10815 & n10816 ) ;
  assign n10818 = n5915 | n10817 ;
  assign n10819 = ( ~n10656 & n10817 ) | ( ~n10656 & n10818 ) | ( n10817 & n10818 ) ;
  assign n10820 = x14 & ~n10819 ;
  assign n10821 = ( ~x14 & n10813 ) | ( ~x14 & n10819 ) | ( n10813 & n10819 ) ;
  assign n10822 = ( ~n10814 & n10820 ) | ( ~n10814 & n10821 ) | ( n10820 & n10821 ) ;
  assign n10823 = n5584 & n10277 ;
  assign n10824 = x17 & n10823 ;
  assign n10825 = n5413 & n10291 ;
  assign n10826 = n5417 | n10825 ;
  assign n10827 = ( n10275 & n10825 ) | ( n10275 & n10826 ) | ( n10825 & n10826 ) ;
  assign n10828 = n5418 | n10827 ;
  assign n10829 = ( n10563 & n10827 ) | ( n10563 & n10828 ) | ( n10827 & n10828 ) ;
  assign n10830 = x17 & ~n10829 ;
  assign n10831 = ( ~x17 & n10823 ) | ( ~x17 & n10829 ) | ( n10823 & n10829 ) ;
  assign n10832 = ( ~n10824 & n10830 ) | ( ~n10824 & n10831 ) | ( n10830 & n10831 ) ;
  assign n10833 = x21 | n10285 ;
  assign n10834 = n4879 & n10487 ;
  assign n10835 = n4878 & ~n10279 ;
  assign n10836 = n5232 & n10281 ;
  assign n10837 = n4874 & ~n10283 ;
  assign n10838 = n10836 | n10837 ;
  assign n10839 = n10835 | n10838 ;
  assign n10840 = n10834 | n10839 ;
  assign n10841 = ~n10772 & n10775 ;
  assign n10842 = ~x20 & n10285 ;
  assign n10843 = n10841 | n10842 ;
  assign n10844 = ( ~n10833 & n10840 ) | ( ~n10833 & n10843 ) | ( n10840 & n10843 ) ;
  assign n10845 = ( n10833 & n10840 ) | ( n10833 & n10843 ) | ( n10840 & n10843 ) ;
  assign n10846 = ( n10833 & n10844 ) | ( n10833 & ~n10845 ) | ( n10844 & ~n10845 ) ;
  assign n10847 = ( ~n10780 & n10832 ) | ( ~n10780 & n10846 ) | ( n10832 & n10846 ) ;
  assign n10848 = ( n10780 & n10832 ) | ( n10780 & n10846 ) | ( n10832 & n10846 ) ;
  assign n10849 = ( n10780 & n10847 ) | ( n10780 & ~n10848 ) | ( n10847 & ~n10848 ) ;
  assign n10850 = ( ~n10783 & n10822 ) | ( ~n10783 & n10849 ) | ( n10822 & n10849 ) ;
  assign n10851 = ( n10783 & n10822 ) | ( n10783 & n10849 ) | ( n10822 & n10849 ) ;
  assign n10852 = ( n10783 & n10850 ) | ( n10783 & ~n10851 ) | ( n10850 & ~n10851 ) ;
  assign n10853 = ( ~n10798 & n10812 ) | ( ~n10798 & n10852 ) | ( n10812 & n10852 ) ;
  assign n10854 = ( n10798 & n10812 ) | ( n10798 & n10852 ) | ( n10812 & n10852 ) ;
  assign n10855 = ( n10798 & n10853 ) | ( n10798 & ~n10854 ) | ( n10853 & ~n10854 ) ;
  assign n10856 = ( n10259 & ~n10304 ) | ( n10259 & n10348 ) | ( ~n10304 & n10348 ) ;
  assign n10857 = ~n10259 & n10304 ;
  assign n10858 = ( n10259 & n10304 ) | ( n10259 & ~n10348 ) | ( n10304 & ~n10348 ) ;
  assign n10859 = ( n10856 & n10857 ) | ( n10856 & n10858 ) | ( n10857 & n10858 ) ;
  assign n10860 = n7346 & n10859 ;
  assign n10861 = x8 & n10860 ;
  assign n10862 = n7341 & n10263 ;
  assign n10863 = n7345 | n10862 ;
  assign n10864 = ( n10259 & n10862 ) | ( n10259 & n10863 ) | ( n10862 & n10863 ) ;
  assign n10865 = n7644 & n10261 ;
  assign n10866 = n10864 | n10865 ;
  assign n10867 = x8 & ~n10866 ;
  assign n10868 = ( ~x8 & n10860 ) | ( ~x8 & n10866 ) | ( n10860 & n10866 ) ;
  assign n10869 = ( ~n10861 & n10867 ) | ( ~n10861 & n10868 ) | ( n10867 & n10868 ) ;
  assign n10870 = ( ~n10695 & n10708 ) | ( ~n10695 & n10744 ) | ( n10708 & n10744 ) ;
  assign n10871 = ( n10695 & ~n10745 ) | ( n10695 & n10870 ) | ( ~n10745 & n10870 ) ;
  assign n10872 = n10302 & ~n10347 ;
  assign n10873 = ( ~n10265 & n10303 ) | ( ~n10265 & n10801 ) | ( n10303 & n10801 ) ;
  assign n10874 = ( n10263 & n10872 ) | ( n10263 & ~n10873 ) | ( n10872 & ~n10873 ) ;
  assign n10875 = n7346 & n10874 ;
  assign n10876 = x8 & n10875 ;
  assign n10877 = n7341 & n10267 ;
  assign n10878 = n7345 | n10877 ;
  assign n10879 = ( n10263 & n10877 ) | ( n10263 & n10878 ) | ( n10877 & n10878 ) ;
  assign n10880 = n7644 & n10265 ;
  assign n10881 = n10879 | n10880 ;
  assign n10882 = x8 & ~n10881 ;
  assign n10883 = ( ~x8 & n10875 ) | ( ~x8 & n10881 ) | ( n10875 & n10881 ) ;
  assign n10884 = ( ~n10876 & n10882 ) | ( ~n10876 & n10883 ) | ( n10882 & n10883 ) ;
  assign n10885 = n7345 & n10291 ;
  assign n10886 = x8 & n10885 ;
  assign n10887 = n7644 & ~n10279 ;
  assign n10888 = n7341 & n10281 ;
  assign n10889 = n10887 | n10888 ;
  assign n10890 = n7346 | n10889 ;
  assign n10891 = ( n10454 & n10889 ) | ( n10454 & n10890 ) | ( n10889 & n10890 ) ;
  assign n10892 = x8 & ~n10891 ;
  assign n10893 = ( ~x8 & n10885 ) | ( ~x8 & n10891 ) | ( n10885 & n10891 ) ;
  assign n10894 = ( ~n10886 & n10892 ) | ( ~n10886 & n10893 ) | ( n10892 & n10893 ) ;
  assign n10895 = x11 & n10478 ;
  assign n10896 = ~n10477 & n10895 ;
  assign n10897 = n10477 & ~n10895 ;
  assign n10898 = n10896 | n10897 ;
  assign n10899 = n7644 & n10281 ;
  assign n10900 = x8 & n10899 ;
  assign n10901 = n7341 & ~n10283 ;
  assign n10902 = n7345 | n10901 ;
  assign n10903 = ( ~n10279 & n10901 ) | ( ~n10279 & n10902 ) | ( n10901 & n10902 ) ;
  assign n10904 = n7346 | n10903 ;
  assign n10905 = ( n10487 & n10903 ) | ( n10487 & n10904 ) | ( n10903 & n10904 ) ;
  assign n10906 = x8 & ~n10905 ;
  assign n10907 = ( ~x8 & n10899 ) | ( ~x8 & n10905 ) | ( n10899 & n10905 ) ;
  assign n10908 = ( ~n10900 & n10906 ) | ( ~n10900 & n10907 ) | ( n10906 & n10907 ) ;
  assign n10909 = n10478 & n10908 ;
  assign n10910 = ( n7644 & n8768 ) | ( n7644 & n10283 ) | ( n8768 & n10283 ) ;
  assign n10911 = ~n10285 & n10910 ;
  assign n10912 = n7342 & n10286 ;
  assign n10913 = n10911 | n10912 ;
  assign n10914 = n7345 & ~n10283 ;
  assign n10915 = n10913 | n10914 ;
  assign n10916 = n7342 & ~n10285 ;
  assign n10917 = x8 & n10916 ;
  assign n10918 = n10915 | n10917 ;
  assign n10919 = x8 & ~n10918 ;
  assign n10920 = n7346 & n10464 ;
  assign n10921 = n7345 & n10281 ;
  assign n10922 = n7644 & ~n10283 ;
  assign n10923 = n7341 & ~n10285 ;
  assign n10924 = n10922 | n10923 ;
  assign n10925 = n10921 | n10924 ;
  assign n10926 = n10920 | n10925 ;
  assign n10927 = n10919 & ~n10926 ;
  assign n10928 = ( n10478 & n10908 ) | ( n10478 & ~n10927 ) | ( n10908 & ~n10927 ) ;
  assign n10929 = ( n10478 & ~n10908 ) | ( n10478 & n10927 ) | ( ~n10908 & n10927 ) ;
  assign n10930 = ( ~n10909 & n10928 ) | ( ~n10909 & n10929 ) | ( n10928 & n10929 ) ;
  assign n10931 = ( n10908 & n10909 ) | ( n10908 & ~n10930 ) | ( n10909 & ~n10930 ) ;
  assign n10932 = ( n10894 & n10898 ) | ( n10894 & n10931 ) | ( n10898 & n10931 ) ;
  assign n10933 = n7346 & ~n10516 ;
  assign n10934 = x8 & n10933 ;
  assign n10935 = n7341 & ~n10279 ;
  assign n10936 = n7345 | n10935 ;
  assign n10937 = ( n10277 & n10935 ) | ( n10277 & n10936 ) | ( n10935 & n10936 ) ;
  assign n10938 = n7644 & n10291 ;
  assign n10939 = n10937 | n10938 ;
  assign n10940 = x8 & ~n10939 ;
  assign n10941 = ( ~x8 & n10933 ) | ( ~x8 & n10939 ) | ( n10933 & n10939 ) ;
  assign n10942 = ( ~n10934 & n10940 ) | ( ~n10934 & n10941 ) | ( n10940 & n10941 ) ;
  assign n10943 = x11 & ~n10480 ;
  assign n10944 = ~n10471 & n10943 ;
  assign n10945 = n10471 & ~n10943 ;
  assign n10946 = n10944 | n10945 ;
  assign n10947 = ( n10932 & n10942 ) | ( n10932 & n10946 ) | ( n10942 & n10946 ) ;
  assign n10948 = n7644 & n10277 ;
  assign n10949 = x8 & n10948 ;
  assign n10950 = n7341 & n10291 ;
  assign n10951 = n7345 | n10950 ;
  assign n10952 = ( n10275 & n10950 ) | ( n10275 & n10951 ) | ( n10950 & n10951 ) ;
  assign n10953 = n7346 | n10952 ;
  assign n10954 = ( n10563 & n10952 ) | ( n10563 & n10953 ) | ( n10952 & n10953 ) ;
  assign n10955 = x8 & ~n10954 ;
  assign n10956 = ( ~x8 & n10948 ) | ( ~x8 & n10954 ) | ( n10948 & n10954 ) ;
  assign n10957 = ( ~n10949 & n10955 ) | ( ~n10949 & n10956 ) | ( n10955 & n10956 ) ;
  assign n10958 = x12 | n10285 ;
  assign n10959 = ~x11 & n10285 ;
  assign n10960 = n10481 | n10959 ;
  assign n10961 = ( ~n10494 & n10958 ) | ( ~n10494 & n10960 ) | ( n10958 & n10960 ) ;
  assign n10962 = ( n10494 & n10958 ) | ( n10494 & n10960 ) | ( n10958 & n10960 ) ;
  assign n10963 = ( n10494 & n10961 ) | ( n10494 & ~n10962 ) | ( n10961 & ~n10962 ) ;
  assign n10964 = ( n10947 & n10957 ) | ( n10947 & n10963 ) | ( n10957 & n10963 ) ;
  assign n10965 = n7346 & n10577 ;
  assign n10966 = x8 & n10965 ;
  assign n10967 = n7341 & n10277 ;
  assign n10968 = n7345 | n10967 ;
  assign n10969 = ( n10273 & n10967 ) | ( n10273 & n10968 ) | ( n10967 & n10968 ) ;
  assign n10970 = n7644 & n10275 ;
  assign n10971 = n10969 | n10970 ;
  assign n10972 = x8 & ~n10971 ;
  assign n10973 = ( ~x8 & n10965 ) | ( ~x8 & n10971 ) | ( n10965 & n10971 ) ;
  assign n10974 = ( ~n10966 & n10972 ) | ( ~n10966 & n10973 ) | ( n10972 & n10973 ) ;
  assign n10975 = ( ~n10462 & n10499 ) | ( ~n10462 & n10510 ) | ( n10499 & n10510 ) ;
  assign n10976 = ( n10462 & ~n10511 ) | ( n10462 & n10975 ) | ( ~n10511 & n10975 ) ;
  assign n10977 = ( n10964 & n10974 ) | ( n10964 & n10976 ) | ( n10974 & n10976 ) ;
  assign n10978 = n7644 & n10273 ;
  assign n10979 = x8 & n10978 ;
  assign n10980 = n7341 & n10275 ;
  assign n10981 = n7345 | n10980 ;
  assign n10982 = ( ~n10297 & n10980 ) | ( ~n10297 & n10981 ) | ( n10980 & n10981 ) ;
  assign n10983 = n7346 | n10982 ;
  assign n10984 = ( ~n10617 & n10982 ) | ( ~n10617 & n10983 ) | ( n10982 & n10983 ) ;
  assign n10985 = x8 & ~n10984 ;
  assign n10986 = ( ~x8 & n10978 ) | ( ~x8 & n10984 ) | ( n10978 & n10984 ) ;
  assign n10987 = ( ~n10979 & n10985 ) | ( ~n10979 & n10986 ) | ( n10985 & n10986 ) ;
  assign n10988 = ( ~n10511 & n10524 ) | ( ~n10511 & n10535 ) | ( n10524 & n10535 ) ;
  assign n10989 = ( n10511 & ~n10536 ) | ( n10511 & n10988 ) | ( ~n10536 & n10988 ) ;
  assign n10990 = ( n10977 & n10987 ) | ( n10977 & n10989 ) | ( n10987 & n10989 ) ;
  assign n10991 = ( ~n10536 & n10557 ) | ( ~n10536 & n10571 ) | ( n10557 & n10571 ) ;
  assign n10992 = ( n10536 & ~n10572 ) | ( n10536 & n10991 ) | ( ~n10572 & n10991 ) ;
  assign n10993 = n7644 & ~n10297 ;
  assign n10994 = x8 & n10993 ;
  assign n10995 = n7341 & n10273 ;
  assign n10996 = n7345 | n10995 ;
  assign n10997 = ( n10271 & n10995 ) | ( n10271 & n10996 ) | ( n10995 & n10996 ) ;
  assign n10998 = n7346 | n10997 ;
  assign n10999 = ( ~n10656 & n10997 ) | ( ~n10656 & n10998 ) | ( n10997 & n10998 ) ;
  assign n11000 = x8 & ~n10999 ;
  assign n11001 = ( ~x8 & n10993 ) | ( ~x8 & n10999 ) | ( n10993 & n10999 ) ;
  assign n11002 = ( ~n10994 & n11000 ) | ( ~n10994 & n11001 ) | ( n11000 & n11001 ) ;
  assign n11003 = ( n10990 & n10992 ) | ( n10990 & n11002 ) | ( n10992 & n11002 ) ;
  assign n11004 = ( ~n10572 & n10585 ) | ( ~n10572 & n10611 ) | ( n10585 & n10611 ) ;
  assign n11005 = ( n10572 & ~n10612 ) | ( n10572 & n11004 ) | ( ~n10612 & n11004 ) ;
  assign n11006 = n7644 & n10271 ;
  assign n11007 = x8 & n11006 ;
  assign n11008 = n7341 & ~n10297 ;
  assign n11009 = n7345 | n11008 ;
  assign n11010 = ( ~n10269 & n11008 ) | ( ~n10269 & n11009 ) | ( n11008 & n11009 ) ;
  assign n11011 = n7346 | n11010 ;
  assign n11012 = ( ~n10698 & n11010 ) | ( ~n10698 & n11011 ) | ( n11010 & n11011 ) ;
  assign n11013 = x8 & ~n11012 ;
  assign n11014 = ( ~x8 & n11006 ) | ( ~x8 & n11012 ) | ( n11006 & n11012 ) ;
  assign n11015 = ( ~n11007 & n11013 ) | ( ~n11007 & n11014 ) | ( n11013 & n11014 ) ;
  assign n11016 = ( n11003 & n11005 ) | ( n11003 & n11015 ) | ( n11005 & n11015 ) ;
  assign n11017 = ( ~n10612 & n10625 ) | ( ~n10612 & n10651 ) | ( n10625 & n10651 ) ;
  assign n11018 = ( n10612 & ~n10652 ) | ( n10612 & n11017 ) | ( ~n10652 & n11017 ) ;
  assign n11019 = n7346 & ~n10787 ;
  assign n11020 = x8 & n11019 ;
  assign n11021 = n7341 & n10271 ;
  assign n11022 = n7345 | n11021 ;
  assign n11023 = ( n10267 & n11021 ) | ( n10267 & n11022 ) | ( n11021 & n11022 ) ;
  assign n11024 = n7644 & ~n10269 ;
  assign n11025 = n11023 | n11024 ;
  assign n11026 = x8 & ~n11025 ;
  assign n11027 = ( ~x8 & n11019 ) | ( ~x8 & n11025 ) | ( n11019 & n11025 ) ;
  assign n11028 = ( ~n11020 & n11026 ) | ( ~n11020 & n11027 ) | ( n11026 & n11027 ) ;
  assign n11029 = ( n11016 & n11018 ) | ( n11016 & n11028 ) | ( n11018 & n11028 ) ;
  assign n11030 = ( ~n10652 & n10666 ) | ( ~n10652 & n10694 ) | ( n10666 & n10694 ) ;
  assign n11031 = ( n10652 & ~n10695 ) | ( n10652 & n11030 ) | ( ~n10695 & n11030 ) ;
  assign n11032 = n7644 & n10267 ;
  assign n11033 = x8 & n11032 ;
  assign n11034 = n7341 & ~n10269 ;
  assign n11035 = n7345 | n11034 ;
  assign n11036 = ( n10265 & n11034 ) | ( n10265 & n11035 ) | ( n11034 & n11035 ) ;
  assign n11037 = n7346 | n11036 ;
  assign n11038 = ( n10804 & n11036 ) | ( n10804 & n11037 ) | ( n11036 & n11037 ) ;
  assign n11039 = x8 & ~n11038 ;
  assign n11040 = ( ~x8 & n11032 ) | ( ~x8 & n11038 ) | ( n11032 & n11038 ) ;
  assign n11041 = ( ~n11033 & n11039 ) | ( ~n11033 & n11040 ) | ( n11039 & n11040 ) ;
  assign n11042 = ( n11029 & n11031 ) | ( n11029 & n11041 ) | ( n11031 & n11041 ) ;
  assign n11043 = ( n10871 & n10884 ) | ( n10871 & n11042 ) | ( n10884 & n11042 ) ;
  assign n11044 = ( ~n10745 & n10784 ) | ( ~n10745 & n10797 ) | ( n10784 & n10797 ) ;
  assign n11045 = ( n10745 & ~n10798 ) | ( n10745 & n11044 ) | ( ~n10798 & n11044 ) ;
  assign n11046 = ( n10261 & ~n10303 ) | ( n10261 & n10347 ) | ( ~n10303 & n10347 ) ;
  assign n11047 = n10261 & ~n10303 ;
  assign n11048 = ( n10261 & n10303 ) | ( n10261 & ~n10347 ) | ( n10303 & ~n10347 ) ;
  assign n11049 = ( n11046 & ~n11047 ) | ( n11046 & n11048 ) | ( ~n11047 & n11048 ) ;
  assign n11050 = n7346 & n11049 ;
  assign n11051 = x8 & n11050 ;
  assign n11052 = n7341 & n10265 ;
  assign n11053 = n7345 | n11052 ;
  assign n11054 = ( n10261 & n11052 ) | ( n10261 & n11053 ) | ( n11052 & n11053 ) ;
  assign n11055 = n7644 & n10263 ;
  assign n11056 = n11054 | n11055 ;
  assign n11057 = x8 & ~n11056 ;
  assign n11058 = ( ~x8 & n11050 ) | ( ~x8 & n11056 ) | ( n11050 & n11056 ) ;
  assign n11059 = ( ~n11051 & n11057 ) | ( ~n11051 & n11058 ) | ( n11057 & n11058 ) ;
  assign n11060 = ( n11043 & n11045 ) | ( n11043 & n11059 ) | ( n11045 & n11059 ) ;
  assign n11061 = ( n10855 & n10869 ) | ( n10855 & n11060 ) | ( n10869 & n11060 ) ;
  assign n11062 = ( n10257 & ~n10305 ) | ( n10257 & n10349 ) | ( ~n10305 & n10349 ) ;
  assign n11063 = n10257 & ~n10305 ;
  assign n11064 = ( n10257 & n10305 ) | ( n10257 & ~n10349 ) | ( n10305 & ~n10349 ) ;
  assign n11065 = ( n11062 & ~n11063 ) | ( n11062 & n11064 ) | ( ~n11063 & n11064 ) ;
  assign n11066 = n7346 & n11065 ;
  assign n11067 = x8 & n11066 ;
  assign n11068 = n7341 & n10261 ;
  assign n11069 = n7345 | n11068 ;
  assign n11070 = ( n10257 & n11068 ) | ( n10257 & n11069 ) | ( n11068 & n11069 ) ;
  assign n11071 = n7644 & n10259 ;
  assign n11072 = n11070 | n11071 ;
  assign n11073 = x8 & ~n11072 ;
  assign n11074 = ( ~x8 & n11066 ) | ( ~x8 & n11072 ) | ( n11066 & n11072 ) ;
  assign n11075 = ( ~n11067 & n11073 ) | ( ~n11067 & n11074 ) | ( n11073 & n11074 ) ;
  assign n11076 = n6571 & n10874 ;
  assign n11077 = x11 & n11076 ;
  assign n11078 = n6567 & n10267 ;
  assign n11079 = n6570 | n11078 ;
  assign n11080 = ( n10263 & n11078 ) | ( n10263 & n11079 ) | ( n11078 & n11079 ) ;
  assign n11081 = n6796 & n10265 ;
  assign n11082 = n11080 | n11081 ;
  assign n11083 = x11 & ~n11082 ;
  assign n11084 = ( ~x11 & n11076 ) | ( ~x11 & n11082 ) | ( n11076 & n11082 ) ;
  assign n11085 = ( ~n11077 & n11083 ) | ( ~n11077 & n11084 ) | ( n11083 & n11084 ) ;
  assign n11086 = n5584 & n10275 ;
  assign n11087 = x17 & n11086 ;
  assign n11088 = n5413 & n10277 ;
  assign n11089 = n5417 | n11088 ;
  assign n11090 = ( n10273 & n11088 ) | ( n10273 & n11089 ) | ( n11088 & n11089 ) ;
  assign n11091 = n5418 | n11090 ;
  assign n11092 = ( n10577 & n11090 ) | ( n10577 & n11091 ) | ( n11090 & n11091 ) ;
  assign n11093 = x17 & ~n11092 ;
  assign n11094 = ( ~x17 & n11086 ) | ( ~x17 & n11092 ) | ( n11086 & n11092 ) ;
  assign n11095 = ( ~n11087 & n11093 ) | ( ~n11087 & n11094 ) | ( n11093 & n11094 ) ;
  assign n11096 = n4878 & n10291 ;
  assign n11097 = x20 & n11096 ;
  assign n11098 = n5232 & ~n10279 ;
  assign n11099 = n4874 & n10281 ;
  assign n11100 = n11098 | n11099 ;
  assign n11101 = n4879 | n11100 ;
  assign n11102 = ( n10454 & n11100 ) | ( n10454 & n11101 ) | ( n11100 & n11101 ) ;
  assign n11103 = x20 & ~n11102 ;
  assign n11104 = ( ~x20 & n11096 ) | ( ~x20 & n11102 ) | ( n11096 & n11102 ) ;
  assign n11105 = ( ~n11097 & n11103 ) | ( ~n11097 & n11104 ) | ( n11103 & n11104 ) ;
  assign n11106 = x20 & ~n10833 ;
  assign n11107 = n10841 | n11106 ;
  assign n11108 = n4589 & ~n10285 ;
  assign n11109 = n10840 & n11108 ;
  assign n11110 = n10840 & ~n11108 ;
  assign n11111 = ( n11107 & n11109 ) | ( n11107 & ~n11110 ) | ( n11109 & ~n11110 ) ;
  assign n11112 = n4591 & n10283 ;
  assign n11113 = n4637 & ~n10285 ;
  assign n11114 = ( ~n10285 & n11112 ) | ( ~n10285 & n11113 ) | ( n11112 & n11113 ) ;
  assign n11115 = ( n4590 & n4649 ) | ( n4590 & n10285 ) | ( n4649 & n10285 ) ;
  assign n11116 = ~n10283 & n11115 ;
  assign n11117 = n11114 | n11116 ;
  assign n11118 = n4590 & ~n10285 ;
  assign n11119 = n11117 | n11118 ;
  assign n11120 = ( x23 & ~n11117 ) | ( x23 & n11118 ) | ( ~n11117 & n11118 ) ;
  assign n11121 = x23 & ~n11117 ;
  assign n11122 = ( n11119 & ~n11120 ) | ( n11119 & n11121 ) | ( ~n11120 & n11121 ) ;
  assign n11123 = ( ~n11105 & n11111 ) | ( ~n11105 & n11122 ) | ( n11111 & n11122 ) ;
  assign n11124 = ( n11105 & n11111 ) | ( n11105 & n11122 ) | ( n11111 & n11122 ) ;
  assign n11125 = ( n11105 & n11123 ) | ( n11105 & ~n11124 ) | ( n11123 & ~n11124 ) ;
  assign n11126 = ( ~n10848 & n11095 ) | ( ~n10848 & n11125 ) | ( n11095 & n11125 ) ;
  assign n11127 = ( n10848 & n11095 ) | ( n10848 & n11125 ) | ( n11095 & n11125 ) ;
  assign n11128 = ( n10848 & n11126 ) | ( n10848 & ~n11127 ) | ( n11126 & ~n11127 ) ;
  assign n11129 = n6332 & n10271 ;
  assign n11130 = x14 & n11129 ;
  assign n11131 = n5909 & ~n10297 ;
  assign n11132 = n5914 | n11131 ;
  assign n11133 = ( ~n10269 & n11131 ) | ( ~n10269 & n11132 ) | ( n11131 & n11132 ) ;
  assign n11134 = n5915 | n11133 ;
  assign n11135 = ( ~n10698 & n11133 ) | ( ~n10698 & n11134 ) | ( n11133 & n11134 ) ;
  assign n11136 = x14 & ~n11135 ;
  assign n11137 = ( ~x14 & n11129 ) | ( ~x14 & n11135 ) | ( n11129 & n11135 ) ;
  assign n11138 = ( ~n11130 & n11136 ) | ( ~n11130 & n11137 ) | ( n11136 & n11137 ) ;
  assign n11139 = ( ~n10851 & n11128 ) | ( ~n10851 & n11138 ) | ( n11128 & n11138 ) ;
  assign n11140 = ( n10851 & n11128 ) | ( n10851 & n11138 ) | ( n11128 & n11138 ) ;
  assign n11141 = ( n10851 & n11139 ) | ( n10851 & ~n11140 ) | ( n11139 & ~n11140 ) ;
  assign n11142 = ( ~n10854 & n11085 ) | ( ~n10854 & n11141 ) | ( n11085 & n11141 ) ;
  assign n11143 = ( n10854 & n11085 ) | ( n10854 & n11141 ) | ( n11085 & n11141 ) ;
  assign n11144 = ( n10854 & n11142 ) | ( n10854 & ~n11143 ) | ( n11142 & ~n11143 ) ;
  assign n11145 = ( n11061 & n11075 ) | ( n11061 & n11144 ) | ( n11075 & n11144 ) ;
  assign n11146 = n10255 & n10350 ;
  assign n11147 = ( n10255 & n10306 ) | ( n10255 & ~n10350 ) | ( n10306 & ~n10350 ) ;
  assign n11148 = ( ~n10307 & n11146 ) | ( ~n10307 & n11147 ) | ( n11146 & n11147 ) ;
  assign n11149 = n7346 & n11148 ;
  assign n11150 = x8 & n11149 ;
  assign n11151 = n7341 & n10259 ;
  assign n11152 = n7345 | n11151 ;
  assign n11153 = ( n10255 & n11151 ) | ( n10255 & n11152 ) | ( n11151 & n11152 ) ;
  assign n11154 = n7644 & n10257 ;
  assign n11155 = n11153 | n11154 ;
  assign n11156 = x8 & ~n11155 ;
  assign n11157 = ( ~x8 & n11149 ) | ( ~x8 & n11155 ) | ( n11149 & n11155 ) ;
  assign n11158 = ( ~n11150 & n11156 ) | ( ~n11150 & n11157 ) | ( n11156 & n11157 ) ;
  assign n11159 = n6796 & n10263 ;
  assign n11160 = x11 & n11159 ;
  assign n11161 = n6567 & n10265 ;
  assign n11162 = n6570 | n11161 ;
  assign n11163 = ( n10261 & n11161 ) | ( n10261 & n11162 ) | ( n11161 & n11162 ) ;
  assign n11164 = n6571 | n11163 ;
  assign n11165 = ( n11049 & n11163 ) | ( n11049 & n11164 ) | ( n11163 & n11164 ) ;
  assign n11166 = x11 & ~n11165 ;
  assign n11167 = ( ~x11 & n11159 ) | ( ~x11 & n11165 ) | ( n11159 & n11165 ) ;
  assign n11168 = ( ~n11160 & n11166 ) | ( ~n11160 & n11167 ) | ( n11166 & n11167 ) ;
  assign n11169 = n5584 & n10273 ;
  assign n11170 = x17 & n11169 ;
  assign n11171 = n5413 & n10275 ;
  assign n11172 = n5417 | n11171 ;
  assign n11173 = ( ~n10297 & n11171 ) | ( ~n10297 & n11172 ) | ( n11171 & n11172 ) ;
  assign n11174 = n5418 | n11173 ;
  assign n11175 = ( ~n10617 & n11173 ) | ( ~n10617 & n11174 ) | ( n11173 & n11174 ) ;
  assign n11176 = x17 & ~n11175 ;
  assign n11177 = ( ~x17 & n11169 ) | ( ~x17 & n11175 ) | ( n11169 & n11175 ) ;
  assign n11178 = ( ~n11170 & n11176 ) | ( ~n11170 & n11177 ) | ( n11176 & n11177 ) ;
  assign n11179 = n4879 & ~n10516 ;
  assign n11180 = x20 & n11179 ;
  assign n11181 = n4874 & ~n10279 ;
  assign n11182 = n4878 | n11181 ;
  assign n11183 = ( n10277 & n11181 ) | ( n10277 & n11182 ) | ( n11181 & n11182 ) ;
  assign n11184 = n5232 & n10291 ;
  assign n11185 = n11183 | n11184 ;
  assign n11186 = x20 & ~n11185 ;
  assign n11187 = ( ~x20 & n11179 ) | ( ~x20 & n11185 ) | ( n11179 & n11185 ) ;
  assign n11188 = ( ~n11180 & n11186 ) | ( ~n11180 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = x23 & n11119 ;
  assign n11190 = n4591 & n10464 ;
  assign n11191 = n4649 & n10281 ;
  assign n11192 = n4637 & ~n10283 ;
  assign n11193 = n4584 & ~n10285 ;
  assign n11194 = n11192 | n11193 ;
  assign n11195 = n11191 | n11194 ;
  assign n11196 = n11190 | n11195 ;
  assign n11197 = n11189 & ~n11196 ;
  assign n11198 = ~n11189 & n11196 ;
  assign n11199 = n11197 | n11198 ;
  assign n11200 = ( ~n11124 & n11188 ) | ( ~n11124 & n11199 ) | ( n11188 & n11199 ) ;
  assign n11201 = ( n11124 & n11188 ) | ( n11124 & n11199 ) | ( n11188 & n11199 ) ;
  assign n11202 = ( n11124 & n11200 ) | ( n11124 & ~n11201 ) | ( n11200 & ~n11201 ) ;
  assign n11203 = ( ~n11127 & n11178 ) | ( ~n11127 & n11202 ) | ( n11178 & n11202 ) ;
  assign n11204 = ( n11127 & n11178 ) | ( n11127 & n11202 ) | ( n11178 & n11202 ) ;
  assign n11205 = ( n11127 & n11203 ) | ( n11127 & ~n11204 ) | ( n11203 & ~n11204 ) ;
  assign n11206 = n5915 & ~n10787 ;
  assign n11207 = x14 & n11206 ;
  assign n11208 = n5909 & n10271 ;
  assign n11209 = n5914 | n11208 ;
  assign n11210 = ( n10267 & n11208 ) | ( n10267 & n11209 ) | ( n11208 & n11209 ) ;
  assign n11211 = n6332 & ~n10269 ;
  assign n11212 = n11210 | n11211 ;
  assign n11213 = x14 & ~n11212 ;
  assign n11214 = ( ~x14 & n11206 ) | ( ~x14 & n11212 ) | ( n11206 & n11212 ) ;
  assign n11215 = ( ~n11207 & n11213 ) | ( ~n11207 & n11214 ) | ( n11213 & n11214 ) ;
  assign n11216 = ( ~n11140 & n11205 ) | ( ~n11140 & n11215 ) | ( n11205 & n11215 ) ;
  assign n11217 = ( n11140 & n11205 ) | ( n11140 & n11215 ) | ( n11205 & n11215 ) ;
  assign n11218 = ( n11140 & n11216 ) | ( n11140 & ~n11217 ) | ( n11216 & ~n11217 ) ;
  assign n11219 = ( n11143 & n11168 ) | ( n11143 & n11218 ) | ( n11168 & n11218 ) ;
  assign n11220 = ( ~n11143 & n11168 ) | ( ~n11143 & n11218 ) | ( n11168 & n11218 ) ;
  assign n11221 = ( n11143 & ~n11219 ) | ( n11143 & n11220 ) | ( ~n11219 & n11220 ) ;
  assign n11222 = ( n11145 & n11158 ) | ( n11145 & n11221 ) | ( n11158 & n11221 ) ;
  assign n11223 = n6571 & n10859 ;
  assign n11224 = x11 & n11223 ;
  assign n11225 = n6567 & n10263 ;
  assign n11226 = n6570 | n11225 ;
  assign n11227 = ( n10259 & n11225 ) | ( n10259 & n11226 ) | ( n11225 & n11226 ) ;
  assign n11228 = n6796 & n10261 ;
  assign n11229 = n11227 | n11228 ;
  assign n11230 = x11 & ~n11229 ;
  assign n11231 = ( ~x11 & n11223 ) | ( ~x11 & n11229 ) | ( n11223 & n11229 ) ;
  assign n11232 = ( ~n11224 & n11230 ) | ( ~n11224 & n11231 ) | ( n11230 & n11231 ) ;
  assign n11233 = n6332 & n10267 ;
  assign n11234 = x14 & n11233 ;
  assign n11235 = n5909 & ~n10269 ;
  assign n11236 = n5914 | n11235 ;
  assign n11237 = ( n10265 & n11235 ) | ( n10265 & n11236 ) | ( n11235 & n11236 ) ;
  assign n11238 = n5915 | n11237 ;
  assign n11239 = ( n10804 & n11237 ) | ( n10804 & n11238 ) | ( n11237 & n11238 ) ;
  assign n11240 = x14 & ~n11239 ;
  assign n11241 = ( ~x14 & n11233 ) | ( ~x14 & n11239 ) | ( n11233 & n11239 ) ;
  assign n11242 = ( ~n11234 & n11240 ) | ( ~n11234 & n11241 ) | ( n11240 & n11241 ) ;
  assign n11243 = n5584 & ~n10297 ;
  assign n11244 = x17 & n11243 ;
  assign n11245 = n5413 & n10273 ;
  assign n11246 = n5417 | n11245 ;
  assign n11247 = ( n10271 & n11245 ) | ( n10271 & n11246 ) | ( n11245 & n11246 ) ;
  assign n11248 = n5418 | n11247 ;
  assign n11249 = ( ~n10656 & n11247 ) | ( ~n10656 & n11248 ) | ( n11247 & n11248 ) ;
  assign n11250 = x17 & ~n11249 ;
  assign n11251 = ( ~x17 & n11243 ) | ( ~x17 & n11249 ) | ( n11243 & n11249 ) ;
  assign n11252 = ( ~n11244 & n11250 ) | ( ~n11244 & n11251 ) | ( n11250 & n11251 ) ;
  assign n11253 = n5232 & n10277 ;
  assign n11254 = x20 & n11253 ;
  assign n11255 = n4874 & n10291 ;
  assign n11256 = n4878 | n11255 ;
  assign n11257 = ( n10275 & n11255 ) | ( n10275 & n11256 ) | ( n11255 & n11256 ) ;
  assign n11258 = n4879 | n11257 ;
  assign n11259 = ( n10563 & n11257 ) | ( n10563 & n11258 ) | ( n11257 & n11258 ) ;
  assign n11260 = x20 & ~n11259 ;
  assign n11261 = ( ~x20 & n11253 ) | ( ~x20 & n11259 ) | ( n11253 & n11259 ) ;
  assign n11262 = ( ~n11254 & n11260 ) | ( ~n11254 & n11261 ) | ( n11260 & n11261 ) ;
  assign n11263 = n4591 & n10487 ;
  assign n11264 = n4649 & ~n10279 ;
  assign n11265 = n4637 & n10281 ;
  assign n11266 = n4584 & ~n10283 ;
  assign n11267 = n11265 | n11266 ;
  assign n11268 = n11264 | n11267 ;
  assign n11269 = n11263 | n11268 ;
  assign n11270 = x23 & ~n11119 ;
  assign n11271 = ~n11196 & n11270 ;
  assign n11272 = n53 & ~n10285 ;
  assign n11273 = n11271 | n11272 ;
  assign n11274 = n4202 & ~n10285 ;
  assign n11275 = n68 & ~n10285 ;
  assign n11276 = ( n11271 & n11274 ) | ( n11271 & n11275 ) | ( n11274 & n11275 ) ;
  assign n11277 = ( x23 & ~n11273 ) | ( x23 & n11276 ) | ( ~n11273 & n11276 ) ;
  assign n11278 = ~n11269 & n11277 ;
  assign n11279 = n11269 & ~n11277 ;
  assign n11280 = n11278 | n11279 ;
  assign n11281 = ( ~n11201 & n11262 ) | ( ~n11201 & n11280 ) | ( n11262 & n11280 ) ;
  assign n11282 = ( n11201 & n11262 ) | ( n11201 & n11280 ) | ( n11262 & n11280 ) ;
  assign n11283 = ( n11201 & n11281 ) | ( n11201 & ~n11282 ) | ( n11281 & ~n11282 ) ;
  assign n11284 = ( ~n11204 & n11252 ) | ( ~n11204 & n11283 ) | ( n11252 & n11283 ) ;
  assign n11285 = ( n11204 & n11252 ) | ( n11204 & n11283 ) | ( n11252 & n11283 ) ;
  assign n11286 = ( n11204 & n11284 ) | ( n11204 & ~n11285 ) | ( n11284 & ~n11285 ) ;
  assign n11287 = ( ~n11217 & n11242 ) | ( ~n11217 & n11286 ) | ( n11242 & n11286 ) ;
  assign n11288 = ( n11217 & n11242 ) | ( n11217 & n11286 ) | ( n11242 & n11286 ) ;
  assign n11289 = ( n11217 & n11287 ) | ( n11217 & ~n11288 ) | ( n11287 & ~n11288 ) ;
  assign n11290 = ( ~n11219 & n11232 ) | ( ~n11219 & n11289 ) | ( n11232 & n11289 ) ;
  assign n11291 = ( n11219 & n11232 ) | ( n11219 & n11289 ) | ( n11232 & n11289 ) ;
  assign n11292 = ( n11219 & n11290 ) | ( n11219 & ~n11291 ) | ( n11290 & ~n11291 ) ;
  assign n11293 = n7644 & n10255 ;
  assign n11294 = x8 & n11293 ;
  assign n11295 = n10253 & ~n10351 ;
  assign n11296 = ( n10253 & ~n10307 ) | ( n10253 & n10351 ) | ( ~n10307 & n10351 ) ;
  assign n11297 = ( ~n10308 & n11295 ) | ( ~n10308 & n11296 ) | ( n11295 & n11296 ) ;
  assign n11298 = n7341 & n10257 ;
  assign n11299 = n7345 | n11298 ;
  assign n11300 = ( ~n10253 & n11298 ) | ( ~n10253 & n11299 ) | ( n11298 & n11299 ) ;
  assign n11301 = n7346 | n11300 ;
  assign n11302 = ( ~n11297 & n11300 ) | ( ~n11297 & n11301 ) | ( n11300 & n11301 ) ;
  assign n11303 = x8 & ~n11302 ;
  assign n11304 = ( ~x8 & n11293 ) | ( ~x8 & n11302 ) | ( n11293 & n11302 ) ;
  assign n11305 = ( ~n11294 & n11303 ) | ( ~n11294 & n11304 ) | ( n11303 & n11304 ) ;
  assign n11306 = ( n11222 & n11292 ) | ( n11222 & n11305 ) | ( n11292 & n11305 ) ;
  assign n11307 = n10251 & n10352 ;
  assign n11308 = ( ~n10251 & n10308 ) | ( ~n10251 & n10352 ) | ( n10308 & n10352 ) ;
  assign n11309 = ( n10309 & ~n11307 ) | ( n10309 & n11308 ) | ( ~n11307 & n11308 ) ;
  assign n11310 = n7346 & ~n11309 ;
  assign n11311 = x8 & n11310 ;
  assign n11312 = n7341 & n10255 ;
  assign n11313 = n7345 | n11312 ;
  assign n11314 = ( n10251 & n11312 ) | ( n10251 & n11313 ) | ( n11312 & n11313 ) ;
  assign n11315 = n7644 & ~n10253 ;
  assign n11316 = n11314 | n11315 ;
  assign n11317 = x8 & ~n11316 ;
  assign n11318 = ( ~x8 & n11310 ) | ( ~x8 & n11316 ) | ( n11310 & n11316 ) ;
  assign n11319 = ( ~n11311 & n11317 ) | ( ~n11311 & n11318 ) | ( n11317 & n11318 ) ;
  assign n11320 = n6796 & n10259 ;
  assign n11321 = x11 & n11320 ;
  assign n11322 = n6567 & n10261 ;
  assign n11323 = n6570 | n11322 ;
  assign n11324 = ( n10257 & n11322 ) | ( n10257 & n11323 ) | ( n11322 & n11323 ) ;
  assign n11325 = n6571 | n11324 ;
  assign n11326 = ( n11065 & n11324 ) | ( n11065 & n11325 ) | ( n11324 & n11325 ) ;
  assign n11327 = x11 & ~n11326 ;
  assign n11328 = ( ~x11 & n11320 ) | ( ~x11 & n11326 ) | ( n11320 & n11326 ) ;
  assign n11329 = ( ~n11321 & n11327 ) | ( ~n11321 & n11328 ) | ( n11327 & n11328 ) ;
  assign n11330 = n6332 & n10265 ;
  assign n11331 = x14 & n11330 ;
  assign n11332 = n5909 & n10267 ;
  assign n11333 = n5914 | n11332 ;
  assign n11334 = ( n10263 & n11332 ) | ( n10263 & n11333 ) | ( n11332 & n11333 ) ;
  assign n11335 = n5915 | n11334 ;
  assign n11336 = ( n10874 & n11334 ) | ( n10874 & n11335 ) | ( n11334 & n11335 ) ;
  assign n11337 = x14 & ~n11336 ;
  assign n11338 = ( ~x14 & n11330 ) | ( ~x14 & n11336 ) | ( n11330 & n11336 ) ;
  assign n11339 = ( ~n11331 & n11337 ) | ( ~n11331 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11340 = n5584 & n10271 ;
  assign n11341 = x17 & n11340 ;
  assign n11342 = n5413 & ~n10297 ;
  assign n11343 = n5417 | n11342 ;
  assign n11344 = ( ~n10269 & n11342 ) | ( ~n10269 & n11343 ) | ( n11342 & n11343 ) ;
  assign n11345 = n5418 | n11344 ;
  assign n11346 = ( ~n10698 & n11344 ) | ( ~n10698 & n11345 ) | ( n11344 & n11345 ) ;
  assign n11347 = x17 & ~n11346 ;
  assign n11348 = ( ~x17 & n11340 ) | ( ~x17 & n11346 ) | ( n11340 & n11346 ) ;
  assign n11349 = ( ~n11341 & n11347 ) | ( ~n11341 & n11348 ) | ( n11347 & n11348 ) ;
  assign n11350 = n5232 & n10275 ;
  assign n11351 = x20 & n11350 ;
  assign n11352 = n4874 & n10277 ;
  assign n11353 = n4878 | n11352 ;
  assign n11354 = ( n10273 & n11352 ) | ( n10273 & n11353 ) | ( n11352 & n11353 ) ;
  assign n11355 = n4879 | n11354 ;
  assign n11356 = ( n10577 & n11354 ) | ( n10577 & n11355 ) | ( n11354 & n11355 ) ;
  assign n11357 = x20 & ~n11356 ;
  assign n11358 = ( ~x20 & n11350 ) | ( ~x20 & n11356 ) | ( n11350 & n11356 ) ;
  assign n11359 = ( ~n11351 & n11357 ) | ( ~n11351 & n11358 ) | ( n11357 & n11358 ) ;
  assign n11360 = n4649 & n10291 ;
  assign n11361 = x23 & n11360 ;
  assign n11362 = n4637 & ~n10279 ;
  assign n11363 = n4584 & n10281 ;
  assign n11364 = n11362 | n11363 ;
  assign n11365 = n4591 | n11364 ;
  assign n11366 = ( n10454 & n11364 ) | ( n10454 & n11365 ) | ( n11364 & n11365 ) ;
  assign n11367 = x23 & ~n11366 ;
  assign n11368 = ( ~x23 & n11360 ) | ( ~x23 & n11366 ) | ( n11360 & n11366 ) ;
  assign n11369 = ( ~n11361 & n11367 ) | ( ~n11361 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11370 = n11269 & n11275 ;
  assign n11371 = n11269 & ~n11275 ;
  assign n11372 = ( n11273 & n11370 ) | ( n11273 & ~n11371 ) | ( n11370 & ~n11371 ) ;
  assign n11373 = n4200 | n4203 ;
  assign n11374 = ( n4200 & n10283 ) | ( n4200 & n11373 ) | ( n10283 & n11373 ) ;
  assign n11375 = ~n10285 & n11374 ;
  assign n11376 = ( n4202 & n4215 ) | ( n4202 & n10285 ) | ( n4215 & n10285 ) ;
  assign n11377 = ~n10283 & n11376 ;
  assign n11378 = n11375 | n11377 ;
  assign n11379 = n11274 | n11378 ;
  assign n11380 = ( x26 & n11274 ) | ( x26 & ~n11378 ) | ( n11274 & ~n11378 ) ;
  assign n11381 = x26 & ~n11378 ;
  assign n11382 = ( n11379 & ~n11380 ) | ( n11379 & n11381 ) | ( ~n11380 & n11381 ) ;
  assign n11383 = ( ~n11369 & n11372 ) | ( ~n11369 & n11382 ) | ( n11372 & n11382 ) ;
  assign n11384 = ( n11369 & n11372 ) | ( n11369 & n11382 ) | ( n11372 & n11382 ) ;
  assign n11385 = ( n11369 & n11383 ) | ( n11369 & ~n11384 ) | ( n11383 & ~n11384 ) ;
  assign n11386 = ( ~n11282 & n11359 ) | ( ~n11282 & n11385 ) | ( n11359 & n11385 ) ;
  assign n11387 = ( n11282 & n11359 ) | ( n11282 & n11385 ) | ( n11359 & n11385 ) ;
  assign n11388 = ( n11282 & n11386 ) | ( n11282 & ~n11387 ) | ( n11386 & ~n11387 ) ;
  assign n11389 = ( ~n11285 & n11349 ) | ( ~n11285 & n11388 ) | ( n11349 & n11388 ) ;
  assign n11390 = ( n11285 & n11349 ) | ( n11285 & n11388 ) | ( n11349 & n11388 ) ;
  assign n11391 = ( n11285 & n11389 ) | ( n11285 & ~n11390 ) | ( n11389 & ~n11390 ) ;
  assign n11392 = ( n11288 & n11339 ) | ( n11288 & n11391 ) | ( n11339 & n11391 ) ;
  assign n11393 = ( ~n11288 & n11339 ) | ( ~n11288 & n11391 ) | ( n11339 & n11391 ) ;
  assign n11394 = ( n11288 & ~n11392 ) | ( n11288 & n11393 ) | ( ~n11392 & n11393 ) ;
  assign n11395 = ( ~n11291 & n11329 ) | ( ~n11291 & n11394 ) | ( n11329 & n11394 ) ;
  assign n11396 = ( n11291 & n11329 ) | ( n11291 & n11394 ) | ( n11329 & n11394 ) ;
  assign n11397 = ( n11291 & n11395 ) | ( n11291 & ~n11396 ) | ( n11395 & ~n11396 ) ;
  assign n11398 = ( n11306 & n11319 ) | ( n11306 & n11397 ) | ( n11319 & n11397 ) ;
  assign n11399 = n6796 & n10257 ;
  assign n11400 = x11 & n11399 ;
  assign n11401 = n6567 & n10259 ;
  assign n11402 = n6570 | n11401 ;
  assign n11403 = ( n10255 & n11401 ) | ( n10255 & n11402 ) | ( n11401 & n11402 ) ;
  assign n11404 = n6571 | n11403 ;
  assign n11405 = ( n11148 & n11403 ) | ( n11148 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11406 = x11 & ~n11405 ;
  assign n11407 = ( ~x11 & n11399 ) | ( ~x11 & n11405 ) | ( n11399 & n11405 ) ;
  assign n11408 = ( ~n11400 & n11406 ) | ( ~n11400 & n11407 ) | ( n11406 & n11407 ) ;
  assign n11409 = n6332 & n10263 ;
  assign n11410 = x14 & n11409 ;
  assign n11411 = n5909 & n10265 ;
  assign n11412 = n5914 | n11411 ;
  assign n11413 = ( n10261 & n11411 ) | ( n10261 & n11412 ) | ( n11411 & n11412 ) ;
  assign n11414 = n5915 | n11413 ;
  assign n11415 = ( n11049 & n11413 ) | ( n11049 & n11414 ) | ( n11413 & n11414 ) ;
  assign n11416 = x14 & ~n11415 ;
  assign n11417 = ( ~x14 & n11409 ) | ( ~x14 & n11415 ) | ( n11409 & n11415 ) ;
  assign n11418 = ( ~n11410 & n11416 ) | ( ~n11410 & n11417 ) | ( n11416 & n11417 ) ;
  assign n11419 = n5584 & ~n10269 ;
  assign n11420 = x17 & n11419 ;
  assign n11421 = n5413 & n10271 ;
  assign n11422 = n5417 | n11421 ;
  assign n11423 = ( n10267 & n11421 ) | ( n10267 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11424 = n5418 | n11423 ;
  assign n11425 = ( ~n10787 & n11423 ) | ( ~n10787 & n11424 ) | ( n11423 & n11424 ) ;
  assign n11426 = x17 & ~n11425 ;
  assign n11427 = ( ~x17 & n11419 ) | ( ~x17 & n11425 ) | ( n11419 & n11425 ) ;
  assign n11428 = ( ~n11420 & n11426 ) | ( ~n11420 & n11427 ) | ( n11426 & n11427 ) ;
  assign n11429 = n5232 & n10273 ;
  assign n11430 = x20 & n11429 ;
  assign n11431 = n4874 & n10275 ;
  assign n11432 = n4878 | n11431 ;
  assign n11433 = ( ~n10297 & n11431 ) | ( ~n10297 & n11432 ) | ( n11431 & n11432 ) ;
  assign n11434 = n4879 | n11433 ;
  assign n11435 = ( ~n10617 & n11433 ) | ( ~n10617 & n11434 ) | ( n11433 & n11434 ) ;
  assign n11436 = x20 & ~n11435 ;
  assign n11437 = ( ~x20 & n11429 ) | ( ~x20 & n11435 ) | ( n11429 & n11435 ) ;
  assign n11438 = ( ~n11430 & n11436 ) | ( ~n11430 & n11437 ) | ( n11436 & n11437 ) ;
  assign n11439 = n4637 & n10291 ;
  assign n11440 = x23 & n11439 ;
  assign n11441 = n4584 & ~n10279 ;
  assign n11442 = n4649 | n11441 ;
  assign n11443 = ( n10277 & n11441 ) | ( n10277 & n11442 ) | ( n11441 & n11442 ) ;
  assign n11444 = n4591 | n11443 ;
  assign n11445 = ( ~n10516 & n11443 ) | ( ~n10516 & n11444 ) | ( n11443 & n11444 ) ;
  assign n11446 = x23 & ~n11445 ;
  assign n11447 = ( ~x23 & n11439 ) | ( ~x23 & n11445 ) | ( n11439 & n11445 ) ;
  assign n11448 = ( ~n11440 & n11446 ) | ( ~n11440 & n11447 ) | ( n11446 & n11447 ) ;
  assign n11449 = n4203 & n10464 ;
  assign n11450 = n4215 & n10281 ;
  assign n11451 = n4200 & ~n10283 ;
  assign n11452 = n2083 & ~n10285 ;
  assign n11453 = n11451 | n11452 ;
  assign n11454 = n11450 | n11453 ;
  assign n11455 = n11449 | n11454 ;
  assign n11456 = x26 & ~n11455 ;
  assign n11457 = ( x26 & n11379 ) | ( x26 & ~n11455 ) | ( n11379 & ~n11455 ) ;
  assign n11458 = ~n11379 & n11456 ;
  assign n11459 = ( x26 & n11455 ) | ( x26 & ~n11458 ) | ( n11455 & ~n11458 ) ;
  assign n11460 = ( n11456 & ~n11457 ) | ( n11456 & n11459 ) | ( ~n11457 & n11459 ) ;
  assign n11461 = ( n11384 & n11448 ) | ( n11384 & n11460 ) | ( n11448 & n11460 ) ;
  assign n11462 = ( ~n11384 & n11448 ) | ( ~n11384 & n11460 ) | ( n11448 & n11460 ) ;
  assign n11463 = ( n11384 & ~n11461 ) | ( n11384 & n11462 ) | ( ~n11461 & n11462 ) ;
  assign n11464 = ( ~n11387 & n11438 ) | ( ~n11387 & n11463 ) | ( n11438 & n11463 ) ;
  assign n11465 = ( n11387 & n11438 ) | ( n11387 & n11463 ) | ( n11438 & n11463 ) ;
  assign n11466 = ( n11387 & n11464 ) | ( n11387 & ~n11465 ) | ( n11464 & ~n11465 ) ;
  assign n11467 = ( ~n11390 & n11428 ) | ( ~n11390 & n11466 ) | ( n11428 & n11466 ) ;
  assign n11468 = ( n11390 & n11428 ) | ( n11390 & n11466 ) | ( n11428 & n11466 ) ;
  assign n11469 = ( n11390 & n11467 ) | ( n11390 & ~n11468 ) | ( n11467 & ~n11468 ) ;
  assign n11470 = ( ~n11392 & n11418 ) | ( ~n11392 & n11469 ) | ( n11418 & n11469 ) ;
  assign n11471 = ( n11392 & n11418 ) | ( n11392 & n11469 ) | ( n11418 & n11469 ) ;
  assign n11472 = ( n11392 & n11470 ) | ( n11392 & ~n11471 ) | ( n11470 & ~n11471 ) ;
  assign n11473 = ( ~n11396 & n11408 ) | ( ~n11396 & n11472 ) | ( n11408 & n11472 ) ;
  assign n11474 = ( n11396 & n11408 ) | ( n11396 & n11472 ) | ( n11408 & n11472 ) ;
  assign n11475 = ( n11396 & n11473 ) | ( n11396 & ~n11474 ) | ( n11473 & ~n11474 ) ;
  assign n11476 = ( n10449 & n11398 ) | ( n10449 & n11475 ) | ( n11398 & n11475 ) ;
  assign n11477 = n7345 & n10312 ;
  assign n11478 = n7644 & ~n10249 ;
  assign n11479 = n7341 & n10251 ;
  assign n11480 = n11478 | n11479 ;
  assign n11481 = n11477 | n11480 ;
  assign n11482 = x8 & n11481 ;
  assign n11483 = ( ~n10310 & n10312 ) | ( ~n10310 & n10354 ) | ( n10312 & n10354 ) ;
  assign n11484 = n10310 & ~n10312 ;
  assign n11485 = ( n10310 & n10312 ) | ( n10310 & n10354 ) | ( n10312 & n10354 ) ;
  assign n11486 = ( n11483 & n11484 ) | ( n11483 & ~n11485 ) | ( n11484 & ~n11485 ) ;
  assign n11487 = n7346 & ~n11486 ;
  assign n11488 = x8 & ~n11487 ;
  assign n11489 = ( ~x8 & n11481 ) | ( ~x8 & n11487 ) | ( n11481 & n11487 ) ;
  assign n11490 = ( ~n11482 & n11488 ) | ( ~n11482 & n11489 ) | ( n11488 & n11489 ) ;
  assign n11491 = n6571 & ~n11297 ;
  assign n11492 = x11 & n11491 ;
  assign n11493 = n6567 & n10257 ;
  assign n11494 = n6570 | n11493 ;
  assign n11495 = ( ~n10253 & n11493 ) | ( ~n10253 & n11494 ) | ( n11493 & n11494 ) ;
  assign n11496 = n6796 & n10255 ;
  assign n11497 = n11495 | n11496 ;
  assign n11498 = x11 & ~n11497 ;
  assign n11499 = ( ~x11 & n11491 ) | ( ~x11 & n11497 ) | ( n11491 & n11497 ) ;
  assign n11500 = ( ~n11492 & n11498 ) | ( ~n11492 & n11499 ) | ( n11498 & n11499 ) ;
  assign n11501 = n5584 & n10267 ;
  assign n11502 = x17 & n11501 ;
  assign n11503 = n5413 & ~n10269 ;
  assign n11504 = n5417 | n11503 ;
  assign n11505 = ( n10265 & n11503 ) | ( n10265 & n11504 ) | ( n11503 & n11504 ) ;
  assign n11506 = n5418 | n11505 ;
  assign n11507 = ( n10804 & n11505 ) | ( n10804 & n11506 ) | ( n11505 & n11506 ) ;
  assign n11508 = x17 & ~n11507 ;
  assign n11509 = ( ~x17 & n11501 ) | ( ~x17 & n11507 ) | ( n11501 & n11507 ) ;
  assign n11510 = ( ~n11502 & n11508 ) | ( ~n11502 & n11509 ) | ( n11508 & n11509 ) ;
  assign n11511 = n5232 & ~n10297 ;
  assign n11512 = x20 & n11511 ;
  assign n11513 = n4874 & n10273 ;
  assign n11514 = n4878 | n11513 ;
  assign n11515 = ( n10271 & n11513 ) | ( n10271 & n11514 ) | ( n11513 & n11514 ) ;
  assign n11516 = n4879 | n11515 ;
  assign n11517 = ( ~n10656 & n11515 ) | ( ~n10656 & n11516 ) | ( n11515 & n11516 ) ;
  assign n11518 = x20 & ~n11517 ;
  assign n11519 = ( ~x20 & n11511 ) | ( ~x20 & n11517 ) | ( n11511 & n11517 ) ;
  assign n11520 = ( ~n11512 & n11518 ) | ( ~n11512 & n11519 ) | ( n11518 & n11519 ) ;
  assign n11521 = n4637 & n10277 ;
  assign n11522 = x23 & n11521 ;
  assign n11523 = n4584 & n10291 ;
  assign n11524 = n4649 | n11523 ;
  assign n11525 = ( n10275 & n11523 ) | ( n10275 & n11524 ) | ( n11523 & n11524 ) ;
  assign n11526 = n4591 | n11525 ;
  assign n11527 = ( n10563 & n11525 ) | ( n10563 & n11526 ) | ( n11525 & n11526 ) ;
  assign n11528 = x23 & ~n11527 ;
  assign n11529 = ( ~x23 & n11521 ) | ( ~x23 & n11527 ) | ( n11521 & n11527 ) ;
  assign n11530 = ( ~n11522 & n11528 ) | ( ~n11522 & n11529 ) | ( n11528 & n11529 ) ;
  assign n11531 = n4203 & n10487 ;
  assign n11532 = n4215 & ~n10279 ;
  assign n11533 = n4200 & n10281 ;
  assign n11534 = n2083 & ~n10283 ;
  assign n11535 = n11533 | n11534 ;
  assign n11536 = n11532 | n11535 ;
  assign n11537 = n11531 | n11536 ;
  assign n11538 = x27 | n10285 ;
  assign n11539 = ~x26 & n10285 ;
  assign n11540 = n11538 & ~n11539 ;
  assign n11541 = ( n11537 & ~n11538 ) | ( n11537 & n11540 ) | ( ~n11538 & n11540 ) ;
  assign n11542 = ( n11458 & n11538 ) | ( n11458 & n11541 ) | ( n11538 & n11541 ) ;
  assign n11543 = ( n11458 & n11540 ) | ( n11458 & ~n11541 ) | ( n11540 & ~n11541 ) ;
  assign n11544 = ( n11537 & ~n11542 ) | ( n11537 & n11543 ) | ( ~n11542 & n11543 ) ;
  assign n11545 = ( ~n11461 & n11530 ) | ( ~n11461 & n11544 ) | ( n11530 & n11544 ) ;
  assign n11546 = ( n11461 & n11530 ) | ( n11461 & n11544 ) | ( n11530 & n11544 ) ;
  assign n11547 = ( n11461 & n11545 ) | ( n11461 & ~n11546 ) | ( n11545 & ~n11546 ) ;
  assign n11548 = ( ~n11465 & n11520 ) | ( ~n11465 & n11547 ) | ( n11520 & n11547 ) ;
  assign n11549 = ( n11465 & n11520 ) | ( n11465 & n11547 ) | ( n11520 & n11547 ) ;
  assign n11550 = ( n11465 & n11548 ) | ( n11465 & ~n11549 ) | ( n11548 & ~n11549 ) ;
  assign n11551 = ( ~n11468 & n11510 ) | ( ~n11468 & n11550 ) | ( n11510 & n11550 ) ;
  assign n11552 = ( n11468 & n11510 ) | ( n11468 & n11550 ) | ( n11510 & n11550 ) ;
  assign n11553 = ( n11468 & n11551 ) | ( n11468 & ~n11552 ) | ( n11551 & ~n11552 ) ;
  assign n11554 = n6332 & n10261 ;
  assign n11555 = x14 & n11554 ;
  assign n11556 = n5909 & n10263 ;
  assign n11557 = n5914 | n11556 ;
  assign n11558 = ( n10259 & n11556 ) | ( n10259 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11559 = n5915 | n11558 ;
  assign n11560 = ( n10859 & n11558 ) | ( n10859 & n11559 ) | ( n11558 & n11559 ) ;
  assign n11561 = x14 & ~n11560 ;
  assign n11562 = ( ~x14 & n11554 ) | ( ~x14 & n11560 ) | ( n11554 & n11560 ) ;
  assign n11563 = ( ~n11555 & n11561 ) | ( ~n11555 & n11562 ) | ( n11561 & n11562 ) ;
  assign n11564 = ( ~n11471 & n11553 ) | ( ~n11471 & n11563 ) | ( n11553 & n11563 ) ;
  assign n11565 = ( n11471 & n11553 ) | ( n11471 & n11563 ) | ( n11553 & n11563 ) ;
  assign n11566 = ( n11471 & n11564 ) | ( n11471 & ~n11565 ) | ( n11564 & ~n11565 ) ;
  assign n11567 = ( ~n11474 & n11500 ) | ( ~n11474 & n11566 ) | ( n11500 & n11566 ) ;
  assign n11568 = ( n11474 & n11500 ) | ( n11474 & n11566 ) | ( n11500 & n11566 ) ;
  assign n11569 = ( n11474 & n11567 ) | ( n11474 & ~n11568 ) | ( n11567 & ~n11568 ) ;
  assign n11570 = ( n11476 & n11490 ) | ( n11476 & n11569 ) | ( n11490 & n11569 ) ;
  assign n11571 = n6571 & ~n11309 ;
  assign n11572 = x11 & n11571 ;
  assign n11573 = n6567 & n10255 ;
  assign n11574 = n6570 | n11573 ;
  assign n11575 = ( n10251 & n11573 ) | ( n10251 & n11574 ) | ( n11573 & n11574 ) ;
  assign n11576 = n6796 & ~n10253 ;
  assign n11577 = n11575 | n11576 ;
  assign n11578 = x11 & ~n11577 ;
  assign n11579 = ( ~x11 & n11571 ) | ( ~x11 & n11577 ) | ( n11571 & n11577 ) ;
  assign n11580 = ( ~n11572 & n11578 ) | ( ~n11572 & n11579 ) | ( n11578 & n11579 ) ;
  assign n11581 = n6332 & n10259 ;
  assign n11582 = x14 & n11581 ;
  assign n11583 = n5909 & n10261 ;
  assign n11584 = n5914 | n11583 ;
  assign n11585 = ( n10257 & n11583 ) | ( n10257 & n11584 ) | ( n11583 & n11584 ) ;
  assign n11586 = n5915 | n11585 ;
  assign n11587 = ( n11065 & n11585 ) | ( n11065 & n11586 ) | ( n11585 & n11586 ) ;
  assign n11588 = x14 & ~n11587 ;
  assign n11589 = ( ~x14 & n11581 ) | ( ~x14 & n11587 ) | ( n11581 & n11587 ) ;
  assign n11590 = ( ~n11582 & n11588 ) | ( ~n11582 & n11589 ) | ( n11588 & n11589 ) ;
  assign n11591 = n5232 & n10271 ;
  assign n11592 = n4879 | n11591 ;
  assign n11593 = ( ~n10698 & n11591 ) | ( ~n10698 & n11592 ) | ( n11591 & n11592 ) ;
  assign n11594 = n4874 & ~n10297 ;
  assign n11595 = ( ~x20 & n11593 ) | ( ~x20 & n11594 ) | ( n11593 & n11594 ) ;
  assign n11596 = n4878 & ~n10269 ;
  assign n11597 = x20 & ~n11594 ;
  assign n11598 = n11596 | n11597 ;
  assign n11599 = ( n11593 & n11596 ) | ( n11593 & n11597 ) | ( n11596 & n11597 ) ;
  assign n11600 = ( n11595 & n11598 ) | ( n11595 & ~n11599 ) | ( n11598 & ~n11599 ) ;
  assign n11601 = n4637 & n10275 ;
  assign n11602 = x23 & n11601 ;
  assign n11603 = n4584 & n10277 ;
  assign n11604 = n4649 | n11603 ;
  assign n11605 = ( n10273 & n11603 ) | ( n10273 & n11604 ) | ( n11603 & n11604 ) ;
  assign n11606 = n4591 | n11605 ;
  assign n11607 = ( n10577 & n11605 ) | ( n10577 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11608 = x23 & ~n11607 ;
  assign n11609 = ( ~x23 & n11601 ) | ( ~x23 & n11607 ) | ( n11601 & n11607 ) ;
  assign n11610 = ( ~n11602 & n11608 ) | ( ~n11602 & n11609 ) | ( n11608 & n11609 ) ;
  assign n11611 = n4215 & n10291 ;
  assign n11612 = x26 & n11611 ;
  assign n11613 = n4200 & ~n10279 ;
  assign n11614 = n2083 & n10281 ;
  assign n11615 = n11613 | n11614 ;
  assign n11616 = n4203 | n11615 ;
  assign n11617 = ( n10454 & n11615 ) | ( n10454 & n11616 ) | ( n11615 & n11616 ) ;
  assign n11618 = x26 & ~n11617 ;
  assign n11619 = ( ~x26 & n11611 ) | ( ~x26 & n11617 ) | ( n11611 & n11617 ) ;
  assign n11620 = ( ~n11612 & n11618 ) | ( ~n11612 & n11619 ) | ( n11618 & n11619 ) ;
  assign n11621 = n3499 & ~n10285 ;
  assign n11622 = n11537 & n11621 ;
  assign n11623 = n11537 & ~n11621 ;
  assign n11624 = ( x26 & n11458 ) | ( x26 & ~n11538 ) | ( n11458 & ~n11538 ) ;
  assign n11625 = ( n11622 & ~n11623 ) | ( n11622 & n11624 ) | ( ~n11623 & n11624 ) ;
  assign n11626 = ( n3500 & n4039 ) | ( n3500 & n10285 ) | ( n4039 & n10285 ) ;
  assign n11627 = ~n10283 & n11626 ;
  assign n11628 = ( n3501 & n6605 ) | ( n3501 & n10283 ) | ( n6605 & n10283 ) ;
  assign n11629 = ~n10285 & n11628 ;
  assign n11630 = n11627 | n11629 ;
  assign n11631 = n3500 & ~n10285 ;
  assign n11632 = n11630 | n11631 ;
  assign n11633 = ( x29 & ~n11630 ) | ( x29 & n11631 ) | ( ~n11630 & n11631 ) ;
  assign n11634 = x29 & ~n11630 ;
  assign n11635 = ( n11632 & ~n11633 ) | ( n11632 & n11634 ) | ( ~n11633 & n11634 ) ;
  assign n11636 = ( ~n11620 & n11625 ) | ( ~n11620 & n11635 ) | ( n11625 & n11635 ) ;
  assign n11637 = ( n11620 & n11625 ) | ( n11620 & n11635 ) | ( n11625 & n11635 ) ;
  assign n11638 = ( n11620 & n11636 ) | ( n11620 & ~n11637 ) | ( n11636 & ~n11637 ) ;
  assign n11639 = ( ~n11546 & n11610 ) | ( ~n11546 & n11638 ) | ( n11610 & n11638 ) ;
  assign n11640 = ( n11546 & n11610 ) | ( n11546 & n11638 ) | ( n11610 & n11638 ) ;
  assign n11641 = ( n11546 & n11639 ) | ( n11546 & ~n11640 ) | ( n11639 & ~n11640 ) ;
  assign n11642 = ( n11549 & n11600 ) | ( n11549 & n11641 ) | ( n11600 & n11641 ) ;
  assign n11643 = ( ~n11549 & n11600 ) | ( ~n11549 & n11641 ) | ( n11600 & n11641 ) ;
  assign n11644 = ( n11549 & ~n11642 ) | ( n11549 & n11643 ) | ( ~n11642 & n11643 ) ;
  assign n11645 = n5584 & n10265 ;
  assign n11646 = x17 & n11645 ;
  assign n11647 = n5413 & n10267 ;
  assign n11648 = n5417 | n11647 ;
  assign n11649 = ( n10263 & n11647 ) | ( n10263 & n11648 ) | ( n11647 & n11648 ) ;
  assign n11650 = n5418 | n11649 ;
  assign n11651 = ( n10874 & n11649 ) | ( n10874 & n11650 ) | ( n11649 & n11650 ) ;
  assign n11652 = x17 & ~n11651 ;
  assign n11653 = ( ~x17 & n11645 ) | ( ~x17 & n11651 ) | ( n11645 & n11651 ) ;
  assign n11654 = ( ~n11646 & n11652 ) | ( ~n11646 & n11653 ) | ( n11652 & n11653 ) ;
  assign n11655 = ( ~n11552 & n11644 ) | ( ~n11552 & n11654 ) | ( n11644 & n11654 ) ;
  assign n11656 = ( n11552 & n11644 ) | ( n11552 & n11654 ) | ( n11644 & n11654 ) ;
  assign n11657 = ( n11552 & n11655 ) | ( n11552 & ~n11656 ) | ( n11655 & ~n11656 ) ;
  assign n11658 = ( ~n11565 & n11590 ) | ( ~n11565 & n11657 ) | ( n11590 & n11657 ) ;
  assign n11659 = ( n11565 & n11590 ) | ( n11565 & n11657 ) | ( n11590 & n11657 ) ;
  assign n11660 = ( n11565 & n11658 ) | ( n11565 & ~n11659 ) | ( n11658 & ~n11659 ) ;
  assign n11661 = ( ~n11568 & n11580 ) | ( ~n11568 & n11660 ) | ( n11580 & n11660 ) ;
  assign n11662 = ( n11568 & n11580 ) | ( n11568 & n11660 ) | ( n11580 & n11660 ) ;
  assign n11663 = ( n11568 & n11661 ) | ( n11568 & ~n11662 ) | ( n11661 & ~n11662 ) ;
  assign n11664 = ( n10436 & n11570 ) | ( n10436 & n11663 ) | ( n11570 & n11663 ) ;
  assign n11665 = ( ~n10436 & n11570 ) | ( ~n10436 & n11663 ) | ( n11570 & n11663 ) ;
  assign n11666 = ( n10436 & ~n11664 ) | ( n10436 & n11665 ) | ( ~n11664 & n11665 ) ;
  assign n11667 = n40 & n10245 ;
  assign n11668 = n8721 & ~n10316 ;
  assign n11669 = n8340 & n10247 ;
  assign n11670 = n11668 | n11669 ;
  assign n11671 = n11667 | n11670 ;
  assign n11672 = x5 & n11671 ;
  assign n11673 = ( ~n10245 & n10317 ) | ( ~n10245 & n10357 ) | ( n10317 & n10357 ) ;
  assign n11674 = n10245 & ~n10317 ;
  assign n11675 = ( n10245 & n10317 ) | ( n10245 & n10357 ) | ( n10317 & n10357 ) ;
  assign n11676 = ( n11673 & n11674 ) | ( n11673 & ~n11675 ) | ( n11674 & ~n11675 ) ;
  assign n11677 = n8341 & ~n11676 ;
  assign n11678 = ( ~x5 & n11671 ) | ( ~x5 & n11677 ) | ( n11671 & n11677 ) ;
  assign n11679 = x5 & ~n11677 ;
  assign n11680 = ( ~n11672 & n11678 ) | ( ~n11672 & n11679 ) | ( n11678 & n11679 ) ;
  assign n11681 = ( ~n11476 & n11490 ) | ( ~n11476 & n11569 ) | ( n11490 & n11569 ) ;
  assign n11682 = ( n11476 & ~n11570 ) | ( n11476 & n11681 ) | ( ~n11570 & n11681 ) ;
  assign n11683 = n40 & ~n10316 ;
  assign n11684 = n8721 & n10247 ;
  assign n11685 = n8340 & n10312 ;
  assign n11686 = n11684 | n11685 ;
  assign n11687 = n11683 | n11686 ;
  assign n11688 = x5 & n11687 ;
  assign n11689 = n10314 & n10357 ;
  assign n11690 = ( ~n10247 & n10317 ) | ( ~n10247 & n10425 ) | ( n10317 & n10425 ) ;
  assign n11691 = ( n10316 & ~n11689 ) | ( n10316 & n11690 ) | ( ~n11689 & n11690 ) ;
  assign n11692 = n8341 & ~n11691 ;
  assign n11693 = ( ~x5 & n11687 ) | ( ~x5 & n11692 ) | ( n11687 & n11692 ) ;
  assign n11694 = x5 & ~n11692 ;
  assign n11695 = ( ~n11688 & n11693 ) | ( ~n11688 & n11694 ) | ( n11693 & n11694 ) ;
  assign n11696 = n40 & n10312 ;
  assign n11697 = x5 & n11696 ;
  assign n11698 = n8721 & ~n10249 ;
  assign n11699 = n8340 & n10251 ;
  assign n11700 = n11698 | n11699 ;
  assign n11701 = n8341 | n11700 ;
  assign n11702 = ( ~n11486 & n11700 ) | ( ~n11486 & n11701 ) | ( n11700 & n11701 ) ;
  assign n11703 = x5 & ~n11702 ;
  assign n11704 = ( ~x5 & n11696 ) | ( ~x5 & n11702 ) | ( n11696 & n11702 ) ;
  assign n11705 = ( ~n11697 & n11703 ) | ( ~n11697 & n11704 ) | ( n11703 & n11704 ) ;
  assign n11706 = ( ~n11222 & n11292 ) | ( ~n11222 & n11305 ) | ( n11292 & n11305 ) ;
  assign n11707 = ( n11222 & ~n11306 ) | ( n11222 & n11706 ) | ( ~n11306 & n11706 ) ;
  assign n11708 = n40 & ~n10249 ;
  assign n11709 = n8721 & n10251 ;
  assign n11710 = n8340 & ~n10253 ;
  assign n11711 = n11709 | n11710 ;
  assign n11712 = n11708 | n11711 ;
  assign n11713 = x5 & n11712 ;
  assign n11714 = n8341 & ~n10441 ;
  assign n11715 = ( ~x5 & n11712 ) | ( ~x5 & n11714 ) | ( n11712 & n11714 ) ;
  assign n11716 = x5 & ~n11714 ;
  assign n11717 = ( ~n11713 & n11715 ) | ( ~n11713 & n11716 ) | ( n11715 & n11716 ) ;
  assign n11718 = ( ~n11145 & n11158 ) | ( ~n11145 & n11221 ) | ( n11158 & n11221 ) ;
  assign n11719 = ( n11145 & ~n11222 ) | ( n11145 & n11718 ) | ( ~n11222 & n11718 ) ;
  assign n11720 = n40 & n10251 ;
  assign n11721 = n8721 & ~n10253 ;
  assign n11722 = n8340 & n10255 ;
  assign n11723 = n11721 | n11722 ;
  assign n11724 = n11720 | n11723 ;
  assign n11725 = x5 & n11724 ;
  assign n11726 = n8341 & ~n11309 ;
  assign n11727 = ( ~x5 & n11724 ) | ( ~x5 & n11726 ) | ( n11724 & n11726 ) ;
  assign n11728 = x5 & ~n11726 ;
  assign n11729 = ( ~n11725 & n11727 ) | ( ~n11725 & n11728 ) | ( n11727 & n11728 ) ;
  assign n11730 = n40 & ~n10253 ;
  assign n11731 = n8721 & n10255 ;
  assign n11732 = n8340 & n10257 ;
  assign n11733 = n11731 | n11732 ;
  assign n11734 = n11730 | n11733 ;
  assign n11735 = x5 & n11734 ;
  assign n11736 = n8341 & ~n11297 ;
  assign n11737 = ( ~x5 & n11734 ) | ( ~x5 & n11736 ) | ( n11734 & n11736 ) ;
  assign n11738 = x5 & ~n11736 ;
  assign n11739 = ( ~n11735 & n11737 ) | ( ~n11735 & n11738 ) | ( n11737 & n11738 ) ;
  assign n11740 = ( ~n10855 & n10869 ) | ( ~n10855 & n11060 ) | ( n10869 & n11060 ) ;
  assign n11741 = ( n10855 & ~n11061 ) | ( n10855 & n11740 ) | ( ~n11061 & n11740 ) ;
  assign n11742 = n40 & n10255 ;
  assign n11743 = n8721 & n10257 ;
  assign n11744 = n8340 & n10259 ;
  assign n11745 = n11743 | n11744 ;
  assign n11746 = n11742 | n11745 ;
  assign n11747 = x5 & n11746 ;
  assign n11748 = n8341 & n11148 ;
  assign n11749 = ( ~x5 & n11746 ) | ( ~x5 & n11748 ) | ( n11746 & n11748 ) ;
  assign n11750 = x5 & ~n11748 ;
  assign n11751 = ( ~n11747 & n11749 ) | ( ~n11747 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11752 = ( ~n11043 & n11045 ) | ( ~n11043 & n11059 ) | ( n11045 & n11059 ) ;
  assign n11753 = ( n11043 & ~n11060 ) | ( n11043 & n11752 ) | ( ~n11060 & n11752 ) ;
  assign n11754 = n40 & n10257 ;
  assign n11755 = n8721 & n10259 ;
  assign n11756 = n8340 & n10261 ;
  assign n11757 = n11755 | n11756 ;
  assign n11758 = n11754 | n11757 ;
  assign n11759 = x5 & n11758 ;
  assign n11760 = n8341 & n11065 ;
  assign n11761 = ( ~x5 & n11758 ) | ( ~x5 & n11760 ) | ( n11758 & n11760 ) ;
  assign n11762 = x5 & ~n11760 ;
  assign n11763 = ( ~n11759 & n11761 ) | ( ~n11759 & n11762 ) | ( n11761 & n11762 ) ;
  assign n11764 = ( ~n10871 & n10884 ) | ( ~n10871 & n11042 ) | ( n10884 & n11042 ) ;
  assign n11765 = ( n10871 & ~n11043 ) | ( n10871 & n11764 ) | ( ~n11043 & n11764 ) ;
  assign n11766 = n40 & n10259 ;
  assign n11767 = n8721 & n10261 ;
  assign n11768 = n8340 & n10263 ;
  assign n11769 = n11767 | n11768 ;
  assign n11770 = n11766 | n11769 ;
  assign n11771 = x5 & n11770 ;
  assign n11772 = n8341 & n10859 ;
  assign n11773 = ( ~x5 & n11770 ) | ( ~x5 & n11772 ) | ( n11770 & n11772 ) ;
  assign n11774 = x5 & ~n11772 ;
  assign n11775 = ( ~n11771 & n11773 ) | ( ~n11771 & n11774 ) | ( n11773 & n11774 ) ;
  assign n11776 = ( ~n11029 & n11031 ) | ( ~n11029 & n11041 ) | ( n11031 & n11041 ) ;
  assign n11777 = ( n11029 & ~n11042 ) | ( n11029 & n11776 ) | ( ~n11042 & n11776 ) ;
  assign n11778 = n40 & n10261 ;
  assign n11779 = n8721 & n10263 ;
  assign n11780 = n8340 & n10265 ;
  assign n11781 = n11779 | n11780 ;
  assign n11782 = n11778 | n11781 ;
  assign n11783 = x5 & n11782 ;
  assign n11784 = n8341 & n11049 ;
  assign n11785 = ( ~x5 & n11782 ) | ( ~x5 & n11784 ) | ( n11782 & n11784 ) ;
  assign n11786 = x5 & ~n11784 ;
  assign n11787 = ( ~n11783 & n11785 ) | ( ~n11783 & n11786 ) | ( n11785 & n11786 ) ;
  assign n11788 = ( ~n11016 & n11018 ) | ( ~n11016 & n11028 ) | ( n11018 & n11028 ) ;
  assign n11789 = ( n11016 & ~n11029 ) | ( n11016 & n11788 ) | ( ~n11029 & n11788 ) ;
  assign n11790 = n40 & n10291 ;
  assign n11791 = x5 & n11790 ;
  assign n11792 = n8721 & ~n10279 ;
  assign n11793 = n8340 & n10281 ;
  assign n11794 = n11792 | n11793 ;
  assign n11795 = n8341 | n11794 ;
  assign n11796 = ( n10454 & n11794 ) | ( n10454 & n11795 ) | ( n11794 & n11795 ) ;
  assign n11797 = x5 & ~n11796 ;
  assign n11798 = ( ~x5 & n11790 ) | ( ~x5 & n11796 ) | ( n11790 & n11796 ) ;
  assign n11799 = ( ~n11791 & n11797 ) | ( ~n11791 & n11798 ) | ( n11797 & n11798 ) ;
  assign n11800 = n10915 & ~n10917 ;
  assign n11801 = ( ~n10915 & n10918 ) | ( ~n10915 & n11800 ) | ( n10918 & n11800 ) ;
  assign n11802 = n8341 | n8721 ;
  assign n11803 = ( n8721 & n10283 ) | ( n8721 & n11802 ) | ( n10283 & n11802 ) ;
  assign n11804 = ~n10285 & n11803 ;
  assign n11805 = ( n36 & n40 ) | ( n36 & n10285 ) | ( n40 & n10285 ) ;
  assign n11806 = ~n10283 & n11805 ;
  assign n11807 = n11804 | n11806 ;
  assign n11808 = x5 & n36 ;
  assign n11809 = ~n10285 & n11808 ;
  assign n11810 = n11807 | n11809 ;
  assign n11811 = x5 & ~n11810 ;
  assign n11812 = n8341 & n10464 ;
  assign n11813 = n40 & n10281 ;
  assign n11814 = n8721 & ~n10283 ;
  assign n11815 = n8340 & ~n10285 ;
  assign n11816 = n11814 | n11815 ;
  assign n11817 = n11813 | n11816 ;
  assign n11818 = n11812 | n11817 ;
  assign n11819 = n11811 & ~n11818 ;
  assign n11820 = n10916 & ~n11819 ;
  assign n11821 = n8341 & n10487 ;
  assign n11822 = n40 & ~n10279 ;
  assign n11823 = n8721 & n10281 ;
  assign n11824 = n8340 & ~n10283 ;
  assign n11825 = n11823 | n11824 ;
  assign n11826 = n11822 | n11825 ;
  assign n11827 = n11821 | n11826 ;
  assign n11828 = x5 & ~n11819 ;
  assign n11829 = ( n10916 & n11827 ) | ( n10916 & ~n11828 ) | ( n11827 & ~n11828 ) ;
  assign n11830 = ( n10916 & ~n11827 ) | ( n10916 & n11828 ) | ( ~n11827 & n11828 ) ;
  assign n11831 = ( ~n11820 & n11829 ) | ( ~n11820 & n11830 ) | ( n11829 & n11830 ) ;
  assign n11832 = ( n10916 & n11820 ) | ( n10916 & ~n11827 ) | ( n11820 & ~n11827 ) ;
  assign n11833 = ( n11819 & ~n11831 ) | ( n11819 & n11832 ) | ( ~n11831 & n11832 ) ;
  assign n11834 = ( n11799 & n11801 ) | ( n11799 & n11833 ) | ( n11801 & n11833 ) ;
  assign n11835 = n40 & n10277 ;
  assign n11836 = n8721 & n10291 ;
  assign n11837 = n8340 & ~n10279 ;
  assign n11838 = n11836 | n11837 ;
  assign n11839 = n11835 | n11838 ;
  assign n11840 = x5 & n11839 ;
  assign n11841 = n8341 & ~n10516 ;
  assign n11842 = ( ~x5 & n11839 ) | ( ~x5 & n11841 ) | ( n11839 & n11841 ) ;
  assign n11843 = x5 & ~n11841 ;
  assign n11844 = ( ~n11840 & n11842 ) | ( ~n11840 & n11843 ) | ( n11842 & n11843 ) ;
  assign n11845 = ~x8 & n10926 ;
  assign n11846 = ( x8 & n10918 ) | ( x8 & n10926 ) | ( n10918 & n10926 ) ;
  assign n11847 = n10918 & n10926 ;
  assign n11848 = ( n11845 & n11846 ) | ( n11845 & ~n11847 ) | ( n11846 & ~n11847 ) ;
  assign n11849 = ( n11834 & n11844 ) | ( n11834 & n11848 ) | ( n11844 & n11848 ) ;
  assign n11850 = n40 & n10275 ;
  assign n11851 = n8721 & n10277 ;
  assign n11852 = n8340 & n10291 ;
  assign n11853 = n11851 | n11852 ;
  assign n11854 = n11850 | n11853 ;
  assign n11855 = x5 & n11854 ;
  assign n11856 = n8341 & n10563 ;
  assign n11857 = ( ~x5 & n11854 ) | ( ~x5 & n11856 ) | ( n11854 & n11856 ) ;
  assign n11858 = x5 & ~n11856 ;
  assign n11859 = ( ~n11855 & n11857 ) | ( ~n11855 & n11858 ) | ( n11857 & n11858 ) ;
  assign n11860 = ( n10930 & n11849 ) | ( n10930 & n11859 ) | ( n11849 & n11859 ) ;
  assign n11861 = n40 & n10273 ;
  assign n11862 = n8721 & n10275 ;
  assign n11863 = n8340 & n10277 ;
  assign n11864 = n11862 | n11863 ;
  assign n11865 = n11861 | n11864 ;
  assign n11866 = x5 & n11865 ;
  assign n11867 = n8341 & n10577 ;
  assign n11868 = ( ~x5 & n11865 ) | ( ~x5 & n11867 ) | ( n11865 & n11867 ) ;
  assign n11869 = x5 & ~n11867 ;
  assign n11870 = ( ~n11866 & n11868 ) | ( ~n11866 & n11869 ) | ( n11868 & n11869 ) ;
  assign n11871 = ( ~n10894 & n10898 ) | ( ~n10894 & n10931 ) | ( n10898 & n10931 ) ;
  assign n11872 = ( n10894 & ~n10932 ) | ( n10894 & n11871 ) | ( ~n10932 & n11871 ) ;
  assign n11873 = ( n11860 & n11870 ) | ( n11860 & n11872 ) | ( n11870 & n11872 ) ;
  assign n11874 = n40 & ~n10297 ;
  assign n11875 = n8721 & n10273 ;
  assign n11876 = n8340 & n10275 ;
  assign n11877 = n11875 | n11876 ;
  assign n11878 = n11874 | n11877 ;
  assign n11879 = x5 & n11878 ;
  assign n11880 = n8341 & ~n10617 ;
  assign n11881 = ( ~x5 & n11878 ) | ( ~x5 & n11880 ) | ( n11878 & n11880 ) ;
  assign n11882 = x5 & ~n11880 ;
  assign n11883 = ( ~n11879 & n11881 ) | ( ~n11879 & n11882 ) | ( n11881 & n11882 ) ;
  assign n11884 = ( ~n10932 & n10942 ) | ( ~n10932 & n10946 ) | ( n10942 & n10946 ) ;
  assign n11885 = ( n10932 & ~n10947 ) | ( n10932 & n11884 ) | ( ~n10947 & n11884 ) ;
  assign n11886 = ( n11873 & n11883 ) | ( n11873 & n11885 ) | ( n11883 & n11885 ) ;
  assign n11887 = n40 & n10271 ;
  assign n11888 = n8721 & ~n10297 ;
  assign n11889 = n8340 & n10273 ;
  assign n11890 = n11888 | n11889 ;
  assign n11891 = n11887 | n11890 ;
  assign n11892 = x5 & n11891 ;
  assign n11893 = n8341 & ~n10656 ;
  assign n11894 = ( ~x5 & n11891 ) | ( ~x5 & n11893 ) | ( n11891 & n11893 ) ;
  assign n11895 = x5 & ~n11893 ;
  assign n11896 = ( ~n11892 & n11894 ) | ( ~n11892 & n11895 ) | ( n11894 & n11895 ) ;
  assign n11897 = ( ~n10947 & n10957 ) | ( ~n10947 & n10963 ) | ( n10957 & n10963 ) ;
  assign n11898 = ( n10947 & ~n10964 ) | ( n10947 & n11897 ) | ( ~n10964 & n11897 ) ;
  assign n11899 = ( n11886 & n11896 ) | ( n11886 & n11898 ) | ( n11896 & n11898 ) ;
  assign n11900 = ( ~n10964 & n10974 ) | ( ~n10964 & n10976 ) | ( n10974 & n10976 ) ;
  assign n11901 = ( n10964 & ~n10977 ) | ( n10964 & n11900 ) | ( ~n10977 & n11900 ) ;
  assign n11902 = n40 & ~n10269 ;
  assign n11903 = n8721 & n10271 ;
  assign n11904 = n8340 & ~n10297 ;
  assign n11905 = n11903 | n11904 ;
  assign n11906 = n11902 | n11905 ;
  assign n11907 = x5 & n11906 ;
  assign n11908 = n8341 & ~n10698 ;
  assign n11909 = ( ~x5 & n11906 ) | ( ~x5 & n11908 ) | ( n11906 & n11908 ) ;
  assign n11910 = x5 & ~n11908 ;
  assign n11911 = ( ~n11907 & n11909 ) | ( ~n11907 & n11910 ) | ( n11909 & n11910 ) ;
  assign n11912 = ( n11899 & n11901 ) | ( n11899 & n11911 ) | ( n11901 & n11911 ) ;
  assign n11913 = n40 & n10267 ;
  assign n11914 = n8721 & ~n10269 ;
  assign n11915 = n8340 & n10271 ;
  assign n11916 = n11914 | n11915 ;
  assign n11917 = n11913 | n11916 ;
  assign n11918 = x5 & n11917 ;
  assign n11919 = n8341 & ~n10787 ;
  assign n11920 = ( ~x5 & n11917 ) | ( ~x5 & n11919 ) | ( n11917 & n11919 ) ;
  assign n11921 = x5 & ~n11919 ;
  assign n11922 = ( ~n11918 & n11920 ) | ( ~n11918 & n11921 ) | ( n11920 & n11921 ) ;
  assign n11923 = ( ~n10977 & n10987 ) | ( ~n10977 & n10989 ) | ( n10987 & n10989 ) ;
  assign n11924 = ( n10977 & ~n10990 ) | ( n10977 & n11923 ) | ( ~n10990 & n11923 ) ;
  assign n11925 = ( n11912 & n11922 ) | ( n11912 & n11924 ) | ( n11922 & n11924 ) ;
  assign n11926 = n40 & n10265 ;
  assign n11927 = n8721 & n10267 ;
  assign n11928 = n8340 & ~n10269 ;
  assign n11929 = n11927 | n11928 ;
  assign n11930 = n11926 | n11929 ;
  assign n11931 = x5 & n11930 ;
  assign n11932 = n8341 & n10804 ;
  assign n11933 = ( ~x5 & n11930 ) | ( ~x5 & n11932 ) | ( n11930 & n11932 ) ;
  assign n11934 = x5 & ~n11932 ;
  assign n11935 = ( ~n11931 & n11933 ) | ( ~n11931 & n11934 ) | ( n11933 & n11934 ) ;
  assign n11936 = ( ~n10990 & n10992 ) | ( ~n10990 & n11002 ) | ( n10992 & n11002 ) ;
  assign n11937 = ( n10990 & ~n11003 ) | ( n10990 & n11936 ) | ( ~n11003 & n11936 ) ;
  assign n11938 = ( n11925 & n11935 ) | ( n11925 & n11937 ) | ( n11935 & n11937 ) ;
  assign n11939 = n40 & n10263 ;
  assign n11940 = n8721 & n10265 ;
  assign n11941 = n8340 & n10267 ;
  assign n11942 = n11940 | n11941 ;
  assign n11943 = n11939 | n11942 ;
  assign n11944 = x5 & n11943 ;
  assign n11945 = n8341 & n10874 ;
  assign n11946 = ( ~x5 & n11943 ) | ( ~x5 & n11945 ) | ( n11943 & n11945 ) ;
  assign n11947 = x5 & ~n11945 ;
  assign n11948 = ( ~n11944 & n11946 ) | ( ~n11944 & n11947 ) | ( n11946 & n11947 ) ;
  assign n11949 = ( ~n11003 & n11005 ) | ( ~n11003 & n11015 ) | ( n11005 & n11015 ) ;
  assign n11950 = ( n11003 & ~n11016 ) | ( n11003 & n11949 ) | ( ~n11016 & n11949 ) ;
  assign n11951 = ( n11938 & n11948 ) | ( n11938 & n11950 ) | ( n11948 & n11950 ) ;
  assign n11952 = ( n11787 & n11789 ) | ( n11787 & n11951 ) | ( n11789 & n11951 ) ;
  assign n11953 = ( n11775 & n11777 ) | ( n11775 & n11952 ) | ( n11777 & n11952 ) ;
  assign n11954 = ( n11763 & n11765 ) | ( n11763 & n11953 ) | ( n11765 & n11953 ) ;
  assign n11955 = ( n11751 & n11753 ) | ( n11751 & n11954 ) | ( n11753 & n11954 ) ;
  assign n11956 = ( n11739 & n11741 ) | ( n11739 & n11955 ) | ( n11741 & n11955 ) ;
  assign n11957 = ( ~n11061 & n11075 ) | ( ~n11061 & n11144 ) | ( n11075 & n11144 ) ;
  assign n11958 = ( n11061 & ~n11145 ) | ( n11061 & n11957 ) | ( ~n11145 & n11957 ) ;
  assign n11959 = ( n11729 & n11956 ) | ( n11729 & n11958 ) | ( n11956 & n11958 ) ;
  assign n11960 = ( n11717 & n11719 ) | ( n11717 & n11959 ) | ( n11719 & n11959 ) ;
  assign n11961 = ( n11705 & n11707 ) | ( n11705 & n11960 ) | ( n11707 & n11960 ) ;
  assign n11962 = n40 & n10247 ;
  assign n11963 = n8721 & n10312 ;
  assign n11964 = n8340 & ~n10249 ;
  assign n11965 = n11963 | n11964 ;
  assign n11966 = n11962 | n11965 ;
  assign n11967 = x5 & n11966 ;
  assign n11968 = n8341 & n10428 ;
  assign n11969 = ( ~x5 & n11966 ) | ( ~x5 & n11968 ) | ( n11966 & n11968 ) ;
  assign n11970 = x5 & ~n11968 ;
  assign n11971 = ( ~n11967 & n11969 ) | ( ~n11967 & n11970 ) | ( n11969 & n11970 ) ;
  assign n11972 = ( ~n11306 & n11319 ) | ( ~n11306 & n11397 ) | ( n11319 & n11397 ) ;
  assign n11973 = ( n11306 & ~n11398 ) | ( n11306 & n11972 ) | ( ~n11398 & n11972 ) ;
  assign n11974 = ( n11961 & n11971 ) | ( n11961 & n11973 ) | ( n11971 & n11973 ) ;
  assign n11975 = ( ~n10449 & n11398 ) | ( ~n10449 & n11475 ) | ( n11398 & n11475 ) ;
  assign n11976 = ( n10449 & ~n11476 ) | ( n10449 & n11975 ) | ( ~n11476 & n11975 ) ;
  assign n11977 = ( n11695 & n11974 ) | ( n11695 & n11976 ) | ( n11974 & n11976 ) ;
  assign n11978 = ( n11680 & n11682 ) | ( n11680 & n11977 ) | ( n11682 & n11977 ) ;
  assign n11979 = ( n10422 & n11666 ) | ( n10422 & n11978 ) | ( n11666 & n11978 ) ;
  assign n11980 = n40 & n10243 ;
  assign n11981 = n8721 & ~n10320 ;
  assign n11982 = n8340 & n10245 ;
  assign n11983 = n11981 | n11982 ;
  assign n11984 = n11980 | n11983 ;
  assign n11985 = x5 & n11984 ;
  assign n11986 = n10243 & n10359 ;
  assign n11987 = n10243 & ~n10321 ;
  assign n11988 = ( ~n10243 & n10321 ) | ( ~n10243 & n10359 ) | ( n10321 & n10359 ) ;
  assign n11989 = ( ~n11986 & n11987 ) | ( ~n11986 & n11988 ) | ( n11987 & n11988 ) ;
  assign n11990 = n8341 & ~n11989 ;
  assign n11991 = ( ~x5 & n11984 ) | ( ~x5 & n11990 ) | ( n11984 & n11990 ) ;
  assign n11992 = x5 & ~n11990 ;
  assign n11993 = ( ~n11985 & n11991 ) | ( ~n11985 & n11992 ) | ( n11991 & n11992 ) ;
  assign n11994 = n7346 & ~n11691 ;
  assign n11995 = x8 & n11994 ;
  assign n11996 = n7341 & n10312 ;
  assign n11997 = n7345 | n11996 ;
  assign n11998 = ( ~n10316 & n11996 ) | ( ~n10316 & n11997 ) | ( n11996 & n11997 ) ;
  assign n11999 = n7644 & n10247 ;
  assign n12000 = n11998 | n11999 ;
  assign n12001 = x8 & ~n12000 ;
  assign n12002 = ( ~x8 & n11994 ) | ( ~x8 & n12000 ) | ( n11994 & n12000 ) ;
  assign n12003 = ( ~n11995 & n12001 ) | ( ~n11995 & n12002 ) | ( n12001 & n12002 ) ;
  assign n12004 = n6796 & n10251 ;
  assign n12005 = x11 & n12004 ;
  assign n12006 = n6567 & ~n10253 ;
  assign n12007 = n6570 | n12006 ;
  assign n12008 = ( ~n10249 & n12006 ) | ( ~n10249 & n12007 ) | ( n12006 & n12007 ) ;
  assign n12009 = n6571 | n12008 ;
  assign n12010 = ( ~n10441 & n12008 ) | ( ~n10441 & n12009 ) | ( n12008 & n12009 ) ;
  assign n12011 = x11 & ~n12010 ;
  assign n12012 = ( ~x11 & n12004 ) | ( ~x11 & n12010 ) | ( n12004 & n12010 ) ;
  assign n12013 = ( ~n12005 & n12011 ) | ( ~n12005 & n12012 ) | ( n12011 & n12012 ) ;
  assign n12014 = n6332 & n10257 ;
  assign n12015 = x14 & n12014 ;
  assign n12016 = n5909 & n10259 ;
  assign n12017 = n5914 | n12016 ;
  assign n12018 = ( n10255 & n12016 ) | ( n10255 & n12017 ) | ( n12016 & n12017 ) ;
  assign n12019 = n5915 | n12018 ;
  assign n12020 = ( n11148 & n12018 ) | ( n11148 & n12019 ) | ( n12018 & n12019 ) ;
  assign n12021 = x14 & ~n12020 ;
  assign n12022 = ( ~x14 & n12014 ) | ( ~x14 & n12020 ) | ( n12014 & n12020 ) ;
  assign n12023 = ( ~n12015 & n12021 ) | ( ~n12015 & n12022 ) | ( n12021 & n12022 ) ;
  assign n12024 = n5584 & n10263 ;
  assign n12025 = x17 & n12024 ;
  assign n12026 = n5413 & n10265 ;
  assign n12027 = n5417 | n12026 ;
  assign n12028 = ( n10261 & n12026 ) | ( n10261 & n12027 ) | ( n12026 & n12027 ) ;
  assign n12029 = n5418 | n12028 ;
  assign n12030 = ( n11049 & n12028 ) | ( n11049 & n12029 ) | ( n12028 & n12029 ) ;
  assign n12031 = x17 & ~n12030 ;
  assign n12032 = ( ~x17 & n12024 ) | ( ~x17 & n12030 ) | ( n12024 & n12030 ) ;
  assign n12033 = ( ~n12025 & n12031 ) | ( ~n12025 & n12032 ) | ( n12031 & n12032 ) ;
  assign n12034 = n4879 & ~n10787 ;
  assign n12035 = x20 & n12034 ;
  assign n12036 = n4874 & n10271 ;
  assign n12037 = n4878 | n12036 ;
  assign n12038 = ( n10267 & n12036 ) | ( n10267 & n12037 ) | ( n12036 & n12037 ) ;
  assign n12039 = n5232 & ~n10269 ;
  assign n12040 = n12038 | n12039 ;
  assign n12041 = x20 & ~n12040 ;
  assign n12042 = ( ~x20 & n12034 ) | ( ~x20 & n12040 ) | ( n12034 & n12040 ) ;
  assign n12043 = ( ~n12035 & n12041 ) | ( ~n12035 & n12042 ) | ( n12041 & n12042 ) ;
  assign n12044 = n4637 & n10273 ;
  assign n12045 = x23 & n12044 ;
  assign n12046 = n4584 & n10275 ;
  assign n12047 = n4649 | n12046 ;
  assign n12048 = ( ~n10297 & n12046 ) | ( ~n10297 & n12047 ) | ( n12046 & n12047 ) ;
  assign n12049 = n4591 | n12048 ;
  assign n12050 = ( ~n10617 & n12048 ) | ( ~n10617 & n12049 ) | ( n12048 & n12049 ) ;
  assign n12051 = x23 & ~n12050 ;
  assign n12052 = ( ~x23 & n12044 ) | ( ~x23 & n12050 ) | ( n12044 & n12050 ) ;
  assign n12053 = ( ~n12045 & n12051 ) | ( ~n12045 & n12052 ) | ( n12051 & n12052 ) ;
  assign n12054 = n3541 & n10464 ;
  assign n12055 = n4039 & n10281 ;
  assign n12056 = n3501 & ~n10283 ;
  assign n12057 = n3536 & ~n10285 ;
  assign n12058 = n12056 | n12057 ;
  assign n12059 = n12055 | n12058 ;
  assign n12060 = n12054 | n12059 ;
  assign n12061 = x29 & n11632 ;
  assign n12062 = ~n12060 & n12061 ;
  assign n12063 = n12060 & ~n12061 ;
  assign n12064 = n12062 | n12063 ;
  assign n12065 = n4215 & n10277 ;
  assign n12066 = n4200 & n10291 ;
  assign n12067 = n2083 & ~n10279 ;
  assign n12068 = n12066 | n12067 ;
  assign n12069 = n12065 | n12068 ;
  assign n12070 = x26 & n12069 ;
  assign n12071 = n4203 & ~n10516 ;
  assign n12072 = ( ~x26 & n12069 ) | ( ~x26 & n12071 ) | ( n12069 & n12071 ) ;
  assign n12073 = x26 & ~n12071 ;
  assign n12074 = ( ~n12070 & n12072 ) | ( ~n12070 & n12073 ) | ( n12072 & n12073 ) ;
  assign n12075 = ( ~n11637 & n12064 ) | ( ~n11637 & n12074 ) | ( n12064 & n12074 ) ;
  assign n12076 = ( n11637 & n12064 ) | ( n11637 & n12074 ) | ( n12064 & n12074 ) ;
  assign n12077 = ( n11637 & n12075 ) | ( n11637 & ~n12076 ) | ( n12075 & ~n12076 ) ;
  assign n12078 = ( ~n11640 & n12053 ) | ( ~n11640 & n12077 ) | ( n12053 & n12077 ) ;
  assign n12079 = ( n11640 & n12053 ) | ( n11640 & n12077 ) | ( n12053 & n12077 ) ;
  assign n12080 = ( n11640 & n12078 ) | ( n11640 & ~n12079 ) | ( n12078 & ~n12079 ) ;
  assign n12081 = ( ~n11642 & n12043 ) | ( ~n11642 & n12080 ) | ( n12043 & n12080 ) ;
  assign n12082 = ( n11642 & n12043 ) | ( n11642 & n12080 ) | ( n12043 & n12080 ) ;
  assign n12083 = ( n11642 & n12081 ) | ( n11642 & ~n12082 ) | ( n12081 & ~n12082 ) ;
  assign n12084 = ( ~n11656 & n12033 ) | ( ~n11656 & n12083 ) | ( n12033 & n12083 ) ;
  assign n12085 = ( n11656 & n12033 ) | ( n11656 & n12083 ) | ( n12033 & n12083 ) ;
  assign n12086 = ( n11656 & n12084 ) | ( n11656 & ~n12085 ) | ( n12084 & ~n12085 ) ;
  assign n12087 = ( ~n11659 & n12023 ) | ( ~n11659 & n12086 ) | ( n12023 & n12086 ) ;
  assign n12088 = ( n11659 & n12023 ) | ( n11659 & n12086 ) | ( n12023 & n12086 ) ;
  assign n12089 = ( n11659 & n12087 ) | ( n11659 & ~n12088 ) | ( n12087 & ~n12088 ) ;
  assign n12090 = ( ~n11662 & n12013 ) | ( ~n11662 & n12089 ) | ( n12013 & n12089 ) ;
  assign n12091 = ( n11662 & n12013 ) | ( n11662 & n12089 ) | ( n12013 & n12089 ) ;
  assign n12092 = ( n11662 & n12090 ) | ( n11662 & ~n12091 ) | ( n12090 & ~n12091 ) ;
  assign n12093 = ( n11664 & ~n12003 ) | ( n11664 & n12092 ) | ( ~n12003 & n12092 ) ;
  assign n12094 = ( n11664 & n12003 ) | ( n11664 & n12092 ) | ( n12003 & n12092 ) ;
  assign n12095 = ( n12003 & n12093 ) | ( n12003 & ~n12094 ) | ( n12093 & ~n12094 ) ;
  assign n12096 = ( n11979 & n11993 ) | ( n11979 & n12095 ) | ( n11993 & n12095 ) ;
  assign n12097 = n40 & n10241 ;
  assign n12098 = n8721 & n10243 ;
  assign n12099 = n8340 & ~n10320 ;
  assign n12100 = n12098 | n12099 ;
  assign n12101 = n12097 | n12100 ;
  assign n12102 = x5 & n12101 ;
  assign n12103 = n10322 & ~n10361 ;
  assign n12104 = ( ~n10243 & n10323 ) | ( ~n10243 & n11986 ) | ( n10323 & n11986 ) ;
  assign n12105 = ( n10241 & n12103 ) | ( n10241 & ~n12104 ) | ( n12103 & ~n12104 ) ;
  assign n12106 = n8341 & n12105 ;
  assign n12107 = ( ~x5 & n12101 ) | ( ~x5 & n12106 ) | ( n12101 & n12106 ) ;
  assign n12108 = x5 & ~n12106 ;
  assign n12109 = ( ~n12102 & n12107 ) | ( ~n12102 & n12108 ) | ( n12107 & n12108 ) ;
  assign n12110 = n7644 & ~n10316 ;
  assign n12111 = x8 & n12110 ;
  assign n12112 = n7341 & n10247 ;
  assign n12113 = n7345 | n12112 ;
  assign n12114 = ( n10245 & n12112 ) | ( n10245 & n12113 ) | ( n12112 & n12113 ) ;
  assign n12115 = n7346 | n12114 ;
  assign n12116 = ( ~n11676 & n12114 ) | ( ~n11676 & n12115 ) | ( n12114 & n12115 ) ;
  assign n12117 = x8 & ~n12116 ;
  assign n12118 = ( ~x8 & n12110 ) | ( ~x8 & n12116 ) | ( n12110 & n12116 ) ;
  assign n12119 = ( ~n12111 & n12117 ) | ( ~n12111 & n12118 ) | ( n12117 & n12118 ) ;
  assign n12120 = n6570 & n10312 ;
  assign n12121 = x11 & n12120 ;
  assign n12122 = n6796 & ~n10249 ;
  assign n12123 = n6567 & n10251 ;
  assign n12124 = n12122 | n12123 ;
  assign n12125 = n6571 | n12124 ;
  assign n12126 = ( ~n11486 & n12124 ) | ( ~n11486 & n12125 ) | ( n12124 & n12125 ) ;
  assign n12127 = x11 & ~n12126 ;
  assign n12128 = ( ~x11 & n12120 ) | ( ~x11 & n12126 ) | ( n12120 & n12126 ) ;
  assign n12129 = ( ~n12121 & n12127 ) | ( ~n12121 & n12128 ) | ( n12127 & n12128 ) ;
  assign n12130 = n6332 & n10255 ;
  assign n12131 = x14 & n12130 ;
  assign n12132 = n5909 & n10257 ;
  assign n12133 = n5914 | n12132 ;
  assign n12134 = ( ~n10253 & n12132 ) | ( ~n10253 & n12133 ) | ( n12132 & n12133 ) ;
  assign n12135 = n5915 | n12134 ;
  assign n12136 = ( ~n11297 & n12134 ) | ( ~n11297 & n12135 ) | ( n12134 & n12135 ) ;
  assign n12137 = x14 & ~n12136 ;
  assign n12138 = ( ~x14 & n12130 ) | ( ~x14 & n12136 ) | ( n12130 & n12136 ) ;
  assign n12139 = ( ~n12131 & n12137 ) | ( ~n12131 & n12138 ) | ( n12137 & n12138 ) ;
  assign n12140 = n5584 & n10261 ;
  assign n12141 = x17 & n12140 ;
  assign n12142 = n5413 & n10263 ;
  assign n12143 = n5417 | n12142 ;
  assign n12144 = ( n10259 & n12142 ) | ( n10259 & n12143 ) | ( n12142 & n12143 ) ;
  assign n12145 = n5418 | n12144 ;
  assign n12146 = ( n10859 & n12144 ) | ( n10859 & n12145 ) | ( n12144 & n12145 ) ;
  assign n12147 = x17 & ~n12146 ;
  assign n12148 = ( ~x17 & n12140 ) | ( ~x17 & n12146 ) | ( n12140 & n12146 ) ;
  assign n12149 = ( ~n12141 & n12147 ) | ( ~n12141 & n12148 ) | ( n12147 & n12148 ) ;
  assign n12150 = n5232 & n10267 ;
  assign n12151 = x20 & n12150 ;
  assign n12152 = n4874 & ~n10269 ;
  assign n12153 = n4878 | n12152 ;
  assign n12154 = ( n10265 & n12152 ) | ( n10265 & n12153 ) | ( n12152 & n12153 ) ;
  assign n12155 = n4879 | n12154 ;
  assign n12156 = ( n10804 & n12154 ) | ( n10804 & n12155 ) | ( n12154 & n12155 ) ;
  assign n12157 = x20 & ~n12156 ;
  assign n12158 = ( ~x20 & n12150 ) | ( ~x20 & n12156 ) | ( n12150 & n12156 ) ;
  assign n12159 = ( ~n12151 & n12157 ) | ( ~n12151 & n12158 ) | ( n12157 & n12158 ) ;
  assign n12160 = n4637 & ~n10297 ;
  assign n12161 = x23 & n12160 ;
  assign n12162 = n4584 & n10273 ;
  assign n12163 = n4649 | n12162 ;
  assign n12164 = ( n10271 & n12162 ) | ( n10271 & n12163 ) | ( n12162 & n12163 ) ;
  assign n12165 = n4591 | n12164 ;
  assign n12166 = ( ~n10656 & n12164 ) | ( ~n10656 & n12165 ) | ( n12164 & n12165 ) ;
  assign n12167 = x23 & ~n12166 ;
  assign n12168 = ( ~x23 & n12160 ) | ( ~x23 & n12166 ) | ( n12160 & n12166 ) ;
  assign n12169 = ( ~n12161 & n12167 ) | ( ~n12161 & n12168 ) | ( n12167 & n12168 ) ;
  assign n12170 = n3501 & n10281 ;
  assign n12171 = x29 & n12170 ;
  assign n12172 = n3536 & ~n10283 ;
  assign n12173 = n4039 | n12172 ;
  assign n12174 = ( ~n10279 & n12172 ) | ( ~n10279 & n12173 ) | ( n12172 & n12173 ) ;
  assign n12175 = n3541 | n12174 ;
  assign n12176 = ( n10487 & n12174 ) | ( n10487 & n12175 ) | ( n12174 & n12175 ) ;
  assign n12177 = x29 & ~n12176 ;
  assign n12178 = ( ~x29 & n12170 ) | ( ~x29 & n12176 ) | ( n12170 & n12176 ) ;
  assign n12179 = ( ~n12171 & n12177 ) | ( ~n12171 & n12178 ) | ( n12177 & n12178 ) ;
  assign n12180 = x29 & ~n11632 ;
  assign n12181 = ~n12060 & n12180 ;
  assign n12182 = n389 & ~n10285 ;
  assign n12183 = ( n12179 & n12181 ) | ( n12179 & n12182 ) | ( n12181 & n12182 ) ;
  assign n12184 = ( ~n12179 & n12181 ) | ( ~n12179 & n12182 ) | ( n12181 & n12182 ) ;
  assign n12185 = ( n12179 & ~n12183 ) | ( n12179 & n12184 ) | ( ~n12183 & n12184 ) ;
  assign n12186 = n4215 & n10275 ;
  assign n12187 = n4200 & n10277 ;
  assign n12188 = n2083 & n10291 ;
  assign n12189 = n12187 | n12188 ;
  assign n12190 = n12186 | n12189 ;
  assign n12191 = x26 & n12190 ;
  assign n12192 = n4203 & n10563 ;
  assign n12193 = ( ~x26 & n12190 ) | ( ~x26 & n12192 ) | ( n12190 & n12192 ) ;
  assign n12194 = x26 & ~n12192 ;
  assign n12195 = ( ~n12191 & n12193 ) | ( ~n12191 & n12194 ) | ( n12193 & n12194 ) ;
  assign n12196 = ( ~n12076 & n12185 ) | ( ~n12076 & n12195 ) | ( n12185 & n12195 ) ;
  assign n12197 = ( n12076 & n12185 ) | ( n12076 & n12195 ) | ( n12185 & n12195 ) ;
  assign n12198 = ( n12076 & n12196 ) | ( n12076 & ~n12197 ) | ( n12196 & ~n12197 ) ;
  assign n12199 = ( ~n12079 & n12169 ) | ( ~n12079 & n12198 ) | ( n12169 & n12198 ) ;
  assign n12200 = ( n12079 & n12169 ) | ( n12079 & n12198 ) | ( n12169 & n12198 ) ;
  assign n12201 = ( n12079 & n12199 ) | ( n12079 & ~n12200 ) | ( n12199 & ~n12200 ) ;
  assign n12202 = ( ~n12082 & n12159 ) | ( ~n12082 & n12201 ) | ( n12159 & n12201 ) ;
  assign n12203 = ( n12082 & n12159 ) | ( n12082 & n12201 ) | ( n12159 & n12201 ) ;
  assign n12204 = ( n12082 & n12202 ) | ( n12082 & ~n12203 ) | ( n12202 & ~n12203 ) ;
  assign n12205 = ( ~n12085 & n12149 ) | ( ~n12085 & n12204 ) | ( n12149 & n12204 ) ;
  assign n12206 = ( n12085 & n12149 ) | ( n12085 & n12204 ) | ( n12149 & n12204 ) ;
  assign n12207 = ( n12085 & n12205 ) | ( n12085 & ~n12206 ) | ( n12205 & ~n12206 ) ;
  assign n12208 = ( ~n12088 & n12139 ) | ( ~n12088 & n12207 ) | ( n12139 & n12207 ) ;
  assign n12209 = ( n12088 & n12139 ) | ( n12088 & n12207 ) | ( n12139 & n12207 ) ;
  assign n12210 = ( n12088 & n12208 ) | ( n12088 & ~n12209 ) | ( n12208 & ~n12209 ) ;
  assign n12211 = ( ~n12091 & n12129 ) | ( ~n12091 & n12210 ) | ( n12129 & n12210 ) ;
  assign n12212 = ( n12091 & n12129 ) | ( n12091 & n12210 ) | ( n12129 & n12210 ) ;
  assign n12213 = ( n12091 & n12211 ) | ( n12091 & ~n12212 ) | ( n12211 & ~n12212 ) ;
  assign n12214 = ( ~n12094 & n12119 ) | ( ~n12094 & n12213 ) | ( n12119 & n12213 ) ;
  assign n12215 = ( n12094 & n12119 ) | ( n12094 & n12213 ) | ( n12119 & n12213 ) ;
  assign n12216 = ( n12094 & n12214 ) | ( n12094 & ~n12215 ) | ( n12214 & ~n12215 ) ;
  assign n12217 = ( ~n12096 & n12109 ) | ( ~n12096 & n12216 ) | ( n12109 & n12216 ) ;
  assign n12218 = ( n12096 & n12109 ) | ( n12096 & n12216 ) | ( n12109 & n12216 ) ;
  assign n12219 = ( n12096 & n12217 ) | ( n12096 & ~n12218 ) | ( n12217 & ~n12218 ) ;
  assign n12220 = n10326 & n10362 ;
  assign n12221 = ( n10324 & n10326 ) | ( n10324 & ~n10362 ) | ( n10326 & ~n10362 ) ;
  assign n12222 = ( ~n10327 & n12220 ) | ( ~n10327 & n12221 ) | ( n12220 & n12221 ) ;
  assign n12223 = n9593 & n10326 ;
  assign n12224 = n9592 | n12223 ;
  assign n12225 = ( n12222 & n12223 ) | ( n12222 & n12224 ) | ( n12223 & n12224 ) ;
  assign n12226 = n41 & n10239 ;
  assign n12227 = ( x2 & ~n12225 ) | ( x2 & n12226 ) | ( ~n12225 & n12226 ) ;
  assign n12228 = ~x2 & n12225 ;
  assign n12229 = ~n9154 & n10241 ;
  assign n12230 = n12226 & ~n12229 ;
  assign n12231 = ( x2 & n12229 ) | ( x2 & n12230 ) | ( n12229 & n12230 ) ;
  assign n12232 = ( n12227 & n12228 ) | ( n12227 & ~n12231 ) | ( n12228 & ~n12231 ) ;
  assign n12233 = n41 & n10247 ;
  assign n12234 = n9592 | n12233 ;
  assign n12235 = ( ~n11691 & n12233 ) | ( ~n11691 & n12234 ) | ( n12233 & n12234 ) ;
  assign n12236 = n9593 & ~n10316 ;
  assign n12237 = ( x2 & ~n12235 ) | ( x2 & n12236 ) | ( ~n12235 & n12236 ) ;
  assign n12238 = ~x2 & n12235 ;
  assign n12239 = n9600 & n10312 ;
  assign n12240 = ( x2 & n12236 ) | ( x2 & n12239 ) | ( n12236 & n12239 ) ;
  assign n12241 = ( n12237 & n12238 ) | ( n12237 & ~n12240 ) | ( n12238 & ~n12240 ) ;
  assign n12242 = ( ~n11717 & n11719 ) | ( ~n11717 & n11959 ) | ( n11719 & n11959 ) ;
  assign n12243 = ( n11717 & ~n11960 ) | ( n11717 & n12242 ) | ( ~n11960 & n12242 ) ;
  assign n12244 = n9592 & ~n11486 ;
  assign n12245 = n9593 & n10312 ;
  assign n12246 = n41 & ~n10249 ;
  assign n12247 = n12245 | n12246 ;
  assign n12248 = x2 | n12247 ;
  assign n12249 = ( ~n12244 & n12247 ) | ( ~n12244 & n12248 ) | ( n12247 & n12248 ) ;
  assign n12250 = n9591 & ~n11486 ;
  assign n12251 = n12249 | n12250 ;
  assign n12252 = n9600 & n10251 ;
  assign n12253 = ( x2 & n12247 ) | ( x2 & n12252 ) | ( n12247 & n12252 ) ;
  assign n12254 = n12251 & ~n12253 ;
  assign n12255 = ( ~n11739 & n11741 ) | ( ~n11739 & n11955 ) | ( n11741 & n11955 ) ;
  assign n12256 = ( n11739 & ~n11956 ) | ( n11739 & n12255 ) | ( ~n11956 & n12255 ) ;
  assign n12257 = n9592 & ~n10698 ;
  assign n12258 = n9593 & ~n10269 ;
  assign n12259 = n41 & n10271 ;
  assign n12260 = n12258 | n12259 ;
  assign n12261 = x2 | n12260 ;
  assign n12262 = ( ~n12257 & n12260 ) | ( ~n12257 & n12261 ) | ( n12260 & n12261 ) ;
  assign n12263 = n9591 & ~n10698 ;
  assign n12264 = n12262 | n12263 ;
  assign n12265 = n9600 & ~n10297 ;
  assign n12266 = ( x2 & n12260 ) | ( x2 & n12265 ) | ( n12260 & n12265 ) ;
  assign n12267 = n12264 & ~n12266 ;
  assign n12268 = ( ~n11860 & n11870 ) | ( ~n11860 & n11872 ) | ( n11870 & n11872 ) ;
  assign n12269 = ( n11860 & ~n11873 ) | ( n11860 & n12268 ) | ( ~n11873 & n12268 ) ;
  assign n12270 = n9593 & n10271 ;
  assign n12271 = n41 & ~n10297 ;
  assign n12272 = n12270 | n12271 ;
  assign n12273 = n9639 | n12272 ;
  assign n12274 = ~x2 & n10656 ;
  assign n12275 = n9158 | n10656 ;
  assign n12276 = ( n12273 & ~n12274 ) | ( n12273 & n12275 ) | ( ~n12274 & n12275 ) ;
  assign n12277 = n9600 & n10273 ;
  assign n12278 = ( x2 & n12272 ) | ( x2 & n12277 ) | ( n12272 & n12277 ) ;
  assign n12279 = n12276 & ~n12278 ;
  assign n12280 = ( n10930 & ~n11849 ) | ( n10930 & n11859 ) | ( ~n11849 & n11859 ) ;
  assign n12281 = ( n11849 & ~n11860 ) | ( n11849 & n12280 ) | ( ~n11860 & n12280 ) ;
  assign n12282 = n41 & n10275 ;
  assign n12283 = x2 & n12282 ;
  assign n12284 = n9600 & n10277 ;
  assign n12285 = n9593 | n12284 ;
  assign n12286 = ( n10273 & n12284 ) | ( n10273 & n12285 ) | ( n12284 & n12285 ) ;
  assign n12287 = n9592 | n12286 ;
  assign n12288 = ( n10577 & n12286 ) | ( n10577 & n12287 ) | ( n12286 & n12287 ) ;
  assign n12289 = x2 & ~n12288 ;
  assign n12290 = ( ~x2 & n12282 ) | ( ~x2 & n12288 ) | ( n12282 & n12288 ) ;
  assign n12291 = ( ~n12283 & n12289 ) | ( ~n12283 & n12290 ) | ( n12289 & n12290 ) ;
  assign n12292 = ( ~n11799 & n11801 ) | ( ~n11799 & n11833 ) | ( n11801 & n11833 ) ;
  assign n12293 = ( n11799 & ~n11834 ) | ( n11799 & n12292 ) | ( ~n11834 & n12292 ) ;
  assign n12294 = n41 & n10277 ;
  assign n12295 = x2 & n12294 ;
  assign n12296 = n9600 & n10291 ;
  assign n12297 = n9593 | n12296 ;
  assign n12298 = ( n10275 & n12296 ) | ( n10275 & n12297 ) | ( n12296 & n12297 ) ;
  assign n12299 = n9592 | n12298 ;
  assign n12300 = ( n10563 & n12298 ) | ( n10563 & n12299 ) | ( n12298 & n12299 ) ;
  assign n12301 = x2 & ~n12300 ;
  assign n12302 = ( ~x2 & n12294 ) | ( ~x2 & n12300 ) | ( n12294 & n12300 ) ;
  assign n12303 = ( ~n12295 & n12301 ) | ( ~n12295 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12304 = n9593 & n10291 ;
  assign n12305 = n41 & ~n10279 ;
  assign n12306 = n12304 | n12305 ;
  assign n12307 = x2 & n12306 ;
  assign n12308 = ~x2 & n12306 ;
  assign n12309 = n9600 & n10281 ;
  assign n12310 = ( x2 & n9590 ) | ( x2 & ~n10454 ) | ( n9590 & ~n10454 ) ;
  assign n12311 = n9591 & n10454 ;
  assign n12312 = ( ~n12309 & n12310 ) | ( ~n12309 & n12311 ) | ( n12310 & n12311 ) ;
  assign n12313 = ( ~n12307 & n12308 ) | ( ~n12307 & n12312 ) | ( n12308 & n12312 ) ;
  assign n12314 = ~n11807 & n11809 ;
  assign n12315 = n11807 & ~n11809 ;
  assign n12316 = n12314 | n12315 ;
  assign n12317 = n9593 & ~n10279 ;
  assign n12318 = n9592 | n12317 ;
  assign n12319 = ( n10487 & n12317 ) | ( n10487 & n12318 ) | ( n12317 & n12318 ) ;
  assign n12320 = n41 & n10281 ;
  assign n12321 = n12319 | n12320 ;
  assign n12322 = x0 & n10285 ;
  assign n12323 = n10281 & n12322 ;
  assign n12324 = n36 | n10285 ;
  assign n12325 = x2 | n9154 ;
  assign n12326 = n12324 & ~n12325 ;
  assign n12327 = ( ~n34 & n35 ) | ( ~n34 & n9155 ) | ( n35 & n9155 ) ;
  assign n12328 = ( n10283 & ~n10286 ) | ( n10283 & n12327 ) | ( ~n10286 & n12327 ) ;
  assign n12329 = ( n12324 & n12326 ) | ( n12324 & n12328 ) | ( n12326 & n12328 ) ;
  assign n12330 = ~n12323 & n12329 ;
  assign n12331 = ( x2 & n12321 ) | ( x2 & n12330 ) | ( n12321 & n12330 ) ;
  assign n12332 = x2 | n10285 ;
  assign n12333 = n12321 & n12332 ;
  assign n12334 = n12331 & ~n12333 ;
  assign n12335 = ( n12313 & n12316 ) | ( n12313 & n12334 ) | ( n12316 & n12334 ) ;
  assign n12336 = n9593 & n10277 ;
  assign n12337 = n9592 | n12336 ;
  assign n12338 = ( ~n10516 & n12336 ) | ( ~n10516 & n12337 ) | ( n12336 & n12337 ) ;
  assign n12339 = n41 & n10291 ;
  assign n12340 = ( x2 & ~n12338 ) | ( x2 & n12339 ) | ( ~n12338 & n12339 ) ;
  assign n12341 = ~x2 & n12338 ;
  assign n12342 = n9600 & ~n10279 ;
  assign n12343 = ( x2 & n12339 ) | ( x2 & n12342 ) | ( n12339 & n12342 ) ;
  assign n12344 = ( n12340 & n12341 ) | ( n12340 & ~n12343 ) | ( n12341 & ~n12343 ) ;
  assign n12345 = x5 & n11810 ;
  assign n12346 = ~n11818 & n12345 ;
  assign n12347 = n11818 & ~n12345 ;
  assign n12348 = n12346 | n12347 ;
  assign n12349 = ( n12335 & n12344 ) | ( n12335 & n12348 ) | ( n12344 & n12348 ) ;
  assign n12350 = ( n11831 & n12303 ) | ( n11831 & n12349 ) | ( n12303 & n12349 ) ;
  assign n12351 = ( n12291 & n12293 ) | ( n12291 & n12350 ) | ( n12293 & n12350 ) ;
  assign n12352 = n41 & n10273 ;
  assign n12353 = x2 & n12352 ;
  assign n12354 = n9600 & n10275 ;
  assign n12355 = n9593 | n12354 ;
  assign n12356 = ( ~n10297 & n12354 ) | ( ~n10297 & n12355 ) | ( n12354 & n12355 ) ;
  assign n12357 = n9592 | n12356 ;
  assign n12358 = ( ~n10617 & n12356 ) | ( ~n10617 & n12357 ) | ( n12356 & n12357 ) ;
  assign n12359 = x2 & ~n12358 ;
  assign n12360 = ( ~x2 & n12352 ) | ( ~x2 & n12358 ) | ( n12352 & n12358 ) ;
  assign n12361 = ( ~n12353 & n12359 ) | ( ~n12353 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12362 = ( ~n11834 & n11844 ) | ( ~n11834 & n11848 ) | ( n11844 & n11848 ) ;
  assign n12363 = ( n11834 & ~n11849 ) | ( n11834 & n12362 ) | ( ~n11849 & n12362 ) ;
  assign n12364 = ( n12351 & n12361 ) | ( n12351 & n12363 ) | ( n12361 & n12363 ) ;
  assign n12365 = ( n12279 & n12281 ) | ( n12279 & n12364 ) | ( n12281 & n12364 ) ;
  assign n12366 = ( n12267 & n12269 ) | ( n12267 & n12365 ) | ( n12269 & n12365 ) ;
  assign n12367 = ( ~n11873 & n11883 ) | ( ~n11873 & n11885 ) | ( n11883 & n11885 ) ;
  assign n12368 = ( n11873 & ~n11886 ) | ( n11873 & n12367 ) | ( ~n11886 & n12367 ) ;
  assign n12369 = n9592 & ~n10787 ;
  assign n12370 = x2 & n12369 ;
  assign n12371 = n9600 & n10271 ;
  assign n12372 = n9593 | n12371 ;
  assign n12373 = ( n10267 & n12371 ) | ( n10267 & n12372 ) | ( n12371 & n12372 ) ;
  assign n12374 = n41 & ~n10269 ;
  assign n12375 = n12373 | n12374 ;
  assign n12376 = x2 & ~n12375 ;
  assign n12377 = ( ~x2 & n12369 ) | ( ~x2 & n12375 ) | ( n12369 & n12375 ) ;
  assign n12378 = ( ~n12370 & n12376 ) | ( ~n12370 & n12377 ) | ( n12376 & n12377 ) ;
  assign n12379 = ( n12366 & n12368 ) | ( n12366 & n12378 ) | ( n12368 & n12378 ) ;
  assign n12380 = n9592 & n10804 ;
  assign n12381 = n9593 & n10265 ;
  assign n12382 = n41 & n10267 ;
  assign n12383 = n12381 | n12382 ;
  assign n12384 = x2 | n12383 ;
  assign n12385 = ( ~n12380 & n12383 ) | ( ~n12380 & n12384 ) | ( n12383 & n12384 ) ;
  assign n12386 = n9591 & n10804 ;
  assign n12387 = n12385 | n12386 ;
  assign n12388 = n9600 & ~n10269 ;
  assign n12389 = ( x2 & n12383 ) | ( x2 & n12388 ) | ( n12383 & n12388 ) ;
  assign n12390 = n12387 & ~n12389 ;
  assign n12391 = ( ~n11886 & n11896 ) | ( ~n11886 & n11898 ) | ( n11896 & n11898 ) ;
  assign n12392 = ( n11886 & ~n11899 ) | ( n11886 & n12391 ) | ( ~n11899 & n12391 ) ;
  assign n12393 = ( n12379 & n12390 ) | ( n12379 & n12392 ) | ( n12390 & n12392 ) ;
  assign n12394 = n9600 & n10267 ;
  assign n12395 = n9593 & n10263 ;
  assign n12396 = n41 & n10265 ;
  assign n12397 = n12395 | n12396 ;
  assign n12398 = ~x2 & n12397 ;
  assign n12399 = ( x2 & n9590 ) | ( x2 & ~n10874 ) | ( n9590 & ~n10874 ) ;
  assign n12400 = n9591 & n10874 ;
  assign n12401 = ( ~n12397 & n12399 ) | ( ~n12397 & n12400 ) | ( n12399 & n12400 ) ;
  assign n12402 = ( ~n12394 & n12398 ) | ( ~n12394 & n12401 ) | ( n12398 & n12401 ) ;
  assign n12403 = ( ~n11899 & n11901 ) | ( ~n11899 & n11911 ) | ( n11901 & n11911 ) ;
  assign n12404 = ( n11899 & ~n11912 ) | ( n11899 & n12403 ) | ( ~n11912 & n12403 ) ;
  assign n12405 = ( n12393 & n12402 ) | ( n12393 & n12404 ) | ( n12402 & n12404 ) ;
  assign n12406 = n9593 & n10261 ;
  assign n12407 = n41 & n10263 ;
  assign n12408 = n12406 | n12407 ;
  assign n12409 = n9639 | n12408 ;
  assign n12410 = x2 | n11049 ;
  assign n12411 = ~n9158 & n11049 ;
  assign n12412 = ( n12409 & n12410 ) | ( n12409 & ~n12411 ) | ( n12410 & ~n12411 ) ;
  assign n12413 = n9600 & n10265 ;
  assign n12414 = ( x2 & n12408 ) | ( x2 & n12413 ) | ( n12408 & n12413 ) ;
  assign n12415 = n12412 & ~n12414 ;
  assign n12416 = ( ~n11912 & n11922 ) | ( ~n11912 & n11924 ) | ( n11922 & n11924 ) ;
  assign n12417 = ( n11912 & ~n11925 ) | ( n11912 & n12416 ) | ( ~n11925 & n12416 ) ;
  assign n12418 = ( n12405 & n12415 ) | ( n12405 & n12417 ) | ( n12415 & n12417 ) ;
  assign n12419 = ( ~n11925 & n11935 ) | ( ~n11925 & n11937 ) | ( n11935 & n11937 ) ;
  assign n12420 = ( n11925 & ~n11938 ) | ( n11925 & n12419 ) | ( ~n11938 & n12419 ) ;
  assign n12421 = n9592 & n10859 ;
  assign n12422 = n9593 & n10259 ;
  assign n12423 = n41 & n10261 ;
  assign n12424 = n12422 | n12423 ;
  assign n12425 = x2 | n12424 ;
  assign n12426 = ( ~n12421 & n12424 ) | ( ~n12421 & n12425 ) | ( n12424 & n12425 ) ;
  assign n12427 = n9591 & n10859 ;
  assign n12428 = n12426 | n12427 ;
  assign n12429 = n9600 & n10263 ;
  assign n12430 = ( x2 & n12424 ) | ( x2 & n12429 ) | ( n12424 & n12429 ) ;
  assign n12431 = n12428 & ~n12430 ;
  assign n12432 = ( n12418 & n12420 ) | ( n12418 & n12431 ) | ( n12420 & n12431 ) ;
  assign n12433 = ( ~n11938 & n11948 ) | ( ~n11938 & n11950 ) | ( n11948 & n11950 ) ;
  assign n12434 = ( n11938 & ~n11951 ) | ( n11938 & n12433 ) | ( ~n11951 & n12433 ) ;
  assign n12435 = n41 & n10259 ;
  assign n12436 = x2 & n12435 ;
  assign n12437 = n9600 & n10261 ;
  assign n12438 = n9593 | n12437 ;
  assign n12439 = ( n10257 & n12437 ) | ( n10257 & n12438 ) | ( n12437 & n12438 ) ;
  assign n12440 = n9592 | n12439 ;
  assign n12441 = ( n11065 & n12439 ) | ( n11065 & n12440 ) | ( n12439 & n12440 ) ;
  assign n12442 = x2 & ~n12441 ;
  assign n12443 = ( ~x2 & n12435 ) | ( ~x2 & n12441 ) | ( n12435 & n12441 ) ;
  assign n12444 = ( ~n12436 & n12442 ) | ( ~n12436 & n12443 ) | ( n12442 & n12443 ) ;
  assign n12445 = ( n12432 & n12434 ) | ( n12432 & n12444 ) | ( n12434 & n12444 ) ;
  assign n12446 = ( ~n11787 & n11789 ) | ( ~n11787 & n11951 ) | ( n11789 & n11951 ) ;
  assign n12447 = ( n11787 & ~n11952 ) | ( n11787 & n12446 ) | ( ~n11952 & n12446 ) ;
  assign n12448 = n9593 & n10255 ;
  assign n12449 = n41 & n10257 ;
  assign n12450 = n12448 | n12449 ;
  assign n12451 = n9600 & n10259 ;
  assign n12452 = ( x2 & n12450 ) | ( x2 & n12451 ) | ( n12450 & n12451 ) ;
  assign n12453 = x0 & n11148 ;
  assign n12454 = x2 | n12453 ;
  assign n12455 = ~x1 & n12453 ;
  assign n12456 = ( n12450 & n12454 ) | ( n12450 & ~n12455 ) | ( n12454 & ~n12455 ) ;
  assign n12457 = ~n12452 & n12456 ;
  assign n12458 = ( n12445 & n12447 ) | ( n12445 & n12457 ) | ( n12447 & n12457 ) ;
  assign n12459 = n9592 & ~n11297 ;
  assign n12460 = n9593 & ~n10253 ;
  assign n12461 = n41 & n10255 ;
  assign n12462 = n12460 | n12461 ;
  assign n12463 = x2 | n12462 ;
  assign n12464 = ( ~n12459 & n12462 ) | ( ~n12459 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = n9591 & ~n11297 ;
  assign n12466 = n12464 | n12465 ;
  assign n12467 = n9600 & n10257 ;
  assign n12468 = ( x2 & n12462 ) | ( x2 & n12467 ) | ( n12462 & n12467 ) ;
  assign n12469 = n12466 & ~n12468 ;
  assign n12470 = ( ~n11775 & n11777 ) | ( ~n11775 & n11952 ) | ( n11777 & n11952 ) ;
  assign n12471 = ( n11775 & ~n11953 ) | ( n11775 & n12470 ) | ( ~n11953 & n12470 ) ;
  assign n12472 = ( n12458 & n12469 ) | ( n12458 & n12471 ) | ( n12469 & n12471 ) ;
  assign n12473 = n9593 & n10251 ;
  assign n12474 = n9592 | n12473 ;
  assign n12475 = ( ~n11309 & n12473 ) | ( ~n11309 & n12474 ) | ( n12473 & n12474 ) ;
  assign n12476 = n41 & ~n10253 ;
  assign n12477 = ( x2 & ~n12475 ) | ( x2 & n12476 ) | ( ~n12475 & n12476 ) ;
  assign n12478 = ~x2 & n12475 ;
  assign n12479 = n9600 & n10255 ;
  assign n12480 = ( x2 & n12476 ) | ( x2 & n12479 ) | ( n12476 & n12479 ) ;
  assign n12481 = ( n12477 & n12478 ) | ( n12477 & ~n12480 ) | ( n12478 & ~n12480 ) ;
  assign n12482 = ( ~n11763 & n11765 ) | ( ~n11763 & n11953 ) | ( n11765 & n11953 ) ;
  assign n12483 = ( n11763 & ~n11954 ) | ( n11763 & n12482 ) | ( ~n11954 & n12482 ) ;
  assign n12484 = ( n12472 & n12481 ) | ( n12472 & n12483 ) | ( n12481 & n12483 ) ;
  assign n12485 = n41 & n10251 ;
  assign n12486 = x2 & n12485 ;
  assign n12487 = n9600 & ~n10253 ;
  assign n12488 = n9593 | n12487 ;
  assign n12489 = ( ~n10249 & n12487 ) | ( ~n10249 & n12488 ) | ( n12487 & n12488 ) ;
  assign n12490 = n9592 | n12489 ;
  assign n12491 = ( ~n10441 & n12489 ) | ( ~n10441 & n12490 ) | ( n12489 & n12490 ) ;
  assign n12492 = x2 & ~n12491 ;
  assign n12493 = ( ~x2 & n12485 ) | ( ~x2 & n12491 ) | ( n12485 & n12491 ) ;
  assign n12494 = ( ~n12486 & n12492 ) | ( ~n12486 & n12493 ) | ( n12492 & n12493 ) ;
  assign n12495 = ( ~n11751 & n11753 ) | ( ~n11751 & n11954 ) | ( n11753 & n11954 ) ;
  assign n12496 = ( n11751 & ~n11955 ) | ( n11751 & n12495 ) | ( ~n11955 & n12495 ) ;
  assign n12497 = ( n12484 & n12494 ) | ( n12484 & n12496 ) | ( n12494 & n12496 ) ;
  assign n12498 = ( n12254 & n12256 ) | ( n12254 & n12497 ) | ( n12256 & n12497 ) ;
  assign n12499 = ( ~n11729 & n11956 ) | ( ~n11729 & n11958 ) | ( n11956 & n11958 ) ;
  assign n12500 = ( n11729 & ~n11959 ) | ( n11729 & n12499 ) | ( ~n11959 & n12499 ) ;
  assign n12501 = n41 & n10312 ;
  assign n12502 = x2 & n12501 ;
  assign n12503 = n9600 & ~n10249 ;
  assign n12504 = n9593 | n12503 ;
  assign n12505 = ( n10247 & n12503 ) | ( n10247 & n12504 ) | ( n12503 & n12504 ) ;
  assign n12506 = n9592 | n12505 ;
  assign n12507 = ( n10428 & n12505 ) | ( n10428 & n12506 ) | ( n12505 & n12506 ) ;
  assign n12508 = x2 & ~n12507 ;
  assign n12509 = ( ~x2 & n12501 ) | ( ~x2 & n12507 ) | ( n12501 & n12507 ) ;
  assign n12510 = ( ~n12502 & n12508 ) | ( ~n12502 & n12509 ) | ( n12508 & n12509 ) ;
  assign n12511 = ( n12498 & n12500 ) | ( n12498 & n12510 ) | ( n12500 & n12510 ) ;
  assign n12512 = ( n12241 & n12243 ) | ( n12241 & n12511 ) | ( n12243 & n12511 ) ;
  assign n12513 = ( ~n11705 & n11707 ) | ( ~n11705 & n11960 ) | ( n11707 & n11960 ) ;
  assign n12514 = ( n11705 & ~n11961 ) | ( n11705 & n12513 ) | ( ~n11961 & n12513 ) ;
  assign n12515 = n9592 & ~n11676 ;
  assign n12516 = n9593 & n10245 ;
  assign n12517 = n41 & ~n10316 ;
  assign n12518 = n12516 | n12517 ;
  assign n12519 = x2 | n12518 ;
  assign n12520 = ( ~n12515 & n12518 ) | ( ~n12515 & n12519 ) | ( n12518 & n12519 ) ;
  assign n12521 = n9591 & ~n11676 ;
  assign n12522 = n12520 | n12521 ;
  assign n12523 = n9600 & n10247 ;
  assign n12524 = ( x2 & n12518 ) | ( x2 & n12523 ) | ( n12518 & n12523 ) ;
  assign n12525 = n12522 & ~n12524 ;
  assign n12526 = ( n12512 & n12514 ) | ( n12512 & n12525 ) | ( n12514 & n12525 ) ;
  assign n12527 = ( ~n11961 & n11971 ) | ( ~n11961 & n11973 ) | ( n11971 & n11973 ) ;
  assign n12528 = ( n11961 & ~n11974 ) | ( n11961 & n12527 ) | ( ~n11974 & n12527 ) ;
  assign n12529 = n9593 & ~n10320 ;
  assign n12530 = x2 & n12529 ;
  assign n12531 = n41 & n10245 ;
  assign n12532 = n9600 & ~n10316 ;
  assign n12533 = n12531 | n12532 ;
  assign n12534 = n9592 | n12533 ;
  assign n12535 = ( ~n10414 & n12533 ) | ( ~n10414 & n12534 ) | ( n12533 & n12534 ) ;
  assign n12536 = x2 & ~n12535 ;
  assign n12537 = ( ~x2 & n12529 ) | ( ~x2 & n12535 ) | ( n12529 & n12535 ) ;
  assign n12538 = ( ~n12530 & n12536 ) | ( ~n12530 & n12537 ) | ( n12536 & n12537 ) ;
  assign n12539 = ( n12526 & n12528 ) | ( n12526 & n12538 ) | ( n12528 & n12538 ) ;
  assign n12540 = n9592 & ~n11989 ;
  assign n12541 = n9593 & n10243 ;
  assign n12542 = n41 & ~n10320 ;
  assign n12543 = n12541 | n12542 ;
  assign n12544 = x2 | n12543 ;
  assign n12545 = ( ~n12540 & n12543 ) | ( ~n12540 & n12544 ) | ( n12543 & n12544 ) ;
  assign n12546 = n9591 & ~n11989 ;
  assign n12547 = n12545 | n12546 ;
  assign n12548 = n9600 & n10245 ;
  assign n12549 = ( x2 & n12543 ) | ( x2 & n12548 ) | ( n12543 & n12548 ) ;
  assign n12550 = n12547 & ~n12549 ;
  assign n12551 = ( ~n11695 & n11974 ) | ( ~n11695 & n11976 ) | ( n11974 & n11976 ) ;
  assign n12552 = ( n11695 & ~n11977 ) | ( n11695 & n12551 ) | ( ~n11977 & n12551 ) ;
  assign n12553 = ( n12539 & n12550 ) | ( n12539 & n12552 ) | ( n12550 & n12552 ) ;
  assign n12554 = n9592 & n12105 ;
  assign n12555 = n9593 & n10241 ;
  assign n12556 = n41 & n10243 ;
  assign n12557 = n12555 | n12556 ;
  assign n12558 = x2 | n12557 ;
  assign n12559 = ( ~n12554 & n12557 ) | ( ~n12554 & n12558 ) | ( n12557 & n12558 ) ;
  assign n12560 = n9591 & n12105 ;
  assign n12561 = n12559 | n12560 ;
  assign n12562 = n9600 & ~n10320 ;
  assign n12563 = ( x2 & n12557 ) | ( x2 & n12562 ) | ( n12557 & n12562 ) ;
  assign n12564 = n12561 & ~n12563 ;
  assign n12565 = ( ~n11680 & n11682 ) | ( ~n11680 & n11977 ) | ( n11682 & n11977 ) ;
  assign n12566 = ( n11680 & ~n11978 ) | ( n11680 & n12565 ) | ( ~n11978 & n12565 ) ;
  assign n12567 = ( n12553 & n12564 ) | ( n12553 & n12566 ) | ( n12564 & n12566 ) ;
  assign n12568 = ( ~n10422 & n11666 ) | ( ~n10422 & n11978 ) | ( n11666 & n11978 ) ;
  assign n12569 = ( n10422 & ~n11979 ) | ( n10422 & n12568 ) | ( ~n11979 & n12568 ) ;
  assign n12570 = n41 & n10241 ;
  assign n12571 = x2 & n12570 ;
  assign n12572 = n10239 & ~n10361 ;
  assign n12573 = ( n10239 & ~n10323 ) | ( n10239 & n10361 ) | ( ~n10323 & n10361 ) ;
  assign n12574 = n10239 & ~n10323 ;
  assign n12575 = ( n12572 & n12573 ) | ( n12572 & ~n12574 ) | ( n12573 & ~n12574 ) ;
  assign n12576 = n9600 & n10243 ;
  assign n12577 = n9593 | n12576 ;
  assign n12578 = ( n10239 & n12576 ) | ( n10239 & n12577 ) | ( n12576 & n12577 ) ;
  assign n12579 = n9592 | n12578 ;
  assign n12580 = ( n12575 & n12578 ) | ( n12575 & n12579 ) | ( n12578 & n12579 ) ;
  assign n12581 = x2 & ~n12580 ;
  assign n12582 = ( ~x2 & n12570 ) | ( ~x2 & n12580 ) | ( n12570 & n12580 ) ;
  assign n12583 = ( ~n12571 & n12581 ) | ( ~n12571 & n12582 ) | ( n12581 & n12582 ) ;
  assign n12584 = ( n12567 & n12569 ) | ( n12567 & n12583 ) | ( n12569 & n12583 ) ;
  assign n12585 = ( ~n11979 & n11993 ) | ( ~n11979 & n12095 ) | ( n11993 & n12095 ) ;
  assign n12586 = ( n11979 & ~n12096 ) | ( n11979 & n12585 ) | ( ~n12096 & n12585 ) ;
  assign n12587 = ( n12232 & n12584 ) | ( n12232 & n12586 ) | ( n12584 & n12586 ) ;
  assign n12588 = ( n10408 & n12219 ) | ( n10408 & n12587 ) | ( n12219 & n12587 ) ;
  assign n12589 = n40 & n10239 ;
  assign n12590 = n8721 & n10241 ;
  assign n12591 = n8340 & n10243 ;
  assign n12592 = n12590 | n12591 ;
  assign n12593 = n12589 | n12592 ;
  assign n12594 = x5 & n12593 ;
  assign n12595 = n8341 & n12575 ;
  assign n12596 = ( ~x5 & n12593 ) | ( ~x5 & n12595 ) | ( n12593 & n12595 ) ;
  assign n12597 = x5 & ~n12595 ;
  assign n12598 = ( ~n12594 & n12596 ) | ( ~n12594 & n12597 ) | ( n12596 & n12597 ) ;
  assign n12599 = n6571 & n10428 ;
  assign n12600 = x11 & n12599 ;
  assign n12601 = n6567 & ~n10249 ;
  assign n12602 = n6570 | n12601 ;
  assign n12603 = ( n10247 & n12601 ) | ( n10247 & n12602 ) | ( n12601 & n12602 ) ;
  assign n12604 = n6796 & n10312 ;
  assign n12605 = n12603 | n12604 ;
  assign n12606 = x11 & ~n12605 ;
  assign n12607 = ( ~x11 & n12599 ) | ( ~x11 & n12605 ) | ( n12599 & n12605 ) ;
  assign n12608 = ( ~n12600 & n12606 ) | ( ~n12600 & n12607 ) | ( n12606 & n12607 ) ;
  assign n12609 = n5915 & ~n11309 ;
  assign n12610 = x14 & n12609 ;
  assign n12611 = n5909 & n10255 ;
  assign n12612 = n5914 | n12611 ;
  assign n12613 = ( n10251 & n12611 ) | ( n10251 & n12612 ) | ( n12611 & n12612 ) ;
  assign n12614 = n6332 & ~n10253 ;
  assign n12615 = n12613 | n12614 ;
  assign n12616 = x14 & ~n12615 ;
  assign n12617 = ( ~x14 & n12609 ) | ( ~x14 & n12615 ) | ( n12609 & n12615 ) ;
  assign n12618 = ( ~n12610 & n12616 ) | ( ~n12610 & n12617 ) | ( n12616 & n12617 ) ;
  assign n12619 = n5232 & n10265 ;
  assign n12620 = x20 & n12619 ;
  assign n12621 = n4874 & n10267 ;
  assign n12622 = n4878 | n12621 ;
  assign n12623 = ( n10263 & n12621 ) | ( n10263 & n12622 ) | ( n12621 & n12622 ) ;
  assign n12624 = n4879 | n12623 ;
  assign n12625 = ( n10874 & n12623 ) | ( n10874 & n12624 ) | ( n12623 & n12624 ) ;
  assign n12626 = x20 & ~n12625 ;
  assign n12627 = ( ~x20 & n12619 ) | ( ~x20 & n12625 ) | ( n12619 & n12625 ) ;
  assign n12628 = ( ~n12620 & n12626 ) | ( ~n12620 & n12627 ) | ( n12626 & n12627 ) ;
  assign n12629 = n4649 & ~n10269 ;
  assign n12630 = n4591 | n12629 ;
  assign n12631 = ( ~n10698 & n12629 ) | ( ~n10698 & n12630 ) | ( n12629 & n12630 ) ;
  assign n12632 = n4584 & ~n10297 ;
  assign n12633 = ( ~x23 & n12631 ) | ( ~x23 & n12632 ) | ( n12631 & n12632 ) ;
  assign n12634 = n4637 & n10271 ;
  assign n12635 = x23 & ~n12632 ;
  assign n12636 = n12634 | n12635 ;
  assign n12637 = ( n12631 & n12634 ) | ( n12631 & n12635 ) | ( n12634 & n12635 ) ;
  assign n12638 = ( n12633 & n12636 ) | ( n12633 & ~n12637 ) | ( n12636 & ~n12637 ) ;
  assign n12639 = n4215 & n10273 ;
  assign n12640 = n4200 & n10275 ;
  assign n12641 = n2083 & n10277 ;
  assign n12642 = n12640 | n12641 ;
  assign n12643 = n12639 | n12642 ;
  assign n12644 = x26 & n12643 ;
  assign n12645 = n4203 & n10577 ;
  assign n12646 = ( ~x26 & n12643 ) | ( ~x26 & n12645 ) | ( n12643 & n12645 ) ;
  assign n12647 = x26 & ~n12645 ;
  assign n12648 = ( ~n12644 & n12646 ) | ( ~n12644 & n12647 ) | ( n12646 & n12647 ) ;
  assign n12649 = n4039 & n10291 ;
  assign n12650 = x29 & n12649 ;
  assign n12651 = n3501 & ~n10279 ;
  assign n12652 = n3536 & n10281 ;
  assign n12653 = n12651 | n12652 ;
  assign n12654 = n3541 | n12653 ;
  assign n12655 = ( n10454 & n12653 ) | ( n10454 & n12654 ) | ( n12653 & n12654 ) ;
  assign n12656 = x29 & ~n12655 ;
  assign n12657 = ( ~x29 & n12649 ) | ( ~x29 & n12655 ) | ( n12649 & n12655 ) ;
  assign n12658 = ( ~n12650 & n12656 ) | ( ~n12650 & n12657 ) | ( n12656 & n12657 ) ;
  assign n12659 = ~n390 & n10283 ;
  assign n12660 = n3270 | n10283 ;
  assign n12661 = ( n3274 & ~n12659 ) | ( n3274 & n12660 ) | ( ~n12659 & n12660 ) ;
  assign n12662 = ~n10285 & n12661 ;
  assign n12663 = n389 & n10286 ;
  assign n12664 = n12662 | n12663 ;
  assign n12665 = n97 | n140 ;
  assign n12666 = n756 | n1593 ;
  assign n12667 = n12665 | n12666 ;
  assign n12668 = n74 | n192 ;
  assign n12669 = n12667 | n12668 ;
  assign n12670 = n762 | n1392 ;
  assign n12671 = n831 | n12670 ;
  assign n12672 = n12669 | n12671 ;
  assign n12673 = n206 | n623 ;
  assign n12674 = n5427 | n12673 ;
  assign n12675 = n12672 | n12674 ;
  assign n12676 = n392 | n431 ;
  assign n12677 = n317 | n12676 ;
  assign n12678 = n2670 | n12677 ;
  assign n12679 = n174 | n370 ;
  assign n12680 = n12678 | n12679 ;
  assign n12681 = n1704 | n12680 ;
  assign n12682 = n605 | n1951 ;
  assign n12683 = n3434 | n12682 ;
  assign n12684 = n3348 | n12683 ;
  assign n12685 = n12681 | n12684 ;
  assign n12686 = n12675 | n12685 ;
  assign n12687 = n491 | n2598 ;
  assign n12688 = n2613 | n12687 ;
  assign n12689 = n345 | n751 ;
  assign n12690 = n700 | n12689 ;
  assign n12691 = n2762 | n12690 ;
  assign n12692 = n233 | n494 ;
  assign n12693 = n2107 | n12692 ;
  assign n12694 = n1977 | n12693 ;
  assign n12695 = n12691 | n12694 ;
  assign n12696 = n2538 | n12695 ;
  assign n12697 = n12688 | n12696 ;
  assign n12698 = n5942 | n12697 ;
  assign n12699 = n12686 | n12698 ;
  assign n12700 = n2848 & ~n12699 ;
  assign n12701 = ~n12664 & n12700 ;
  assign n12702 = n12664 & ~n12700 ;
  assign n12703 = n12701 | n12702 ;
  assign n12704 = n12179 & n12183 ;
  assign n12705 = ( n12658 & ~n12703 ) | ( n12658 & n12704 ) | ( ~n12703 & n12704 ) ;
  assign n12706 = ( n12658 & n12703 ) | ( n12658 & ~n12704 ) | ( n12703 & ~n12704 ) ;
  assign n12707 = ( ~n12658 & n12705 ) | ( ~n12658 & n12706 ) | ( n12705 & n12706 ) ;
  assign n12708 = ( n12197 & n12648 ) | ( n12197 & ~n12707 ) | ( n12648 & ~n12707 ) ;
  assign n12709 = ( n12197 & ~n12648 ) | ( n12197 & n12707 ) | ( ~n12648 & n12707 ) ;
  assign n12710 = ( ~n12197 & n12708 ) | ( ~n12197 & n12709 ) | ( n12708 & n12709 ) ;
  assign n12711 = ( n12200 & n12638 ) | ( n12200 & ~n12710 ) | ( n12638 & ~n12710 ) ;
  assign n12712 = ( n12200 & ~n12638 ) | ( n12200 & n12710 ) | ( ~n12638 & n12710 ) ;
  assign n12713 = ( ~n12200 & n12711 ) | ( ~n12200 & n12712 ) | ( n12711 & n12712 ) ;
  assign n12714 = ( n12203 & ~n12628 ) | ( n12203 & n12713 ) | ( ~n12628 & n12713 ) ;
  assign n12715 = ( n12203 & n12628 ) | ( n12203 & ~n12713 ) | ( n12628 & ~n12713 ) ;
  assign n12716 = ( ~n12203 & n12714 ) | ( ~n12203 & n12715 ) | ( n12714 & n12715 ) ;
  assign n12717 = n5584 & n10259 ;
  assign n12718 = x17 & n12717 ;
  assign n12719 = n5413 & n10261 ;
  assign n12720 = n5417 | n12719 ;
  assign n12721 = ( n10257 & n12719 ) | ( n10257 & n12720 ) | ( n12719 & n12720 ) ;
  assign n12722 = n5418 | n12721 ;
  assign n12723 = ( n11065 & n12721 ) | ( n11065 & n12722 ) | ( n12721 & n12722 ) ;
  assign n12724 = x17 & ~n12723 ;
  assign n12725 = ( ~x17 & n12717 ) | ( ~x17 & n12723 ) | ( n12717 & n12723 ) ;
  assign n12726 = ( ~n12718 & n12724 ) | ( ~n12718 & n12725 ) | ( n12724 & n12725 ) ;
  assign n12727 = ( n12206 & ~n12716 ) | ( n12206 & n12726 ) | ( ~n12716 & n12726 ) ;
  assign n12728 = ( n12206 & n12716 ) | ( n12206 & ~n12726 ) | ( n12716 & ~n12726 ) ;
  assign n12729 = ( ~n12206 & n12727 ) | ( ~n12206 & n12728 ) | ( n12727 & n12728 ) ;
  assign n12730 = ( n12209 & ~n12618 ) | ( n12209 & n12729 ) | ( ~n12618 & n12729 ) ;
  assign n12731 = ( n12209 & n12618 ) | ( n12209 & ~n12729 ) | ( n12618 & ~n12729 ) ;
  assign n12732 = ( ~n12209 & n12730 ) | ( ~n12209 & n12731 ) | ( n12730 & n12731 ) ;
  assign n12733 = ( n12212 & ~n12608 ) | ( n12212 & n12732 ) | ( ~n12608 & n12732 ) ;
  assign n12734 = ( n12212 & n12608 ) | ( n12212 & ~n12732 ) | ( n12608 & ~n12732 ) ;
  assign n12735 = ( ~n12212 & n12733 ) | ( ~n12212 & n12734 ) | ( n12733 & n12734 ) ;
  assign n12736 = n7345 & ~n10320 ;
  assign n12737 = n7644 & n10245 ;
  assign n12738 = n7341 & ~n10316 ;
  assign n12739 = n12737 | n12738 ;
  assign n12740 = n12736 | n12739 ;
  assign n12741 = x8 & n12740 ;
  assign n12742 = n7346 & ~n10414 ;
  assign n12743 = x8 & ~n12742 ;
  assign n12744 = ( ~x8 & n12740 ) | ( ~x8 & n12742 ) | ( n12740 & n12742 ) ;
  assign n12745 = ( ~n12741 & n12743 ) | ( ~n12741 & n12744 ) | ( n12743 & n12744 ) ;
  assign n12746 = ( n12215 & ~n12735 ) | ( n12215 & n12745 ) | ( ~n12735 & n12745 ) ;
  assign n12747 = ( n12215 & n12735 ) | ( n12215 & ~n12745 ) | ( n12735 & ~n12745 ) ;
  assign n12748 = ( ~n12215 & n12746 ) | ( ~n12215 & n12747 ) | ( n12746 & n12747 ) ;
  assign n12749 = ( n12218 & n12598 ) | ( n12218 & ~n12748 ) | ( n12598 & ~n12748 ) ;
  assign n12750 = ( ~n12218 & n12598 ) | ( ~n12218 & n12748 ) | ( n12598 & n12748 ) ;
  assign n12751 = ( ~n12598 & n12749 ) | ( ~n12598 & n12750 ) | ( n12749 & n12750 ) ;
  assign n12752 = ( n10394 & n12588 ) | ( n10394 & ~n12751 ) | ( n12588 & ~n12751 ) ;
  assign n12753 = ( n10237 & n10333 ) | ( n10237 & n10365 ) | ( n10333 & n10365 ) ;
  assign n12754 = n10237 | n10333 ;
  assign n12755 = ( ~n10237 & n10333 ) | ( ~n10237 & n10365 ) | ( n10333 & n10365 ) ;
  assign n12756 = ( ~n12753 & n12754 ) | ( ~n12753 & n12755 ) | ( n12754 & n12755 ) ;
  assign n12757 = n9592 & n12756 ;
  assign n12758 = x2 & n12757 ;
  assign n12759 = n9593 & ~n10237 ;
  assign n12760 = n41 & ~n10332 ;
  assign n12761 = n9600 & n10329 ;
  assign n12762 = n12760 | n12761 ;
  assign n12763 = n12759 | n12762 ;
  assign n12764 = x2 & ~n12763 ;
  assign n12765 = ( ~x2 & n12757 ) | ( ~x2 & n12763 ) | ( n12757 & n12763 ) ;
  assign n12766 = ( ~n12758 & n12764 ) | ( ~n12758 & n12765 ) | ( n12764 & n12765 ) ;
  assign n12767 = n40 & n10326 ;
  assign n12768 = n8721 & n10239 ;
  assign n12769 = n8340 & n10241 ;
  assign n12770 = n12768 | n12769 ;
  assign n12771 = n12767 | n12770 ;
  assign n12772 = x5 & n12771 ;
  assign n12773 = n8341 & n12222 ;
  assign n12774 = ( ~x5 & n12771 ) | ( ~x5 & n12773 ) | ( n12771 & n12773 ) ;
  assign n12775 = x5 & ~n12773 ;
  assign n12776 = ( ~n12772 & n12774 ) | ( ~n12772 & n12775 ) | ( n12774 & n12775 ) ;
  assign n12777 = n6571 & ~n11691 ;
  assign n12778 = x11 & n12777 ;
  assign n12779 = n6567 & n10312 ;
  assign n12780 = n6570 | n12779 ;
  assign n12781 = ( ~n10316 & n12779 ) | ( ~n10316 & n12780 ) | ( n12779 & n12780 ) ;
  assign n12782 = n6796 & n10247 ;
  assign n12783 = n12781 | n12782 ;
  assign n12784 = x11 & ~n12783 ;
  assign n12785 = ( ~x11 & n12777 ) | ( ~x11 & n12783 ) | ( n12777 & n12783 ) ;
  assign n12786 = ( ~n12778 & n12784 ) | ( ~n12778 & n12785 ) | ( n12784 & n12785 ) ;
  assign n12787 = n5584 & n10257 ;
  assign n12788 = x17 & n12787 ;
  assign n12789 = n5413 & n10259 ;
  assign n12790 = n5417 | n12789 ;
  assign n12791 = ( n10255 & n12789 ) | ( n10255 & n12790 ) | ( n12789 & n12790 ) ;
  assign n12792 = n5418 | n12791 ;
  assign n12793 = ( n11148 & n12791 ) | ( n11148 & n12792 ) | ( n12791 & n12792 ) ;
  assign n12794 = x17 & ~n12793 ;
  assign n12795 = ( ~x17 & n12787 ) | ( ~x17 & n12793 ) | ( n12787 & n12793 ) ;
  assign n12796 = ( ~n12788 & n12794 ) | ( ~n12788 & n12795 ) | ( n12794 & n12795 ) ;
  assign n12797 = n5232 & n10263 ;
  assign n12798 = x20 & n12797 ;
  assign n12799 = n4874 & n10265 ;
  assign n12800 = n4878 | n12799 ;
  assign n12801 = ( n10261 & n12799 ) | ( n10261 & n12800 ) | ( n12799 & n12800 ) ;
  assign n12802 = n4879 | n12801 ;
  assign n12803 = ( n11049 & n12801 ) | ( n11049 & n12802 ) | ( n12801 & n12802 ) ;
  assign n12804 = x20 & ~n12803 ;
  assign n12805 = ( ~x20 & n12797 ) | ( ~x20 & n12803 ) | ( n12797 & n12803 ) ;
  assign n12806 = ( ~n12798 & n12804 ) | ( ~n12798 & n12805 ) | ( n12804 & n12805 ) ;
  assign n12807 = n4591 & ~n10787 ;
  assign n12808 = x23 & n12807 ;
  assign n12809 = n4584 & n10271 ;
  assign n12810 = n4649 | n12809 ;
  assign n12811 = ( n10267 & n12809 ) | ( n10267 & n12810 ) | ( n12809 & n12810 ) ;
  assign n12812 = n4637 & ~n10269 ;
  assign n12813 = n12811 | n12812 ;
  assign n12814 = x23 & ~n12813 ;
  assign n12815 = ( ~x23 & n12807 ) | ( ~x23 & n12813 ) | ( n12807 & n12813 ) ;
  assign n12816 = ( ~n12808 & n12814 ) | ( ~n12808 & n12815 ) | ( n12814 & n12815 ) ;
  assign n12817 = n4215 & ~n10297 ;
  assign n12818 = n4200 & n10273 ;
  assign n12819 = n2083 & n10275 ;
  assign n12820 = n12818 | n12819 ;
  assign n12821 = n12817 | n12820 ;
  assign n12822 = x26 & n12821 ;
  assign n12823 = n4203 & ~n10617 ;
  assign n12824 = ( ~x26 & n12821 ) | ( ~x26 & n12823 ) | ( n12821 & n12823 ) ;
  assign n12825 = x26 & ~n12823 ;
  assign n12826 = ( ~n12822 & n12824 ) | ( ~n12822 & n12825 ) | ( n12824 & n12825 ) ;
  assign n12827 = n3501 & n10291 ;
  assign n12828 = x29 & n12827 ;
  assign n12829 = n3536 & ~n10279 ;
  assign n12830 = n4039 | n12829 ;
  assign n12831 = ( n10277 & n12829 ) | ( n10277 & n12830 ) | ( n12829 & n12830 ) ;
  assign n12832 = n3541 | n12831 ;
  assign n12833 = ( ~n10516 & n12831 ) | ( ~n10516 & n12832 ) | ( n12831 & n12832 ) ;
  assign n12834 = x29 & ~n12833 ;
  assign n12835 = ( ~x29 & n12827 ) | ( ~x29 & n12833 ) | ( n12827 & n12833 ) ;
  assign n12836 = ( ~n12828 & n12834 ) | ( ~n12828 & n12835 ) | ( n12834 & n12835 ) ;
  assign n12837 = n314 | n1094 ;
  assign n12838 = n777 | n864 ;
  assign n12839 = n2019 | n12838 ;
  assign n12840 = n12837 | n12839 ;
  assign n12841 = n2463 & ~n12840 ;
  assign n12842 = n534 | n712 ;
  assign n12843 = n2657 | n12842 ;
  assign n12844 = n220 | n405 ;
  assign n12845 = n308 | n378 ;
  assign n12846 = n12844 | n12845 ;
  assign n12847 = n917 | n12846 ;
  assign n12848 = n12682 | n12847 ;
  assign n12849 = n12843 | n12848 ;
  assign n12850 = n12841 & ~n12849 ;
  assign n12851 = n244 | n1041 ;
  assign n12852 = n3385 | n12851 ;
  assign n12853 = n727 | n12852 ;
  assign n12854 = n63 | n786 ;
  assign n12855 = n2603 | n12854 ;
  assign n12856 = n12853 | n12855 ;
  assign n12857 = n12850 & ~n12856 ;
  assign n12858 = n1876 | n12692 ;
  assign n12859 = n1003 | n12858 ;
  assign n12860 = n4952 | n12859 ;
  assign n12861 = n1957 | n2410 ;
  assign n12862 = n12860 | n12861 ;
  assign n12863 = n164 | n323 ;
  assign n12864 = n647 | n12863 ;
  assign n12865 = n6093 | n12864 ;
  assign n12866 = n679 | n700 ;
  assign n12867 = n634 | n12866 ;
  assign n12868 = n12865 | n12867 ;
  assign n12869 = n3337 | n12868 ;
  assign n12870 = n567 | n915 ;
  assign n12871 = n570 | n12870 ;
  assign n12872 = n163 | n265 ;
  assign n12873 = n391 | n12872 ;
  assign n12874 = n12871 | n12873 ;
  assign n12875 = n12869 | n12874 ;
  assign n12876 = n12862 | n12875 ;
  assign n12877 = n144 | n1332 ;
  assign n12878 = n357 | n2087 ;
  assign n12879 = n12877 | n12878 ;
  assign n12880 = n517 | n968 ;
  assign n12881 = n12879 | n12880 ;
  assign n12882 = n454 | n600 ;
  assign n12883 = n12881 | n12882 ;
  assign n12884 = n1407 | n1593 ;
  assign n12885 = n12883 | n12884 ;
  assign n12886 = n1688 | n1977 ;
  assign n12887 = n1519 | n12886 ;
  assign n12888 = n12885 | n12887 ;
  assign n12889 = n12876 | n12888 ;
  assign n12890 = n12857 & ~n12889 ;
  assign n12891 = n3273 & ~n10285 ;
  assign n12892 = n3270 | n12891 ;
  assign n12893 = ( n10281 & n12891 ) | ( n10281 & n12892 ) | ( n12891 & n12892 ) ;
  assign n12894 = n390 | n12893 ;
  assign n12895 = ( n10464 & n12893 ) | ( n10464 & n12894 ) | ( n12893 & n12894 ) ;
  assign n12896 = n3274 & ~n10283 ;
  assign n12897 = n12895 | n12896 ;
  assign n12898 = ( n12702 & ~n12890 ) | ( n12702 & n12897 ) | ( ~n12890 & n12897 ) ;
  assign n12899 = ( n12702 & n12890 ) | ( n12702 & ~n12897 ) | ( n12890 & ~n12897 ) ;
  assign n12900 = ( ~n12702 & n12898 ) | ( ~n12702 & n12899 ) | ( n12898 & n12899 ) ;
  assign n12901 = ( n12705 & n12836 ) | ( n12705 & ~n12900 ) | ( n12836 & ~n12900 ) ;
  assign n12902 = ( n12705 & ~n12836 ) | ( n12705 & n12900 ) | ( ~n12836 & n12900 ) ;
  assign n12903 = ( ~n12705 & n12901 ) | ( ~n12705 & n12902 ) | ( n12901 & n12902 ) ;
  assign n12904 = ( n12708 & n12826 ) | ( n12708 & ~n12903 ) | ( n12826 & ~n12903 ) ;
  assign n12905 = ( n12708 & ~n12826 ) | ( n12708 & n12903 ) | ( ~n12826 & n12903 ) ;
  assign n12906 = ( ~n12708 & n12904 ) | ( ~n12708 & n12905 ) | ( n12904 & n12905 ) ;
  assign n12907 = ( n12711 & n12816 ) | ( n12711 & ~n12906 ) | ( n12816 & ~n12906 ) ;
  assign n12908 = ( n12711 & ~n12816 ) | ( n12711 & n12906 ) | ( ~n12816 & n12906 ) ;
  assign n12909 = ( ~n12711 & n12907 ) | ( ~n12711 & n12908 ) | ( n12907 & n12908 ) ;
  assign n12910 = ( n12715 & n12806 ) | ( n12715 & ~n12909 ) | ( n12806 & ~n12909 ) ;
  assign n12911 = ( n12715 & ~n12806 ) | ( n12715 & n12909 ) | ( ~n12806 & n12909 ) ;
  assign n12912 = ( ~n12715 & n12910 ) | ( ~n12715 & n12911 ) | ( n12910 & n12911 ) ;
  assign n12913 = ( n12727 & n12796 ) | ( n12727 & ~n12912 ) | ( n12796 & ~n12912 ) ;
  assign n12914 = ( n12727 & ~n12796 ) | ( n12727 & n12912 ) | ( ~n12796 & n12912 ) ;
  assign n12915 = ( ~n12727 & n12913 ) | ( ~n12727 & n12914 ) | ( n12913 & n12914 ) ;
  assign n12916 = n6332 & n10251 ;
  assign n12917 = x14 & n12916 ;
  assign n12918 = n5909 & ~n10253 ;
  assign n12919 = n5914 | n12918 ;
  assign n12920 = ( ~n10249 & n12918 ) | ( ~n10249 & n12919 ) | ( n12918 & n12919 ) ;
  assign n12921 = n5915 | n12920 ;
  assign n12922 = ( ~n10441 & n12920 ) | ( ~n10441 & n12921 ) | ( n12920 & n12921 ) ;
  assign n12923 = x14 & ~n12922 ;
  assign n12924 = ( ~x14 & n12916 ) | ( ~x14 & n12922 ) | ( n12916 & n12922 ) ;
  assign n12925 = ( ~n12917 & n12923 ) | ( ~n12917 & n12924 ) | ( n12923 & n12924 ) ;
  assign n12926 = ( n12731 & n12915 ) | ( n12731 & n12925 ) | ( n12915 & n12925 ) ;
  assign n12927 = ( n12731 & ~n12915 ) | ( n12731 & n12925 ) | ( ~n12915 & n12925 ) ;
  assign n12928 = ( n12915 & ~n12926 ) | ( n12915 & n12927 ) | ( ~n12926 & n12927 ) ;
  assign n12929 = ( n12734 & n12786 ) | ( n12734 & ~n12928 ) | ( n12786 & ~n12928 ) ;
  assign n12930 = ( n12734 & ~n12786 ) | ( n12734 & n12928 ) | ( ~n12786 & n12928 ) ;
  assign n12931 = ( ~n12734 & n12929 ) | ( ~n12734 & n12930 ) | ( n12929 & n12930 ) ;
  assign n12932 = n7346 & ~n11989 ;
  assign n12933 = x8 & n12932 ;
  assign n12934 = n7345 & n10243 ;
  assign n12935 = n7644 & ~n10320 ;
  assign n12936 = n7341 & n10245 ;
  assign n12937 = n12935 | n12936 ;
  assign n12938 = n12934 | n12937 ;
  assign n12939 = x8 & ~n12938 ;
  assign n12940 = ( ~x8 & n12932 ) | ( ~x8 & n12938 ) | ( n12932 & n12938 ) ;
  assign n12941 = ( ~n12933 & n12939 ) | ( ~n12933 & n12940 ) | ( n12939 & n12940 ) ;
  assign n12942 = ( n12746 & n12931 ) | ( n12746 & n12941 ) | ( n12931 & n12941 ) ;
  assign n12943 = ( n12746 & ~n12931 ) | ( n12746 & n12941 ) | ( ~n12931 & n12941 ) ;
  assign n12944 = ( n12931 & ~n12942 ) | ( n12931 & n12943 ) | ( ~n12942 & n12943 ) ;
  assign n12945 = ( n12749 & n12776 ) | ( n12749 & ~n12944 ) | ( n12776 & ~n12944 ) ;
  assign n12946 = ( ~n12749 & n12776 ) | ( ~n12749 & n12944 ) | ( n12776 & n12944 ) ;
  assign n12947 = ( ~n12776 & n12945 ) | ( ~n12776 & n12946 ) | ( n12945 & n12946 ) ;
  assign n12948 = ( n12752 & n12766 ) | ( n12752 & ~n12947 ) | ( n12766 & ~n12947 ) ;
  assign n12949 = n41 & ~n10237 ;
  assign n12950 = x2 & n12949 ;
  assign n12951 = n10214 & ~n10366 ;
  assign n12952 = ( n10214 & ~n10334 ) | ( n10214 & n10366 ) | ( ~n10334 & n10366 ) ;
  assign n12953 = ( ~n10335 & n12951 ) | ( ~n10335 & n12952 ) | ( n12951 & n12952 ) ;
  assign n12954 = n9600 & ~n10332 ;
  assign n12955 = n9593 | n12954 ;
  assign n12956 = ( n10214 & n12954 ) | ( n10214 & n12955 ) | ( n12954 & n12955 ) ;
  assign n12957 = n9592 | n12956 ;
  assign n12958 = ( n12953 & n12956 ) | ( n12953 & n12957 ) | ( n12956 & n12957 ) ;
  assign n12959 = x2 & ~n12958 ;
  assign n12960 = ( ~x2 & n12949 ) | ( ~x2 & n12958 ) | ( n12949 & n12958 ) ;
  assign n12961 = ( ~n12950 & n12959 ) | ( ~n12950 & n12960 ) | ( n12959 & n12960 ) ;
  assign n12962 = n40 & n10329 ;
  assign n12963 = n8721 & n10326 ;
  assign n12964 = n8340 & n10239 ;
  assign n12965 = n12963 | n12964 ;
  assign n12966 = n12962 | n12965 ;
  assign n12967 = x5 & n12966 ;
  assign n12968 = n8341 & n10397 ;
  assign n12969 = ( ~x5 & n12966 ) | ( ~x5 & n12968 ) | ( n12966 & n12968 ) ;
  assign n12970 = x5 & ~n12968 ;
  assign n12971 = ( ~n12967 & n12969 ) | ( ~n12967 & n12970 ) | ( n12969 & n12970 ) ;
  assign n12972 = n7346 & n12105 ;
  assign n12973 = x8 & n12972 ;
  assign n12974 = n7341 & ~n10320 ;
  assign n12975 = n7345 | n12974 ;
  assign n12976 = ( n10241 & n12974 ) | ( n10241 & n12975 ) | ( n12974 & n12975 ) ;
  assign n12977 = n7644 & n10243 ;
  assign n12978 = n12976 | n12977 ;
  assign n12979 = x8 & ~n12978 ;
  assign n12980 = ( ~x8 & n12972 ) | ( ~x8 & n12978 ) | ( n12972 & n12978 ) ;
  assign n12981 = ( ~n12973 & n12979 ) | ( ~n12973 & n12980 ) | ( n12979 & n12980 ) ;
  assign n12982 = n6796 & ~n10316 ;
  assign n12983 = x11 & n12982 ;
  assign n12984 = n6567 & n10247 ;
  assign n12985 = n6570 | n12984 ;
  assign n12986 = ( n10245 & n12984 ) | ( n10245 & n12985 ) | ( n12984 & n12985 ) ;
  assign n12987 = n6571 | n12986 ;
  assign n12988 = ( ~n11676 & n12986 ) | ( ~n11676 & n12987 ) | ( n12986 & n12987 ) ;
  assign n12989 = x11 & ~n12988 ;
  assign n12990 = ( ~x11 & n12982 ) | ( ~x11 & n12988 ) | ( n12982 & n12988 ) ;
  assign n12991 = ( ~n12983 & n12989 ) | ( ~n12983 & n12990 ) | ( n12989 & n12990 ) ;
  assign n12992 = n5914 & n10312 ;
  assign n12993 = x14 & n12992 ;
  assign n12994 = n6332 & ~n10249 ;
  assign n12995 = n5909 & n10251 ;
  assign n12996 = n12994 | n12995 ;
  assign n12997 = n5915 | n12996 ;
  assign n12998 = ( ~n11486 & n12996 ) | ( ~n11486 & n12997 ) | ( n12996 & n12997 ) ;
  assign n12999 = x14 & ~n12998 ;
  assign n13000 = ( ~x14 & n12992 ) | ( ~x14 & n12998 ) | ( n12992 & n12998 ) ;
  assign n13001 = ( ~n12993 & n12999 ) | ( ~n12993 & n13000 ) | ( n12999 & n13000 ) ;
  assign n13002 = n5232 & n10261 ;
  assign n13003 = x20 & n13002 ;
  assign n13004 = n4874 & n10263 ;
  assign n13005 = n4878 | n13004 ;
  assign n13006 = ( n10259 & n13004 ) | ( n10259 & n13005 ) | ( n13004 & n13005 ) ;
  assign n13007 = n4879 | n13006 ;
  assign n13008 = ( n10859 & n13006 ) | ( n10859 & n13007 ) | ( n13006 & n13007 ) ;
  assign n13009 = x20 & ~n13008 ;
  assign n13010 = ( ~x20 & n13002 ) | ( ~x20 & n13008 ) | ( n13002 & n13008 ) ;
  assign n13011 = ( ~n13003 & n13009 ) | ( ~n13003 & n13010 ) | ( n13009 & n13010 ) ;
  assign n13012 = n4637 & n10267 ;
  assign n13013 = x23 & n13012 ;
  assign n13014 = n4584 & ~n10269 ;
  assign n13015 = n4649 | n13014 ;
  assign n13016 = ( n10265 & n13014 ) | ( n10265 & n13015 ) | ( n13014 & n13015 ) ;
  assign n13017 = n4591 | n13016 ;
  assign n13018 = ( n10804 & n13016 ) | ( n10804 & n13017 ) | ( n13016 & n13017 ) ;
  assign n13019 = x23 & ~n13018 ;
  assign n13020 = ( ~x23 & n13012 ) | ( ~x23 & n13018 ) | ( n13012 & n13018 ) ;
  assign n13021 = ( ~n13013 & n13019 ) | ( ~n13013 & n13020 ) | ( n13019 & n13020 ) ;
  assign n13022 = n4215 & n10271 ;
  assign n13023 = n4200 & ~n10297 ;
  assign n13024 = n2083 & n10273 ;
  assign n13025 = n13023 | n13024 ;
  assign n13026 = n13022 | n13025 ;
  assign n13027 = x26 & n13026 ;
  assign n13028 = n4203 & ~n10656 ;
  assign n13029 = ( ~x26 & n13026 ) | ( ~x26 & n13028 ) | ( n13026 & n13028 ) ;
  assign n13030 = x26 & ~n13028 ;
  assign n13031 = ( ~n13027 & n13029 ) | ( ~n13027 & n13030 ) | ( n13029 & n13030 ) ;
  assign n13032 = n3501 & n10277 ;
  assign n13033 = x29 & n13032 ;
  assign n13034 = n3536 & n10291 ;
  assign n13035 = n4039 | n13034 ;
  assign n13036 = ( n10275 & n13034 ) | ( n10275 & n13035 ) | ( n13034 & n13035 ) ;
  assign n13037 = n3541 | n13036 ;
  assign n13038 = ( n10563 & n13036 ) | ( n10563 & n13037 ) | ( n13036 & n13037 ) ;
  assign n13039 = x29 & ~n13038 ;
  assign n13040 = ( ~x29 & n13032 ) | ( ~x29 & n13038 ) | ( n13032 & n13038 ) ;
  assign n13041 = ( ~n13033 & n13039 ) | ( ~n13033 & n13040 ) | ( n13039 & n13040 ) ;
  assign n13042 = n454 | n554 ;
  assign n13043 = n656 | n13042 ;
  assign n13044 = n578 | n13043 ;
  assign n13045 = n6134 | n13044 ;
  assign n13046 = n1084 | n3970 ;
  assign n13047 = n265 | n334 ;
  assign n13048 = n13046 | n13047 ;
  assign n13049 = n13045 | n13048 ;
  assign n13050 = n10161 | n13049 ;
  assign n13051 = n3077 | n3441 ;
  assign n13052 = n5077 | n13051 ;
  assign n13053 = n13050 | n13052 ;
  assign n13054 = n3669 | n3950 ;
  assign n13055 = n13053 | n13054 ;
  assign n13056 = n3273 & ~n10283 ;
  assign n13057 = n3270 | n13056 ;
  assign n13058 = ( ~n10279 & n13056 ) | ( ~n10279 & n13057 ) | ( n13056 & n13057 ) ;
  assign n13059 = n390 | n13058 ;
  assign n13060 = ( n10487 & n13058 ) | ( n10487 & n13059 ) | ( n13058 & n13059 ) ;
  assign n13061 = n3274 & n10281 ;
  assign n13062 = n13060 | n13061 ;
  assign n13063 = ( n12898 & n13055 ) | ( n12898 & n13062 ) | ( n13055 & n13062 ) ;
  assign n13064 = ( ~n12898 & n13055 ) | ( ~n12898 & n13062 ) | ( n13055 & n13062 ) ;
  assign n13065 = ( n12898 & ~n13063 ) | ( n12898 & n13064 ) | ( ~n13063 & n13064 ) ;
  assign n13066 = ( ~n12901 & n13041 ) | ( ~n12901 & n13065 ) | ( n13041 & n13065 ) ;
  assign n13067 = ( n12901 & n13041 ) | ( n12901 & n13065 ) | ( n13041 & n13065 ) ;
  assign n13068 = ( n12901 & n13066 ) | ( n12901 & ~n13067 ) | ( n13066 & ~n13067 ) ;
  assign n13069 = ( ~n12904 & n13031 ) | ( ~n12904 & n13068 ) | ( n13031 & n13068 ) ;
  assign n13070 = ( n12904 & n13031 ) | ( n12904 & n13068 ) | ( n13031 & n13068 ) ;
  assign n13071 = ( n12904 & n13069 ) | ( n12904 & ~n13070 ) | ( n13069 & ~n13070 ) ;
  assign n13072 = ( ~n12907 & n13021 ) | ( ~n12907 & n13071 ) | ( n13021 & n13071 ) ;
  assign n13073 = ( n12907 & n13021 ) | ( n12907 & n13071 ) | ( n13021 & n13071 ) ;
  assign n13074 = ( n12907 & n13072 ) | ( n12907 & ~n13073 ) | ( n13072 & ~n13073 ) ;
  assign n13075 = ( ~n12910 & n13011 ) | ( ~n12910 & n13074 ) | ( n13011 & n13074 ) ;
  assign n13076 = ( n12910 & n13011 ) | ( n12910 & n13074 ) | ( n13011 & n13074 ) ;
  assign n13077 = ( n12910 & n13075 ) | ( n12910 & ~n13076 ) | ( n13075 & ~n13076 ) ;
  assign n13078 = n5418 & ~n11297 ;
  assign n13079 = x17 & n13078 ;
  assign n13080 = n5413 & n10257 ;
  assign n13081 = n5417 | n13080 ;
  assign n13082 = ( ~n10253 & n13080 ) | ( ~n10253 & n13081 ) | ( n13080 & n13081 ) ;
  assign n13083 = n5584 & n10255 ;
  assign n13084 = n13082 | n13083 ;
  assign n13085 = x17 & ~n13084 ;
  assign n13086 = ( ~x17 & n13078 ) | ( ~x17 & n13084 ) | ( n13078 & n13084 ) ;
  assign n13087 = ( ~n13079 & n13085 ) | ( ~n13079 & n13086 ) | ( n13085 & n13086 ) ;
  assign n13088 = ( ~n12913 & n13077 ) | ( ~n12913 & n13087 ) | ( n13077 & n13087 ) ;
  assign n13089 = ( n12913 & n13077 ) | ( n12913 & n13087 ) | ( n13077 & n13087 ) ;
  assign n13090 = ( n12913 & n13088 ) | ( n12913 & ~n13089 ) | ( n13088 & ~n13089 ) ;
  assign n13091 = ( ~n12927 & n13001 ) | ( ~n12927 & n13090 ) | ( n13001 & n13090 ) ;
  assign n13092 = ( n12927 & n13001 ) | ( n12927 & n13090 ) | ( n13001 & n13090 ) ;
  assign n13093 = ( n12927 & n13091 ) | ( n12927 & ~n13092 ) | ( n13091 & ~n13092 ) ;
  assign n13094 = ( ~n12929 & n12991 ) | ( ~n12929 & n13093 ) | ( n12991 & n13093 ) ;
  assign n13095 = ( n12929 & n12991 ) | ( n12929 & n13093 ) | ( n12991 & n13093 ) ;
  assign n13096 = ( n12929 & n13094 ) | ( n12929 & ~n13095 ) | ( n13094 & ~n13095 ) ;
  assign n13097 = ( n12943 & ~n12981 ) | ( n12943 & n13096 ) | ( ~n12981 & n13096 ) ;
  assign n13098 = ( n12943 & n12981 ) | ( n12943 & n13096 ) | ( n12981 & n13096 ) ;
  assign n13099 = ( n12981 & n13097 ) | ( n12981 & ~n13098 ) | ( n13097 & ~n13098 ) ;
  assign n13100 = ( ~n12945 & n12971 ) | ( ~n12945 & n13099 ) | ( n12971 & n13099 ) ;
  assign n13101 = ( n12945 & n12971 ) | ( n12945 & n13099 ) | ( n12971 & n13099 ) ;
  assign n13102 = ( n12945 & n13100 ) | ( n12945 & ~n13101 ) | ( n13100 & ~n13101 ) ;
  assign n13103 = ( n12948 & n12961 ) | ( n12948 & n13102 ) | ( n12961 & n13102 ) ;
  assign n13104 = n40 & ~n10332 ;
  assign n13105 = n8721 & n10329 ;
  assign n13106 = n8340 & n10326 ;
  assign n13107 = n13105 | n13106 ;
  assign n13108 = n13104 | n13107 ;
  assign n13109 = x5 & n13108 ;
  assign n13110 = n8341 & ~n10383 ;
  assign n13111 = ( ~x5 & n13108 ) | ( ~x5 & n13110 ) | ( n13108 & n13110 ) ;
  assign n13112 = x5 & ~n13110 ;
  assign n13113 = ( ~n13109 & n13111 ) | ( ~n13109 & n13112 ) | ( n13111 & n13112 ) ;
  assign n13114 = n7644 & n10241 ;
  assign n13115 = x8 & n13114 ;
  assign n13116 = n7341 & n10243 ;
  assign n13117 = n7345 | n13116 ;
  assign n13118 = ( n10239 & n13116 ) | ( n10239 & n13117 ) | ( n13116 & n13117 ) ;
  assign n13119 = n7346 | n13118 ;
  assign n13120 = ( n12575 & n13118 ) | ( n12575 & n13119 ) | ( n13118 & n13119 ) ;
  assign n13121 = x8 & ~n13120 ;
  assign n13122 = ( ~x8 & n13114 ) | ( ~x8 & n13120 ) | ( n13114 & n13120 ) ;
  assign n13123 = ( ~n13115 & n13121 ) | ( ~n13115 & n13122 ) | ( n13121 & n13122 ) ;
  assign n13124 = n6570 & ~n10320 ;
  assign n13125 = x11 & n13124 ;
  assign n13126 = n6796 & n10245 ;
  assign n13127 = n6567 & ~n10316 ;
  assign n13128 = n13126 | n13127 ;
  assign n13129 = n6571 | n13128 ;
  assign n13130 = ( ~n10414 & n13128 ) | ( ~n10414 & n13129 ) | ( n13128 & n13129 ) ;
  assign n13131 = x11 & ~n13130 ;
  assign n13132 = ( ~x11 & n13124 ) | ( ~x11 & n13130 ) | ( n13124 & n13130 ) ;
  assign n13133 = ( ~n13125 & n13131 ) | ( ~n13125 & n13132 ) | ( n13131 & n13132 ) ;
  assign n13134 = n5584 & ~n10253 ;
  assign n13135 = x17 & n13134 ;
  assign n13136 = n5413 & n10255 ;
  assign n13137 = n5417 | n13136 ;
  assign n13138 = ( n10251 & n13136 ) | ( n10251 & n13137 ) | ( n13136 & n13137 ) ;
  assign n13139 = n5418 | n13138 ;
  assign n13140 = ( ~n11309 & n13138 ) | ( ~n11309 & n13139 ) | ( n13138 & n13139 ) ;
  assign n13141 = x17 & ~n13140 ;
  assign n13142 = ( ~x17 & n13134 ) | ( ~x17 & n13140 ) | ( n13134 & n13140 ) ;
  assign n13143 = ( ~n13135 & n13141 ) | ( ~n13135 & n13142 ) | ( n13141 & n13142 ) ;
  assign n13144 = n5232 & n10259 ;
  assign n13145 = x20 & n13144 ;
  assign n13146 = n4874 & n10261 ;
  assign n13147 = n4878 | n13146 ;
  assign n13148 = ( n10257 & n13146 ) | ( n10257 & n13147 ) | ( n13146 & n13147 ) ;
  assign n13149 = n4879 | n13148 ;
  assign n13150 = ( n11065 & n13148 ) | ( n11065 & n13149 ) | ( n13148 & n13149 ) ;
  assign n13151 = x20 & ~n13150 ;
  assign n13152 = ( ~x20 & n13144 ) | ( ~x20 & n13150 ) | ( n13144 & n13150 ) ;
  assign n13153 = ( ~n13145 & n13151 ) | ( ~n13145 & n13152 ) | ( n13151 & n13152 ) ;
  assign n13154 = n4637 & n10265 ;
  assign n13155 = x23 & n13154 ;
  assign n13156 = n4584 & n10267 ;
  assign n13157 = n4649 | n13156 ;
  assign n13158 = ( n10263 & n13156 ) | ( n10263 & n13157 ) | ( n13156 & n13157 ) ;
  assign n13159 = n4591 | n13158 ;
  assign n13160 = ( n10874 & n13158 ) | ( n10874 & n13159 ) | ( n13158 & n13159 ) ;
  assign n13161 = x23 & ~n13160 ;
  assign n13162 = ( ~x23 & n13154 ) | ( ~x23 & n13160 ) | ( n13154 & n13160 ) ;
  assign n13163 = ( ~n13155 & n13161 ) | ( ~n13155 & n13162 ) | ( n13161 & n13162 ) ;
  assign n13164 = n4215 & ~n10269 ;
  assign n13165 = n4200 & n10271 ;
  assign n13166 = n2083 & ~n10297 ;
  assign n13167 = n13165 | n13166 ;
  assign n13168 = n13164 | n13167 ;
  assign n13169 = x26 & n13168 ;
  assign n13170 = n4203 & ~n10698 ;
  assign n13171 = ( ~x26 & n13168 ) | ( ~x26 & n13170 ) | ( n13168 & n13170 ) ;
  assign n13172 = x26 & ~n13170 ;
  assign n13173 = ( ~n13169 & n13171 ) | ( ~n13169 & n13172 ) | ( n13171 & n13172 ) ;
  assign n13174 = n3541 & n10577 ;
  assign n13175 = x29 & n13174 ;
  assign n13176 = n3536 & n10277 ;
  assign n13177 = n4039 | n13176 ;
  assign n13178 = ( n10273 & n13176 ) | ( n10273 & n13177 ) | ( n13176 & n13177 ) ;
  assign n13179 = n3501 & n10275 ;
  assign n13180 = n13178 | n13179 ;
  assign n13181 = x29 & ~n13180 ;
  assign n13182 = ( ~x29 & n13174 ) | ( ~x29 & n13180 ) | ( n13174 & n13180 ) ;
  assign n13183 = ( ~n13175 & n13181 ) | ( ~n13175 & n13182 ) | ( n13181 & n13182 ) ;
  assign n13184 = n3274 & ~n10279 ;
  assign n13185 = n3273 & n10281 ;
  assign n13186 = n13184 | n13185 ;
  assign n13187 = n390 | n13186 ;
  assign n13188 = ( n10454 & n13186 ) | ( n10454 & n13187 ) | ( n13186 & n13187 ) ;
  assign n13189 = n3270 & n10291 ;
  assign n13190 = n13188 | n13189 ;
  assign n13191 = n441 | n500 ;
  assign n13192 = n2214 | n13191 ;
  assign n13193 = n590 | n13192 ;
  assign n13194 = n611 | n1849 ;
  assign n13195 = n13193 | n13194 ;
  assign n13196 = n2770 | n13195 ;
  assign n13197 = n343 | n2666 ;
  assign n13198 = n1732 | n13197 ;
  assign n13199 = n4766 | n13198 ;
  assign n13200 = n1279 | n13199 ;
  assign n13201 = n13196 | n13200 ;
  assign n13202 = n283 | n13201 ;
  assign n13203 = n367 | n1727 ;
  assign n13204 = n2934 | n13203 ;
  assign n13205 = n1997 | n2636 ;
  assign n13206 = n13204 | n13205 ;
  assign n13207 = n337 | n794 ;
  assign n13208 = n151 | n13207 ;
  assign n13209 = n3905 | n13208 ;
  assign n13210 = n620 & ~n13209 ;
  assign n13211 = n428 | n3709 ;
  assign n13212 = n1007 | n13211 ;
  assign n13213 = n2851 | n13212 ;
  assign n13214 = n13210 & ~n13213 ;
  assign n13215 = ~n13206 & n13214 ;
  assign n13216 = n700 | n3519 ;
  assign n13217 = n123 | n290 ;
  assign n13218 = n13216 | n13217 ;
  assign n13219 = n667 | n751 ;
  assign n13220 = n987 | n13219 ;
  assign n13221 = n1415 | n13220 ;
  assign n13222 = n4101 | n13221 ;
  assign n13223 = n13218 | n13222 ;
  assign n13224 = n13215 & ~n13223 ;
  assign n13225 = ~n13202 & n13224 ;
  assign n13226 = ( n13063 & n13190 ) | ( n13063 & ~n13225 ) | ( n13190 & ~n13225 ) ;
  assign n13227 = ( ~n13063 & n13190 ) | ( ~n13063 & n13225 ) | ( n13190 & n13225 ) ;
  assign n13228 = ( ~n13190 & n13226 ) | ( ~n13190 & n13227 ) | ( n13226 & n13227 ) ;
  assign n13229 = ( n13067 & n13183 ) | ( n13067 & ~n13228 ) | ( n13183 & ~n13228 ) ;
  assign n13230 = ( n13067 & ~n13183 ) | ( n13067 & n13228 ) | ( ~n13183 & n13228 ) ;
  assign n13231 = ( ~n13067 & n13229 ) | ( ~n13067 & n13230 ) | ( n13229 & n13230 ) ;
  assign n13232 = ( n13070 & ~n13173 ) | ( n13070 & n13231 ) | ( ~n13173 & n13231 ) ;
  assign n13233 = ( n13070 & n13173 ) | ( n13070 & ~n13231 ) | ( n13173 & ~n13231 ) ;
  assign n13234 = ( ~n13070 & n13232 ) | ( ~n13070 & n13233 ) | ( n13232 & n13233 ) ;
  assign n13235 = ( n13073 & ~n13163 ) | ( n13073 & n13234 ) | ( ~n13163 & n13234 ) ;
  assign n13236 = ( n13073 & n13163 ) | ( n13073 & ~n13234 ) | ( n13163 & ~n13234 ) ;
  assign n13237 = ( ~n13073 & n13235 ) | ( ~n13073 & n13236 ) | ( n13235 & n13236 ) ;
  assign n13238 = ( n13076 & n13153 ) | ( n13076 & ~n13237 ) | ( n13153 & ~n13237 ) ;
  assign n13239 = ( n13076 & ~n13153 ) | ( n13076 & n13237 ) | ( ~n13153 & n13237 ) ;
  assign n13240 = ( ~n13076 & n13238 ) | ( ~n13076 & n13239 ) | ( n13238 & n13239 ) ;
  assign n13241 = ( n13089 & n13143 ) | ( n13089 & ~n13240 ) | ( n13143 & ~n13240 ) ;
  assign n13242 = ( n13089 & ~n13143 ) | ( n13089 & n13240 ) | ( ~n13143 & n13240 ) ;
  assign n13243 = ( ~n13089 & n13241 ) | ( ~n13089 & n13242 ) | ( n13241 & n13242 ) ;
  assign n13244 = n6332 & n10312 ;
  assign n13245 = x14 & n13244 ;
  assign n13246 = n5909 & ~n10249 ;
  assign n13247 = n5914 | n13246 ;
  assign n13248 = ( n10247 & n13246 ) | ( n10247 & n13247 ) | ( n13246 & n13247 ) ;
  assign n13249 = n5915 | n13248 ;
  assign n13250 = ( n10428 & n13248 ) | ( n10428 & n13249 ) | ( n13248 & n13249 ) ;
  assign n13251 = x14 & ~n13250 ;
  assign n13252 = ( ~x14 & n13244 ) | ( ~x14 & n13250 ) | ( n13244 & n13250 ) ;
  assign n13253 = ( ~n13245 & n13251 ) | ( ~n13245 & n13252 ) | ( n13251 & n13252 ) ;
  assign n13254 = ( n13092 & n13243 ) | ( n13092 & n13253 ) | ( n13243 & n13253 ) ;
  assign n13255 = ( n13092 & ~n13243 ) | ( n13092 & n13253 ) | ( ~n13243 & n13253 ) ;
  assign n13256 = ( n13243 & ~n13254 ) | ( n13243 & n13255 ) | ( ~n13254 & n13255 ) ;
  assign n13257 = ( n13095 & n13133 ) | ( n13095 & ~n13256 ) | ( n13133 & ~n13256 ) ;
  assign n13258 = ( n13095 & ~n13133 ) | ( n13095 & n13256 ) | ( ~n13133 & n13256 ) ;
  assign n13259 = ( ~n13095 & n13257 ) | ( ~n13095 & n13258 ) | ( n13257 & n13258 ) ;
  assign n13260 = ( n13098 & n13123 ) | ( n13098 & ~n13259 ) | ( n13123 & ~n13259 ) ;
  assign n13261 = ( n13098 & ~n13123 ) | ( n13098 & n13259 ) | ( ~n13123 & n13259 ) ;
  assign n13262 = ( ~n13098 & n13260 ) | ( ~n13098 & n13261 ) | ( n13260 & n13261 ) ;
  assign n13263 = ( n13101 & n13113 ) | ( n13101 & ~n13262 ) | ( n13113 & ~n13262 ) ;
  assign n13264 = ( n13101 & ~n13113 ) | ( n13101 & n13262 ) | ( ~n13113 & n13262 ) ;
  assign n13265 = ( ~n13101 & n13263 ) | ( ~n13101 & n13264 ) | ( n13263 & n13264 ) ;
  assign n13266 = ( n10379 & n13103 ) | ( n10379 & ~n13265 ) | ( n13103 & ~n13265 ) ;
  assign n13267 = n10235 & ~n10335 ;
  assign n13268 = n220 | n662 ;
  assign n13269 = n87 | n13268 ;
  assign n13270 = n1351 | n13269 ;
  assign n13271 = n3481 & ~n3512 ;
  assign n13272 = ~n13270 & n13271 ;
  assign n13273 = ~n10193 & n13272 ;
  assign n13274 = ~n3529 & n13273 ;
  assign n13275 = n10229 & ~n13274 ;
  assign n13276 = ~n10229 & n13274 ;
  assign n13277 = n13275 | n13276 ;
  assign n13278 = ( ~n10230 & n10234 ) | ( ~n10230 & n13277 ) | ( n10234 & n13277 ) ;
  assign n13279 = ( n10230 & n10234 ) | ( n10230 & n13277 ) | ( n10234 & n13277 ) ;
  assign n13280 = ( n10230 & n13278 ) | ( n10230 & ~n13279 ) | ( n13278 & ~n13279 ) ;
  assign n13281 = n13267 & n13280 ;
  assign n13282 = n10235 | n10367 ;
  assign n13283 = ( ~n13267 & n13280 ) | ( ~n13267 & n13282 ) | ( n13280 & n13282 ) ;
  assign n13284 = n13280 & n13282 ;
  assign n13285 = ( n13281 & n13283 ) | ( n13281 & ~n13284 ) | ( n13283 & ~n13284 ) ;
  assign n13286 = n9592 & ~n13285 ;
  assign n13287 = n9593 & ~n13280 ;
  assign n13288 = n41 & ~n10235 ;
  assign n13289 = n13287 | n13288 ;
  assign n13290 = x2 | n13289 ;
  assign n13291 = ( ~n13286 & n13289 ) | ( ~n13286 & n13290 ) | ( n13289 & n13290 ) ;
  assign n13292 = n9591 & ~n13285 ;
  assign n13293 = n13291 | n13292 ;
  assign n13294 = n9600 & n10214 ;
  assign n13295 = ( x2 & n13289 ) | ( x2 & n13294 ) | ( n13289 & n13294 ) ;
  assign n13296 = n13293 & ~n13295 ;
  assign n13297 = n40 & ~n10237 ;
  assign n13298 = n8721 & ~n10332 ;
  assign n13299 = n8340 & n10329 ;
  assign n13300 = n13298 | n13299 ;
  assign n13301 = n13297 | n13300 ;
  assign n13302 = x5 & n13301 ;
  assign n13303 = n8341 & n12756 ;
  assign n13304 = ( ~x5 & n13301 ) | ( ~x5 & n13303 ) | ( n13301 & n13303 ) ;
  assign n13305 = x5 & ~n13303 ;
  assign n13306 = ( ~n13302 & n13304 ) | ( ~n13302 & n13305 ) | ( n13304 & n13305 ) ;
  assign n13307 = n7644 & n10239 ;
  assign n13308 = x8 & n13307 ;
  assign n13309 = n7341 & n10241 ;
  assign n13310 = n7345 | n13309 ;
  assign n13311 = ( n10326 & n13309 ) | ( n10326 & n13310 ) | ( n13309 & n13310 ) ;
  assign n13312 = n7346 | n13311 ;
  assign n13313 = ( n12222 & n13311 ) | ( n12222 & n13312 ) | ( n13311 & n13312 ) ;
  assign n13314 = x8 & ~n13313 ;
  assign n13315 = ( ~x8 & n13307 ) | ( ~x8 & n13313 ) | ( n13307 & n13313 ) ;
  assign n13316 = ( ~n13308 & n13314 ) | ( ~n13308 & n13315 ) | ( n13314 & n13315 ) ;
  assign n13317 = n5915 & ~n11691 ;
  assign n13318 = x14 & n13317 ;
  assign n13319 = n5909 & n10312 ;
  assign n13320 = n5914 | n13319 ;
  assign n13321 = ( ~n10316 & n13319 ) | ( ~n10316 & n13320 ) | ( n13319 & n13320 ) ;
  assign n13322 = n6332 & n10247 ;
  assign n13323 = n13321 | n13322 ;
  assign n13324 = x14 & ~n13323 ;
  assign n13325 = ( ~x14 & n13317 ) | ( ~x14 & n13323 ) | ( n13317 & n13323 ) ;
  assign n13326 = ( ~n13318 & n13324 ) | ( ~n13318 & n13325 ) | ( n13324 & n13325 ) ;
  assign n13327 = n5584 & n10251 ;
  assign n13328 = x17 & n13327 ;
  assign n13329 = n5413 & ~n10253 ;
  assign n13330 = n5417 | n13329 ;
  assign n13331 = ( ~n10249 & n13329 ) | ( ~n10249 & n13330 ) | ( n13329 & n13330 ) ;
  assign n13332 = n5418 | n13331 ;
  assign n13333 = ( ~n10441 & n13331 ) | ( ~n10441 & n13332 ) | ( n13331 & n13332 ) ;
  assign n13334 = x17 & ~n13333 ;
  assign n13335 = ( ~x17 & n13327 ) | ( ~x17 & n13333 ) | ( n13327 & n13333 ) ;
  assign n13336 = ( ~n13328 & n13334 ) | ( ~n13328 & n13335 ) | ( n13334 & n13335 ) ;
  assign n13337 = n5232 & n10257 ;
  assign n13338 = x20 & n13337 ;
  assign n13339 = n4874 & n10259 ;
  assign n13340 = n4878 | n13339 ;
  assign n13341 = ( n10255 & n13339 ) | ( n10255 & n13340 ) | ( n13339 & n13340 ) ;
  assign n13342 = n4879 | n13341 ;
  assign n13343 = ( n11148 & n13341 ) | ( n11148 & n13342 ) | ( n13341 & n13342 ) ;
  assign n13344 = x20 & ~n13343 ;
  assign n13345 = ( ~x20 & n13337 ) | ( ~x20 & n13343 ) | ( n13337 & n13343 ) ;
  assign n13346 = ( ~n13338 & n13344 ) | ( ~n13338 & n13345 ) | ( n13344 & n13345 ) ;
  assign n13347 = n4637 & n10263 ;
  assign n13348 = x23 & n13347 ;
  assign n13349 = n4584 & n10265 ;
  assign n13350 = n4649 | n13349 ;
  assign n13351 = ( n10261 & n13349 ) | ( n10261 & n13350 ) | ( n13349 & n13350 ) ;
  assign n13352 = n4591 | n13351 ;
  assign n13353 = ( n11049 & n13351 ) | ( n11049 & n13352 ) | ( n13351 & n13352 ) ;
  assign n13354 = x23 & ~n13353 ;
  assign n13355 = ( ~x23 & n13347 ) | ( ~x23 & n13353 ) | ( n13347 & n13353 ) ;
  assign n13356 = ( ~n13348 & n13354 ) | ( ~n13348 & n13355 ) | ( n13354 & n13355 ) ;
  assign n13357 = n4215 & n10267 ;
  assign n13358 = n4200 & ~n10269 ;
  assign n13359 = n2083 & n10271 ;
  assign n13360 = n13358 | n13359 ;
  assign n13361 = n13357 | n13360 ;
  assign n13362 = x26 & n13361 ;
  assign n13363 = n4203 & ~n10787 ;
  assign n13364 = ( ~x26 & n13361 ) | ( ~x26 & n13363 ) | ( n13361 & n13363 ) ;
  assign n13365 = x26 & ~n13363 ;
  assign n13366 = ( ~n13362 & n13364 ) | ( ~n13362 & n13365 ) | ( n13364 & n13365 ) ;
  assign n13367 = n3541 & ~n10617 ;
  assign n13368 = x29 & n13367 ;
  assign n13369 = n3536 & n10275 ;
  assign n13370 = n4039 | n13369 ;
  assign n13371 = ( ~n10297 & n13369 ) | ( ~n10297 & n13370 ) | ( n13369 & n13370 ) ;
  assign n13372 = n3501 & n10273 ;
  assign n13373 = n13371 | n13372 ;
  assign n13374 = x29 & ~n13373 ;
  assign n13375 = ( ~x29 & n13367 ) | ( ~x29 & n13373 ) | ( n13367 & n13373 ) ;
  assign n13376 = ( ~n13368 & n13374 ) | ( ~n13368 & n13375 ) | ( n13374 & n13375 ) ;
  assign n13377 = n3273 & ~n10279 ;
  assign n13378 = n3270 | n13377 ;
  assign n13379 = ( n10277 & n13377 ) | ( n10277 & n13378 ) | ( n13377 & n13378 ) ;
  assign n13380 = n390 | n13379 ;
  assign n13381 = ( ~n10516 & n13379 ) | ( ~n10516 & n13380 ) | ( n13379 & n13380 ) ;
  assign n13382 = n3274 & n10291 ;
  assign n13383 = n13381 | n13382 ;
  assign n13384 = n1379 | n2307 ;
  assign n13385 = n3296 | n3375 ;
  assign n13386 = n13384 | n13385 ;
  assign n13387 = n1852 | n13386 ;
  assign n13388 = n284 | n922 ;
  assign n13389 = n708 | n13388 ;
  assign n13390 = n1448 | n13389 ;
  assign n13391 = n2164 | n2215 ;
  assign n13392 = n13390 | n13391 ;
  assign n13393 = n2500 & ~n13392 ;
  assign n13394 = n680 | n1005 ;
  assign n13395 = n1762 | n2897 ;
  assign n13396 = n13394 | n13395 ;
  assign n13397 = n360 | n533 ;
  assign n13398 = n835 | n13397 ;
  assign n13399 = n379 | n1793 ;
  assign n13400 = n13398 | n13399 ;
  assign n13401 = n13396 | n13400 ;
  assign n13402 = n13393 & ~n13401 ;
  assign n13403 = ~n13387 & n13402 ;
  assign n13404 = n341 | n517 ;
  assign n13405 = n5031 | n13404 ;
  assign n13406 = n335 | n704 ;
  assign n13407 = n4102 | n13406 ;
  assign n13408 = n13405 | n13407 ;
  assign n13409 = n900 | n946 ;
  assign n13410 = n13408 | n13409 ;
  assign n13411 = n2291 | n10140 ;
  assign n13412 = n13410 | n13411 ;
  assign n13413 = n4296 | n5442 ;
  assign n13414 = n314 | n318 ;
  assign n13415 = n13413 | n13414 ;
  assign n13416 = n1054 | n1347 ;
  assign n13417 = n1537 | n2850 ;
  assign n13418 = n13416 | n13417 ;
  assign n13419 = n13415 | n13418 ;
  assign n13420 = n13412 | n13419 ;
  assign n13421 = n3322 | n13420 ;
  assign n13422 = n13403 & ~n13421 ;
  assign n13423 = ( n13226 & n13383 ) | ( n13226 & ~n13422 ) | ( n13383 & ~n13422 ) ;
  assign n13424 = ( n13226 & ~n13383 ) | ( n13226 & n13422 ) | ( ~n13383 & n13422 ) ;
  assign n13425 = ( ~n13226 & n13423 ) | ( ~n13226 & n13424 ) | ( n13423 & n13424 ) ;
  assign n13426 = ( n13229 & n13376 ) | ( n13229 & ~n13425 ) | ( n13376 & ~n13425 ) ;
  assign n13427 = ( n13229 & ~n13376 ) | ( n13229 & n13425 ) | ( ~n13376 & n13425 ) ;
  assign n13428 = ( ~n13229 & n13426 ) | ( ~n13229 & n13427 ) | ( n13426 & n13427 ) ;
  assign n13429 = ( n13233 & n13366 ) | ( n13233 & ~n13428 ) | ( n13366 & ~n13428 ) ;
  assign n13430 = ( n13233 & ~n13366 ) | ( n13233 & n13428 ) | ( ~n13366 & n13428 ) ;
  assign n13431 = ( ~n13233 & n13429 ) | ( ~n13233 & n13430 ) | ( n13429 & n13430 ) ;
  assign n13432 = ( n13236 & n13356 ) | ( n13236 & ~n13431 ) | ( n13356 & ~n13431 ) ;
  assign n13433 = ( n13236 & ~n13356 ) | ( n13236 & n13431 ) | ( ~n13356 & n13431 ) ;
  assign n13434 = ( ~n13236 & n13432 ) | ( ~n13236 & n13433 ) | ( n13432 & n13433 ) ;
  assign n13435 = ( n13238 & ~n13346 ) | ( n13238 & n13434 ) | ( ~n13346 & n13434 ) ;
  assign n13436 = ( n13238 & n13346 ) | ( n13238 & ~n13434 ) | ( n13346 & ~n13434 ) ;
  assign n13437 = ( ~n13238 & n13435 ) | ( ~n13238 & n13436 ) | ( n13435 & n13436 ) ;
  assign n13438 = ( n13241 & n13336 ) | ( n13241 & ~n13437 ) | ( n13336 & ~n13437 ) ;
  assign n13439 = ( n13241 & ~n13336 ) | ( n13241 & n13437 ) | ( ~n13336 & n13437 ) ;
  assign n13440 = ( ~n13241 & n13438 ) | ( ~n13241 & n13439 ) | ( n13438 & n13439 ) ;
  assign n13441 = ( n13255 & n13326 ) | ( n13255 & ~n13440 ) | ( n13326 & ~n13440 ) ;
  assign n13442 = ( n13255 & ~n13326 ) | ( n13255 & n13440 ) | ( ~n13326 & n13440 ) ;
  assign n13443 = ( ~n13255 & n13441 ) | ( ~n13255 & n13442 ) | ( n13441 & n13442 ) ;
  assign n13444 = n6571 & ~n11989 ;
  assign n13445 = x11 & n13444 ;
  assign n13446 = n6570 & n10243 ;
  assign n13447 = n6796 & ~n10320 ;
  assign n13448 = n6567 & n10245 ;
  assign n13449 = n13447 | n13448 ;
  assign n13450 = n13446 | n13449 ;
  assign n13451 = x11 & ~n13450 ;
  assign n13452 = ( ~x11 & n13444 ) | ( ~x11 & n13450 ) | ( n13444 & n13450 ) ;
  assign n13453 = ( ~n13445 & n13451 ) | ( ~n13445 & n13452 ) | ( n13451 & n13452 ) ;
  assign n13454 = ( n13257 & n13443 ) | ( n13257 & n13453 ) | ( n13443 & n13453 ) ;
  assign n13455 = ( n13257 & ~n13443 ) | ( n13257 & n13453 ) | ( ~n13443 & n13453 ) ;
  assign n13456 = ( n13443 & ~n13454 ) | ( n13443 & n13455 ) | ( ~n13454 & n13455 ) ;
  assign n13457 = ( n13260 & n13316 ) | ( n13260 & ~n13456 ) | ( n13316 & ~n13456 ) ;
  assign n13458 = ( ~n13260 & n13316 ) | ( ~n13260 & n13456 ) | ( n13316 & n13456 ) ;
  assign n13459 = ( ~n13316 & n13457 ) | ( ~n13316 & n13458 ) | ( n13457 & n13458 ) ;
  assign n13460 = ( n13263 & ~n13306 ) | ( n13263 & n13459 ) | ( ~n13306 & n13459 ) ;
  assign n13461 = ( n13263 & n13306 ) | ( n13263 & ~n13459 ) | ( n13306 & ~n13459 ) ;
  assign n13462 = ( ~n13263 & n13460 ) | ( ~n13263 & n13461 ) | ( n13460 & n13461 ) ;
  assign n13463 = ( n13266 & n13296 ) | ( n13266 & ~n13462 ) | ( n13296 & ~n13462 ) ;
  assign n13464 = ( n66 & n10230 ) | ( n66 & ~n13276 ) | ( n10230 & ~n13276 ) ;
  assign n13465 = ( ~n10230 & n13275 ) | ( ~n10230 & n13464 ) | ( n13275 & n13464 ) ;
  assign n13466 = n13276 | n13464 ;
  assign n13467 = ( ~n66 & n13465 ) | ( ~n66 & n13466 ) | ( n13465 & n13466 ) ;
  assign n13468 = ~n10234 & n13467 ;
  assign n13469 = n66 & ~n13275 ;
  assign n13470 = n10230 & n13277 ;
  assign n13471 = n13469 | n13470 ;
  assign n13472 = n10234 & ~n13471 ;
  assign n13473 = n13468 | n13472 ;
  assign n13474 = n13267 | n13280 ;
  assign n13475 = n13473 | n13474 ;
  assign n13476 = n13473 & n13474 ;
  assign n13477 = n13475 & ~n13476 ;
  assign n13478 = n13284 & ~n13473 ;
  assign n13479 = n13284 & ~n13478 ;
  assign n13480 = ( n13477 & ~n13478 ) | ( n13477 & n13479 ) | ( ~n13478 & n13479 ) ;
  assign n13481 = n9593 & ~n13473 ;
  assign n13482 = n9592 | n13481 ;
  assign n13483 = ( ~n13480 & n13481 ) | ( ~n13480 & n13482 ) | ( n13481 & n13482 ) ;
  assign n13484 = n41 & ~n13280 ;
  assign n13485 = ( x2 & ~n13483 ) | ( x2 & n13484 ) | ( ~n13483 & n13484 ) ;
  assign n13486 = ~x2 & n13483 ;
  assign n13487 = n9600 & ~n10235 ;
  assign n13488 = ( x2 & n13484 ) | ( x2 & n13487 ) | ( n13484 & n13487 ) ;
  assign n13489 = ( n13485 & n13486 ) | ( n13485 & ~n13488 ) | ( n13486 & ~n13488 ) ;
  assign n13490 = n40 & n10214 ;
  assign n13491 = n8721 & ~n10237 ;
  assign n13492 = n8340 & ~n10332 ;
  assign n13493 = n13491 | n13492 ;
  assign n13494 = n13490 | n13493 ;
  assign n13495 = x5 & n13494 ;
  assign n13496 = n8341 & n12953 ;
  assign n13497 = ( ~x5 & n13494 ) | ( ~x5 & n13496 ) | ( n13494 & n13496 ) ;
  assign n13498 = x5 & ~n13496 ;
  assign n13499 = ( ~n13495 & n13497 ) | ( ~n13495 & n13498 ) | ( n13497 & n13498 ) ;
  assign n13500 = n7644 & n10326 ;
  assign n13501 = x8 & n13500 ;
  assign n13502 = n7341 & n10239 ;
  assign n13503 = n7345 | n13502 ;
  assign n13504 = ( n10329 & n13502 ) | ( n10329 & n13503 ) | ( n13502 & n13503 ) ;
  assign n13505 = n7346 | n13504 ;
  assign n13506 = ( n10397 & n13504 ) | ( n10397 & n13505 ) | ( n13504 & n13505 ) ;
  assign n13507 = x8 & ~n13506 ;
  assign n13508 = ( ~x8 & n13500 ) | ( ~x8 & n13506 ) | ( n13500 & n13506 ) ;
  assign n13509 = ( ~n13501 & n13507 ) | ( ~n13501 & n13508 ) | ( n13507 & n13508 ) ;
  assign n13510 = n6796 & n10243 ;
  assign n13511 = x11 & n13510 ;
  assign n13512 = n6567 & ~n10320 ;
  assign n13513 = n6570 | n13512 ;
  assign n13514 = ( n10241 & n13512 ) | ( n10241 & n13513 ) | ( n13512 & n13513 ) ;
  assign n13515 = n6571 | n13514 ;
  assign n13516 = ( n12105 & n13514 ) | ( n12105 & n13515 ) | ( n13514 & n13515 ) ;
  assign n13517 = x11 & ~n13516 ;
  assign n13518 = ( ~x11 & n13510 ) | ( ~x11 & n13516 ) | ( n13510 & n13516 ) ;
  assign n13519 = ( ~n13511 & n13517 ) | ( ~n13511 & n13518 ) | ( n13517 & n13518 ) ;
  assign n13520 = n6332 & ~n10316 ;
  assign n13521 = x14 & n13520 ;
  assign n13522 = n5909 & n10247 ;
  assign n13523 = n5914 | n13522 ;
  assign n13524 = ( n10245 & n13522 ) | ( n10245 & n13523 ) | ( n13522 & n13523 ) ;
  assign n13525 = n5915 | n13524 ;
  assign n13526 = ( ~n11676 & n13524 ) | ( ~n11676 & n13525 ) | ( n13524 & n13525 ) ;
  assign n13527 = x14 & ~n13526 ;
  assign n13528 = ( ~x14 & n13520 ) | ( ~x14 & n13526 ) | ( n13520 & n13526 ) ;
  assign n13529 = ( ~n13521 & n13527 ) | ( ~n13521 & n13528 ) | ( n13527 & n13528 ) ;
  assign n13530 = n5417 & n10312 ;
  assign n13531 = x17 & n13530 ;
  assign n13532 = n5584 & ~n10249 ;
  assign n13533 = n5413 & n10251 ;
  assign n13534 = n13532 | n13533 ;
  assign n13535 = n5418 | n13534 ;
  assign n13536 = ( ~n11486 & n13534 ) | ( ~n11486 & n13535 ) | ( n13534 & n13535 ) ;
  assign n13537 = x17 & ~n13536 ;
  assign n13538 = ( ~x17 & n13530 ) | ( ~x17 & n13536 ) | ( n13530 & n13536 ) ;
  assign n13539 = ( ~n13531 & n13537 ) | ( ~n13531 & n13538 ) | ( n13537 & n13538 ) ;
  assign n13540 = n4879 & ~n11297 ;
  assign n13541 = x20 & n13540 ;
  assign n13542 = n4874 & n10257 ;
  assign n13543 = n4878 | n13542 ;
  assign n13544 = ( ~n10253 & n13542 ) | ( ~n10253 & n13543 ) | ( n13542 & n13543 ) ;
  assign n13545 = n5232 & n10255 ;
  assign n13546 = n13544 | n13545 ;
  assign n13547 = x20 & ~n13546 ;
  assign n13548 = ( ~x20 & n13540 ) | ( ~x20 & n13546 ) | ( n13540 & n13546 ) ;
  assign n13549 = ( ~n13541 & n13547 ) | ( ~n13541 & n13548 ) | ( n13547 & n13548 ) ;
  assign n13550 = n4637 & n10261 ;
  assign n13551 = x23 & n13550 ;
  assign n13552 = n4584 & n10263 ;
  assign n13553 = n4649 | n13552 ;
  assign n13554 = ( n10259 & n13552 ) | ( n10259 & n13553 ) | ( n13552 & n13553 ) ;
  assign n13555 = n4591 | n13554 ;
  assign n13556 = ( n10859 & n13554 ) | ( n10859 & n13555 ) | ( n13554 & n13555 ) ;
  assign n13557 = x23 & ~n13556 ;
  assign n13558 = ( ~x23 & n13550 ) | ( ~x23 & n13556 ) | ( n13550 & n13556 ) ;
  assign n13559 = ( ~n13551 & n13557 ) | ( ~n13551 & n13558 ) | ( n13557 & n13558 ) ;
  assign n13560 = n3541 & ~n10656 ;
  assign n13561 = x29 & n13560 ;
  assign n13562 = n3536 & n10273 ;
  assign n13563 = n4039 | n13562 ;
  assign n13564 = ( n10271 & n13562 ) | ( n10271 & n13563 ) | ( n13562 & n13563 ) ;
  assign n13565 = n3501 & ~n10297 ;
  assign n13566 = n13564 | n13565 ;
  assign n13567 = x29 & ~n13566 ;
  assign n13568 = ( ~x29 & n13560 ) | ( ~x29 & n13566 ) | ( n13560 & n13566 ) ;
  assign n13569 = ( ~n13561 & n13567 ) | ( ~n13561 & n13568 ) | ( n13567 & n13568 ) ;
  assign n13570 = n390 & n10563 ;
  assign n13571 = n3270 & n10275 ;
  assign n13572 = n3274 & n10277 ;
  assign n13573 = n3273 & n10291 ;
  assign n13574 = n13572 | n13573 ;
  assign n13575 = n13571 | n13574 ;
  assign n13576 = n13570 | n13575 ;
  assign n13577 = n2321 | n3460 ;
  assign n13578 = n545 | n589 ;
  assign n13579 = n1672 | n13578 ;
  assign n13580 = n500 | n794 ;
  assign n13581 = n13579 | n13580 ;
  assign n13582 = ( n3916 & ~n13577 ) | ( n3916 & n13581 ) | ( ~n13577 & n13581 ) ;
  assign n13583 = n13577 | n13582 ;
  assign n13584 = n262 | n2420 ;
  assign n13585 = n1857 | n13584 ;
  assign n13586 = n113 | n218 ;
  assign n13587 = n3037 | n13586 ;
  assign n13588 = n13585 | n13587 ;
  assign n13589 = n225 | n468 ;
  assign n13590 = n324 | n13589 ;
  assign n13591 = n3205 | n13590 ;
  assign n13592 = n6171 | n13591 ;
  assign n13593 = n13588 | n13592 ;
  assign n13594 = n13583 | n13593 ;
  assign n13595 = n276 | n557 ;
  assign n13596 = n3010 | n13595 ;
  assign n13597 = n929 | n2901 ;
  assign n13598 = n1400 | n13597 ;
  assign n13599 = n13596 | n13598 ;
  assign n13600 = n13594 | n13599 ;
  assign n13601 = n303 | n1176 ;
  assign n13602 = n3395 | n13601 ;
  assign n13603 = n3390 | n13602 ;
  assign n13604 = n2027 | n13603 ;
  assign n13605 = n3921 | n13604 ;
  assign n13606 = n176 | n860 ;
  assign n13607 = n254 | n285 ;
  assign n13608 = n13606 | n13607 ;
  assign n13609 = n1663 | n13608 ;
  assign n13610 = n199 | n4253 ;
  assign n13611 = n13609 | n13610 ;
  assign n13612 = n13605 | n13611 ;
  assign n13613 = n6082 | n13612 ;
  assign n13614 = n13600 | n13613 ;
  assign n13615 = n2511 | n3733 ;
  assign n13616 = n5063 | n13615 ;
  assign n13617 = n644 | n722 ;
  assign n13618 = n13616 | n13617 ;
  assign n13619 = n2836 | n3638 ;
  assign n13620 = n3569 | n13619 ;
  assign n13621 = n488 | n662 ;
  assign n13622 = n2648 | n13621 ;
  assign n13623 = n222 | n3052 ;
  assign n13624 = n141 | n13623 ;
  assign n13625 = n13622 | n13624 ;
  assign n13626 = n3566 | n13625 ;
  assign n13627 = n13620 | n13626 ;
  assign n13628 = n13618 | n13627 ;
  assign n13629 = n13614 | n13628 ;
  assign n13630 = ( n13423 & n13576 ) | ( n13423 & n13629 ) | ( n13576 & n13629 ) ;
  assign n13631 = ( ~n13423 & n13576 ) | ( ~n13423 & n13629 ) | ( n13576 & n13629 ) ;
  assign n13632 = ( n13423 & ~n13630 ) | ( n13423 & n13631 ) | ( ~n13630 & n13631 ) ;
  assign n13633 = ( ~n13426 & n13569 ) | ( ~n13426 & n13632 ) | ( n13569 & n13632 ) ;
  assign n13634 = ( n13426 & n13569 ) | ( n13426 & n13632 ) | ( n13569 & n13632 ) ;
  assign n13635 = ( n13426 & n13633 ) | ( n13426 & ~n13634 ) | ( n13633 & ~n13634 ) ;
  assign n13636 = n4203 & n10804 ;
  assign n13637 = x26 & n13636 ;
  assign n13638 = n4215 & n10265 ;
  assign n13639 = n4200 & n10267 ;
  assign n13640 = n2083 & ~n10269 ;
  assign n13641 = n13639 | n13640 ;
  assign n13642 = n13638 | n13641 ;
  assign n13643 = x26 & ~n13642 ;
  assign n13644 = ( ~x26 & n13636 ) | ( ~x26 & n13642 ) | ( n13636 & n13642 ) ;
  assign n13645 = ( ~n13637 & n13643 ) | ( ~n13637 & n13644 ) | ( n13643 & n13644 ) ;
  assign n13646 = ( n13429 & n13635 ) | ( n13429 & n13645 ) | ( n13635 & n13645 ) ;
  assign n13647 = ( ~n13429 & n13635 ) | ( ~n13429 & n13645 ) | ( n13635 & n13645 ) ;
  assign n13648 = ( n13429 & ~n13646 ) | ( n13429 & n13647 ) | ( ~n13646 & n13647 ) ;
  assign n13649 = ( ~n13432 & n13559 ) | ( ~n13432 & n13648 ) | ( n13559 & n13648 ) ;
  assign n13650 = ( n13432 & n13559 ) | ( n13432 & n13648 ) | ( n13559 & n13648 ) ;
  assign n13651 = ( n13432 & n13649 ) | ( n13432 & ~n13650 ) | ( n13649 & ~n13650 ) ;
  assign n13652 = ( ~n13436 & n13549 ) | ( ~n13436 & n13651 ) | ( n13549 & n13651 ) ;
  assign n13653 = ( n13436 & n13549 ) | ( n13436 & n13651 ) | ( n13549 & n13651 ) ;
  assign n13654 = ( n13436 & n13652 ) | ( n13436 & ~n13653 ) | ( n13652 & ~n13653 ) ;
  assign n13655 = ( ~n13438 & n13539 ) | ( ~n13438 & n13654 ) | ( n13539 & n13654 ) ;
  assign n13656 = ( n13438 & n13539 ) | ( n13438 & n13654 ) | ( n13539 & n13654 ) ;
  assign n13657 = ( n13438 & n13655 ) | ( n13438 & ~n13656 ) | ( n13655 & ~n13656 ) ;
  assign n13658 = ( ~n13441 & n13529 ) | ( ~n13441 & n13657 ) | ( n13529 & n13657 ) ;
  assign n13659 = ( n13441 & n13529 ) | ( n13441 & n13657 ) | ( n13529 & n13657 ) ;
  assign n13660 = ( n13441 & n13658 ) | ( n13441 & ~n13659 ) | ( n13658 & ~n13659 ) ;
  assign n13661 = ( ~n13455 & n13519 ) | ( ~n13455 & n13660 ) | ( n13519 & n13660 ) ;
  assign n13662 = ( n13455 & n13519 ) | ( n13455 & n13660 ) | ( n13519 & n13660 ) ;
  assign n13663 = ( n13455 & n13661 ) | ( n13455 & ~n13662 ) | ( n13661 & ~n13662 ) ;
  assign n13664 = ( n13457 & n13509 ) | ( n13457 & n13663 ) | ( n13509 & n13663 ) ;
  assign n13665 = ( ~n13457 & n13509 ) | ( ~n13457 & n13663 ) | ( n13509 & n13663 ) ;
  assign n13666 = ( n13457 & ~n13664 ) | ( n13457 & n13665 ) | ( ~n13664 & n13665 ) ;
  assign n13667 = ( ~n13461 & n13499 ) | ( ~n13461 & n13666 ) | ( n13499 & n13666 ) ;
  assign n13668 = ( n13461 & n13499 ) | ( n13461 & n13666 ) | ( n13499 & n13666 ) ;
  assign n13669 = ( n13461 & n13667 ) | ( n13461 & ~n13668 ) | ( n13667 & ~n13668 ) ;
  assign n13670 = ( n13463 & n13489 ) | ( n13463 & n13669 ) | ( n13489 & n13669 ) ;
  assign n13671 = n13474 & ~n13478 ;
  assign n13672 = n9592 & n13671 ;
  assign n13673 = n41 & ~n13473 ;
  assign n13674 = n9593 | n13673 ;
  assign n13675 = ( n13475 & n13673 ) | ( n13475 & n13674 ) | ( n13673 & n13674 ) ;
  assign n13676 = ( x2 & ~n13672 ) | ( x2 & n13675 ) | ( ~n13672 & n13675 ) ;
  assign n13677 = ~x2 & n13672 ;
  assign n13678 = ( x2 & n9155 ) | ( x2 & ~n13280 ) | ( n9155 & ~n13280 ) ;
  assign n13679 = ( n9600 & n13675 ) | ( n9600 & n13678 ) | ( n13675 & n13678 ) ;
  assign n13680 = ( n13676 & n13677 ) | ( n13676 & ~n13679 ) | ( n13677 & ~n13679 ) ;
  assign n13681 = n40 & ~n10235 ;
  assign n13682 = n8721 & n10214 ;
  assign n13683 = n8340 & ~n10237 ;
  assign n13684 = n13682 | n13683 ;
  assign n13685 = n13681 | n13684 ;
  assign n13686 = x5 & n13685 ;
  assign n13687 = n8341 & n10371 ;
  assign n13688 = ( ~x5 & n13685 ) | ( ~x5 & n13687 ) | ( n13685 & n13687 ) ;
  assign n13689 = x5 & ~n13687 ;
  assign n13690 = ( ~n13686 & n13688 ) | ( ~n13686 & n13689 ) | ( n13688 & n13689 ) ;
  assign n13691 = n7644 & n10329 ;
  assign n13692 = x8 & n13691 ;
  assign n13693 = n7341 & n10326 ;
  assign n13694 = n7345 | n13693 ;
  assign n13695 = ( ~n10332 & n13693 ) | ( ~n10332 & n13694 ) | ( n13693 & n13694 ) ;
  assign n13696 = n7346 | n13695 ;
  assign n13697 = ( ~n10383 & n13695 ) | ( ~n10383 & n13696 ) | ( n13695 & n13696 ) ;
  assign n13698 = x8 & ~n13697 ;
  assign n13699 = ( ~x8 & n13691 ) | ( ~x8 & n13697 ) | ( n13691 & n13697 ) ;
  assign n13700 = ( ~n13692 & n13698 ) | ( ~n13692 & n13699 ) | ( n13698 & n13699 ) ;
  assign n13701 = n6571 & n12575 ;
  assign n13702 = x11 & n13701 ;
  assign n13703 = n6567 & n10243 ;
  assign n13704 = n6570 | n13703 ;
  assign n13705 = ( n10239 & n13703 ) | ( n10239 & n13704 ) | ( n13703 & n13704 ) ;
  assign n13706 = n6796 & n10241 ;
  assign n13707 = n13705 | n13706 ;
  assign n13708 = x11 & ~n13707 ;
  assign n13709 = ( ~x11 & n13701 ) | ( ~x11 & n13707 ) | ( n13701 & n13707 ) ;
  assign n13710 = ( ~n13702 & n13708 ) | ( ~n13702 & n13709 ) | ( n13708 & n13709 ) ;
  assign n13711 = n5914 & ~n10320 ;
  assign n13712 = x14 & n13711 ;
  assign n13713 = n6332 & n10245 ;
  assign n13714 = n5909 & ~n10316 ;
  assign n13715 = n13713 | n13714 ;
  assign n13716 = n5915 | n13715 ;
  assign n13717 = ( ~n10414 & n13715 ) | ( ~n10414 & n13716 ) | ( n13715 & n13716 ) ;
  assign n13718 = x14 & ~n13717 ;
  assign n13719 = ( ~x14 & n13711 ) | ( ~x14 & n13717 ) | ( n13711 & n13717 ) ;
  assign n13720 = ( ~n13712 & n13718 ) | ( ~n13712 & n13719 ) | ( n13718 & n13719 ) ;
  assign n13721 = n5418 & n10428 ;
  assign n13722 = x17 & n13721 ;
  assign n13723 = n5413 & ~n10249 ;
  assign n13724 = n5417 | n13723 ;
  assign n13725 = ( n10247 & n13723 ) | ( n10247 & n13724 ) | ( n13723 & n13724 ) ;
  assign n13726 = n5584 & n10312 ;
  assign n13727 = n13725 | n13726 ;
  assign n13728 = x17 & ~n13727 ;
  assign n13729 = ( ~x17 & n13721 ) | ( ~x17 & n13727 ) | ( n13721 & n13727 ) ;
  assign n13730 = ( ~n13722 & n13728 ) | ( ~n13722 & n13729 ) | ( n13728 & n13729 ) ;
  assign n13731 = n4879 & ~n11309 ;
  assign n13732 = x20 & n13731 ;
  assign n13733 = n4874 & n10255 ;
  assign n13734 = n4878 | n13733 ;
  assign n13735 = ( n10251 & n13733 ) | ( n10251 & n13734 ) | ( n13733 & n13734 ) ;
  assign n13736 = n5232 & ~n10253 ;
  assign n13737 = n13735 | n13736 ;
  assign n13738 = x20 & ~n13737 ;
  assign n13739 = ( ~x20 & n13731 ) | ( ~x20 & n13737 ) | ( n13731 & n13737 ) ;
  assign n13740 = ( ~n13732 & n13738 ) | ( ~n13732 & n13739 ) | ( n13738 & n13739 ) ;
  assign n13741 = n4637 & n10259 ;
  assign n13742 = x23 & n13741 ;
  assign n13743 = n4584 & n10261 ;
  assign n13744 = n4649 | n13743 ;
  assign n13745 = ( n10257 & n13743 ) | ( n10257 & n13744 ) | ( n13743 & n13744 ) ;
  assign n13746 = n4591 | n13745 ;
  assign n13747 = ( n11065 & n13745 ) | ( n11065 & n13746 ) | ( n13745 & n13746 ) ;
  assign n13748 = x23 & ~n13747 ;
  assign n13749 = ( ~x23 & n13741 ) | ( ~x23 & n13747 ) | ( n13741 & n13747 ) ;
  assign n13750 = ( ~n13742 & n13748 ) | ( ~n13742 & n13749 ) | ( n13748 & n13749 ) ;
  assign n13751 = n4039 & ~n10269 ;
  assign n13752 = n3541 | n13751 ;
  assign n13753 = ( ~n10698 & n13751 ) | ( ~n10698 & n13752 ) | ( n13751 & n13752 ) ;
  assign n13754 = n3536 & ~n10297 ;
  assign n13755 = ( ~x29 & n13753 ) | ( ~x29 & n13754 ) | ( n13753 & n13754 ) ;
  assign n13756 = n3501 & n10271 ;
  assign n13757 = x29 & ~n13754 ;
  assign n13758 = n13756 | n13757 ;
  assign n13759 = ( n13753 & n13756 ) | ( n13753 & n13757 ) | ( n13756 & n13757 ) ;
  assign n13760 = ( n13755 & n13758 ) | ( n13755 & ~n13759 ) | ( n13758 & ~n13759 ) ;
  assign n13761 = n3273 & n10277 ;
  assign n13762 = n3270 | n13761 ;
  assign n13763 = ( n10273 & n13761 ) | ( n10273 & n13762 ) | ( n13761 & n13762 ) ;
  assign n13764 = n390 | n13763 ;
  assign n13765 = ( n10577 & n13763 ) | ( n10577 & n13764 ) | ( n13763 & n13764 ) ;
  assign n13766 = n3274 & n10275 ;
  assign n13767 = n13765 | n13766 ;
  assign n13768 = n577 | n12669 ;
  assign n13769 = n87 | n104 ;
  assign n13770 = n239 | n13769 ;
  assign n13771 = n4353 | n4509 ;
  assign n13772 = n2288 | n13771 ;
  assign n13773 = n13770 | n13772 ;
  assign n13774 = n13768 | n13773 ;
  assign n13775 = n1904 | n2058 ;
  assign n13776 = n3638 | n13775 ;
  assign n13777 = n2304 | n13776 ;
  assign n13778 = n13774 | n13777 ;
  assign n13779 = n3961 | n13778 ;
  assign n13780 = n3790 | n13779 ;
  assign n13781 = ( n13630 & n13767 ) | ( n13630 & n13780 ) | ( n13767 & n13780 ) ;
  assign n13782 = ( ~n13630 & n13767 ) | ( ~n13630 & n13780 ) | ( n13767 & n13780 ) ;
  assign n13783 = ( n13630 & ~n13781 ) | ( n13630 & n13782 ) | ( ~n13781 & n13782 ) ;
  assign n13784 = ( ~n13634 & n13760 ) | ( ~n13634 & n13783 ) | ( n13760 & n13783 ) ;
  assign n13785 = ( n13634 & n13760 ) | ( n13634 & n13783 ) | ( n13760 & n13783 ) ;
  assign n13786 = ( n13634 & n13784 ) | ( n13634 & ~n13785 ) | ( n13784 & ~n13785 ) ;
  assign n13787 = n4215 & n10263 ;
  assign n13788 = n4200 & n10265 ;
  assign n13789 = n2083 & n10267 ;
  assign n13790 = n13788 | n13789 ;
  assign n13791 = n13787 | n13790 ;
  assign n13792 = x26 & n13791 ;
  assign n13793 = n4203 & n10874 ;
  assign n13794 = ( ~x26 & n13791 ) | ( ~x26 & n13793 ) | ( n13791 & n13793 ) ;
  assign n13795 = x26 & ~n13793 ;
  assign n13796 = ( ~n13792 & n13794 ) | ( ~n13792 & n13795 ) | ( n13794 & n13795 ) ;
  assign n13797 = ( ~n13646 & n13786 ) | ( ~n13646 & n13796 ) | ( n13786 & n13796 ) ;
  assign n13798 = ( n13646 & n13786 ) | ( n13646 & n13796 ) | ( n13786 & n13796 ) ;
  assign n13799 = ( n13646 & n13797 ) | ( n13646 & ~n13798 ) | ( n13797 & ~n13798 ) ;
  assign n13800 = ( n13650 & n13750 ) | ( n13650 & n13799 ) | ( n13750 & n13799 ) ;
  assign n13801 = ( ~n13650 & n13750 ) | ( ~n13650 & n13799 ) | ( n13750 & n13799 ) ;
  assign n13802 = ( n13650 & ~n13800 ) | ( n13650 & n13801 ) | ( ~n13800 & n13801 ) ;
  assign n13803 = ( ~n13653 & n13740 ) | ( ~n13653 & n13802 ) | ( n13740 & n13802 ) ;
  assign n13804 = ( n13653 & n13740 ) | ( n13653 & n13802 ) | ( n13740 & n13802 ) ;
  assign n13805 = ( n13653 & n13803 ) | ( n13653 & ~n13804 ) | ( n13803 & ~n13804 ) ;
  assign n13806 = ( n13656 & n13730 ) | ( n13656 & n13805 ) | ( n13730 & n13805 ) ;
  assign n13807 = ( ~n13656 & n13730 ) | ( ~n13656 & n13805 ) | ( n13730 & n13805 ) ;
  assign n13808 = ( n13656 & ~n13806 ) | ( n13656 & n13807 ) | ( ~n13806 & n13807 ) ;
  assign n13809 = ( ~n13659 & n13720 ) | ( ~n13659 & n13808 ) | ( n13720 & n13808 ) ;
  assign n13810 = ( n13659 & n13720 ) | ( n13659 & n13808 ) | ( n13720 & n13808 ) ;
  assign n13811 = ( n13659 & n13809 ) | ( n13659 & ~n13810 ) | ( n13809 & ~n13810 ) ;
  assign n13812 = ( ~n13662 & n13710 ) | ( ~n13662 & n13811 ) | ( n13710 & n13811 ) ;
  assign n13813 = ( n13662 & n13710 ) | ( n13662 & n13811 ) | ( n13710 & n13811 ) ;
  assign n13814 = ( n13662 & n13812 ) | ( n13662 & ~n13813 ) | ( n13812 & ~n13813 ) ;
  assign n13815 = ( ~n13664 & n13700 ) | ( ~n13664 & n13814 ) | ( n13700 & n13814 ) ;
  assign n13816 = ( n13664 & n13700 ) | ( n13664 & n13814 ) | ( n13700 & n13814 ) ;
  assign n13817 = ( n13664 & n13815 ) | ( n13664 & ~n13816 ) | ( n13815 & ~n13816 ) ;
  assign n13818 = ( n13668 & n13690 ) | ( n13668 & n13817 ) | ( n13690 & n13817 ) ;
  assign n13819 = ( n13668 & ~n13690 ) | ( n13668 & n13817 ) | ( ~n13690 & n13817 ) ;
  assign n13820 = ( n13690 & ~n13818 ) | ( n13690 & n13819 ) | ( ~n13818 & n13819 ) ;
  assign n13821 = ( n13670 & n13680 ) | ( n13670 & n13820 ) | ( n13680 & n13820 ) ;
  assign n13822 = n40 & ~n13280 ;
  assign n13823 = n8721 & ~n10235 ;
  assign n13824 = n8340 & n10214 ;
  assign n13825 = n13823 | n13824 ;
  assign n13826 = n13822 | n13825 ;
  assign n13827 = x5 & n13826 ;
  assign n13828 = n8341 & ~n13285 ;
  assign n13829 = ( ~x5 & n13826 ) | ( ~x5 & n13828 ) | ( n13826 & n13828 ) ;
  assign n13830 = x5 & ~n13828 ;
  assign n13831 = ( ~n13827 & n13829 ) | ( ~n13827 & n13830 ) | ( n13829 & n13830 ) ;
  assign n13832 = n7345 & ~n10237 ;
  assign n13833 = n7644 & ~n10332 ;
  assign n13834 = n7341 & n10329 ;
  assign n13835 = n13833 | n13834 ;
  assign n13836 = n13832 | n13835 ;
  assign n13837 = x8 & n13836 ;
  assign n13838 = n7346 & n12756 ;
  assign n13839 = ( ~x8 & n13836 ) | ( ~x8 & n13838 ) | ( n13836 & n13838 ) ;
  assign n13840 = x8 & ~n13838 ;
  assign n13841 = ( ~n13837 & n13839 ) | ( ~n13837 & n13840 ) | ( n13839 & n13840 ) ;
  assign n13842 = n6796 & n10239 ;
  assign n13843 = x11 & n13842 ;
  assign n13844 = n6567 & n10241 ;
  assign n13845 = n6570 | n13844 ;
  assign n13846 = ( n10326 & n13844 ) | ( n10326 & n13845 ) | ( n13844 & n13845 ) ;
  assign n13847 = n6571 | n13846 ;
  assign n13848 = ( n12222 & n13846 ) | ( n12222 & n13847 ) | ( n13846 & n13847 ) ;
  assign n13849 = x11 & ~n13848 ;
  assign n13850 = ( ~x11 & n13842 ) | ( ~x11 & n13848 ) | ( n13842 & n13848 ) ;
  assign n13851 = ( ~n13843 & n13849 ) | ( ~n13843 & n13850 ) | ( n13849 & n13850 ) ;
  assign n13852 = n5915 & ~n11989 ;
  assign n13853 = x14 & n13852 ;
  assign n13854 = n5914 & n10243 ;
  assign n13855 = n6332 & ~n10320 ;
  assign n13856 = n5909 & n10245 ;
  assign n13857 = n13855 | n13856 ;
  assign n13858 = n13854 | n13857 ;
  assign n13859 = x14 & ~n13858 ;
  assign n13860 = ( ~x14 & n13852 ) | ( ~x14 & n13858 ) | ( n13852 & n13858 ) ;
  assign n13861 = ( ~n13853 & n13859 ) | ( ~n13853 & n13860 ) | ( n13859 & n13860 ) ;
  assign n13862 = n5584 & n10247 ;
  assign n13863 = x17 & n13862 ;
  assign n13864 = n5413 & n10312 ;
  assign n13865 = n5417 | n13864 ;
  assign n13866 = ( ~n10316 & n13864 ) | ( ~n10316 & n13865 ) | ( n13864 & n13865 ) ;
  assign n13867 = n5418 | n13866 ;
  assign n13868 = ( ~n11691 & n13866 ) | ( ~n11691 & n13867 ) | ( n13866 & n13867 ) ;
  assign n13869 = x17 & ~n13868 ;
  assign n13870 = ( ~x17 & n13862 ) | ( ~x17 & n13868 ) | ( n13862 & n13868 ) ;
  assign n13871 = ( ~n13863 & n13869 ) | ( ~n13863 & n13870 ) | ( n13869 & n13870 ) ;
  assign n13872 = n5232 & n10251 ;
  assign n13873 = x20 & n13872 ;
  assign n13874 = n4874 & ~n10253 ;
  assign n13875 = n4878 | n13874 ;
  assign n13876 = ( ~n10249 & n13874 ) | ( ~n10249 & n13875 ) | ( n13874 & n13875 ) ;
  assign n13877 = n4879 | n13876 ;
  assign n13878 = ( ~n10441 & n13876 ) | ( ~n10441 & n13877 ) | ( n13876 & n13877 ) ;
  assign n13879 = x20 & ~n13878 ;
  assign n13880 = ( ~x20 & n13872 ) | ( ~x20 & n13878 ) | ( n13872 & n13878 ) ;
  assign n13881 = ( ~n13873 & n13879 ) | ( ~n13873 & n13880 ) | ( n13879 & n13880 ) ;
  assign n13882 = n4637 & n10257 ;
  assign n13883 = x23 & n13882 ;
  assign n13884 = n4584 & n10259 ;
  assign n13885 = n4649 | n13884 ;
  assign n13886 = ( n10255 & n13884 ) | ( n10255 & n13885 ) | ( n13884 & n13885 ) ;
  assign n13887 = n4591 | n13886 ;
  assign n13888 = ( n11148 & n13886 ) | ( n11148 & n13887 ) | ( n13886 & n13887 ) ;
  assign n13889 = x23 & ~n13888 ;
  assign n13890 = ( ~x23 & n13882 ) | ( ~x23 & n13888 ) | ( n13882 & n13888 ) ;
  assign n13891 = ( ~n13883 & n13889 ) | ( ~n13883 & n13890 ) | ( n13889 & n13890 ) ;
  assign n13892 = n3541 & ~n10787 ;
  assign n13893 = x29 & n13892 ;
  assign n13894 = n3536 & n10271 ;
  assign n13895 = n4039 | n13894 ;
  assign n13896 = ( n10267 & n13894 ) | ( n10267 & n13895 ) | ( n13894 & n13895 ) ;
  assign n13897 = n3501 & ~n10269 ;
  assign n13898 = n13896 | n13897 ;
  assign n13899 = x29 & ~n13898 ;
  assign n13900 = ( ~x29 & n13892 ) | ( ~x29 & n13898 ) | ( n13892 & n13898 ) ;
  assign n13901 = ( ~n13893 & n13899 ) | ( ~n13893 & n13900 ) | ( n13899 & n13900 ) ;
  assign n13902 = n3273 & n10275 ;
  assign n13903 = n3270 | n13902 ;
  assign n13904 = ( ~n10297 & n13902 ) | ( ~n10297 & n13903 ) | ( n13902 & n13903 ) ;
  assign n13905 = n390 | n13904 ;
  assign n13906 = ( ~n10617 & n13904 ) | ( ~n10617 & n13905 ) | ( n13904 & n13905 ) ;
  assign n13907 = n3274 & n10273 ;
  assign n13908 = n13906 | n13907 ;
  assign n13909 = n3797 | n4953 ;
  assign n13910 = n3874 | n13909 ;
  assign n13911 = n350 | n1257 ;
  assign n13912 = n2566 | n5071 ;
  assign n13913 = n13911 | n13912 ;
  assign n13914 = n2648 | n13913 ;
  assign n13915 = n2251 | n13914 ;
  assign n13916 = n13910 | n13915 ;
  assign n13917 = n113 | n285 ;
  assign n13918 = n1895 | n13917 ;
  assign n13919 = n1178 | n13918 ;
  assign n13920 = n201 | n428 ;
  assign n13921 = n2890 | n13920 ;
  assign n13922 = n13919 | n13921 ;
  assign n13923 = n13916 | n13922 ;
  assign n13924 = n276 | n287 ;
  assign n13925 = n2018 | n13924 ;
  assign n13926 = n2212 | n13925 ;
  assign n13927 = n13923 | n13926 ;
  assign n13928 = n1560 | n1626 ;
  assign n13929 = n1698 | n13580 ;
  assign n13930 = n13928 | n13929 ;
  assign n13931 = n3107 | n13930 ;
  assign n13932 = n13775 | n13931 ;
  assign n13933 = n165 | n742 ;
  assign n13934 = n3562 | n13933 ;
  assign n13935 = n4382 | n13934 ;
  assign n13936 = n13932 | n13935 ;
  assign n13937 = n2970 | n13936 ;
  assign n13938 = n2281 | n13937 ;
  assign n13939 = n13927 | n13938 ;
  assign n13940 = ( n13781 & n13908 ) | ( n13781 & n13939 ) | ( n13908 & n13939 ) ;
  assign n13941 = ( ~n13781 & n13908 ) | ( ~n13781 & n13939 ) | ( n13908 & n13939 ) ;
  assign n13942 = ( n13781 & ~n13940 ) | ( n13781 & n13941 ) | ( ~n13940 & n13941 ) ;
  assign n13943 = ( ~n13785 & n13901 ) | ( ~n13785 & n13942 ) | ( n13901 & n13942 ) ;
  assign n13944 = ( n13785 & n13901 ) | ( n13785 & n13942 ) | ( n13901 & n13942 ) ;
  assign n13945 = ( n13785 & n13943 ) | ( n13785 & ~n13944 ) | ( n13943 & ~n13944 ) ;
  assign n13946 = n4215 & n10261 ;
  assign n13947 = n4200 & n10263 ;
  assign n13948 = n2083 & n10265 ;
  assign n13949 = n13947 | n13948 ;
  assign n13950 = n13946 | n13949 ;
  assign n13951 = x26 & n13950 ;
  assign n13952 = n4203 & n11049 ;
  assign n13953 = ( ~x26 & n13950 ) | ( ~x26 & n13952 ) | ( n13950 & n13952 ) ;
  assign n13954 = x26 & ~n13952 ;
  assign n13955 = ( ~n13951 & n13953 ) | ( ~n13951 & n13954 ) | ( n13953 & n13954 ) ;
  assign n13956 = ( ~n13798 & n13945 ) | ( ~n13798 & n13955 ) | ( n13945 & n13955 ) ;
  assign n13957 = ( n13798 & n13945 ) | ( n13798 & n13955 ) | ( n13945 & n13955 ) ;
  assign n13958 = ( n13798 & n13956 ) | ( n13798 & ~n13957 ) | ( n13956 & ~n13957 ) ;
  assign n13959 = ( ~n13800 & n13891 ) | ( ~n13800 & n13958 ) | ( n13891 & n13958 ) ;
  assign n13960 = ( n13800 & n13891 ) | ( n13800 & n13958 ) | ( n13891 & n13958 ) ;
  assign n13961 = ( n13800 & n13959 ) | ( n13800 & ~n13960 ) | ( n13959 & ~n13960 ) ;
  assign n13962 = ( ~n13804 & n13881 ) | ( ~n13804 & n13961 ) | ( n13881 & n13961 ) ;
  assign n13963 = ( n13804 & n13881 ) | ( n13804 & n13961 ) | ( n13881 & n13961 ) ;
  assign n13964 = ( n13804 & n13962 ) | ( n13804 & ~n13963 ) | ( n13962 & ~n13963 ) ;
  assign n13965 = ( ~n13806 & n13871 ) | ( ~n13806 & n13964 ) | ( n13871 & n13964 ) ;
  assign n13966 = ( n13806 & n13871 ) | ( n13806 & n13964 ) | ( n13871 & n13964 ) ;
  assign n13967 = ( n13806 & n13965 ) | ( n13806 & ~n13966 ) | ( n13965 & ~n13966 ) ;
  assign n13968 = ( n13810 & n13861 ) | ( n13810 & n13967 ) | ( n13861 & n13967 ) ;
  assign n13969 = ( ~n13810 & n13861 ) | ( ~n13810 & n13967 ) | ( n13861 & n13967 ) ;
  assign n13970 = ( n13810 & ~n13968 ) | ( n13810 & n13969 ) | ( ~n13968 & n13969 ) ;
  assign n13971 = ( n13813 & ~n13851 ) | ( n13813 & n13970 ) | ( ~n13851 & n13970 ) ;
  assign n13972 = ( n13813 & n13851 ) | ( n13813 & n13970 ) | ( n13851 & n13970 ) ;
  assign n13973 = ( n13851 & n13971 ) | ( n13851 & ~n13972 ) | ( n13971 & ~n13972 ) ;
  assign n13974 = ( ~n13816 & n13841 ) | ( ~n13816 & n13973 ) | ( n13841 & n13973 ) ;
  assign n13975 = ( n13816 & n13841 ) | ( n13816 & n13973 ) | ( n13841 & n13973 ) ;
  assign n13976 = ( n13816 & n13974 ) | ( n13816 & ~n13975 ) | ( n13974 & ~n13975 ) ;
  assign n13977 = ( ~n13818 & n13831 ) | ( ~n13818 & n13976 ) | ( n13831 & n13976 ) ;
  assign n13978 = ( n13818 & n13831 ) | ( n13818 & n13976 ) | ( n13831 & n13976 ) ;
  assign n13979 = ( n13818 & n13977 ) | ( n13818 & ~n13978 ) | ( n13977 & ~n13978 ) ;
  assign n13980 = ~x1 & n13476 ;
  assign n13981 = ( n9155 & ~n9158 ) | ( n9155 & n9588 ) | ( ~n9158 & n9588 ) ;
  assign n13982 = n13475 | n13981 ;
  assign n13983 = ~x2 & n9154 ;
  assign n13984 = ( ~n9155 & n13473 ) | ( ~n9155 & n13983 ) | ( n13473 & n13983 ) ;
  assign n13985 = n13475 & ~n13984 ;
  assign n13986 = ( n13980 & n13982 ) | ( n13980 & ~n13985 ) | ( n13982 & ~n13985 ) ;
  assign n13987 = n12325 & n13986 ;
  assign n13988 = n9158 & n13476 ;
  assign n13989 = n13987 & ~n13988 ;
  assign n13990 = ( ~n13821 & n13979 ) | ( ~n13821 & n13989 ) | ( n13979 & n13989 ) ;
  assign n13991 = ( n13821 & n13979 ) | ( n13821 & n13989 ) | ( n13979 & n13989 ) ;
  assign n13992 = ( n13821 & n13990 ) | ( n13821 & ~n13991 ) | ( n13990 & ~n13991 ) ;
  assign n13993 = n40 & n13992 ;
  assign n13994 = x5 & n13993 ;
  assign n13995 = ( ~n13670 & n13680 ) | ( ~n13670 & n13820 ) | ( n13680 & n13820 ) ;
  assign n13996 = ( n13670 & ~n13821 ) | ( n13670 & n13995 ) | ( ~n13821 & n13995 ) ;
  assign n13997 = ( ~n13463 & n13489 ) | ( ~n13463 & n13669 ) | ( n13489 & n13669 ) ;
  assign n13998 = ( n13463 & ~n13670 ) | ( n13463 & n13997 ) | ( ~n13670 & n13997 ) ;
  assign n13999 = ( n13266 & ~n13296 ) | ( n13266 & n13462 ) | ( ~n13296 & n13462 ) ;
  assign n14000 = ( ~n13266 & n13463 ) | ( ~n13266 & n13999 ) | ( n13463 & n13999 ) ;
  assign n14001 = ( ~n12948 & n12961 ) | ( ~n12948 & n13102 ) | ( n12961 & n13102 ) ;
  assign n14002 = ( n12948 & ~n13103 ) | ( n12948 & n14001 ) | ( ~n13103 & n14001 ) ;
  assign n14003 = ( n12752 & ~n12766 ) | ( n12752 & n12947 ) | ( ~n12766 & n12947 ) ;
  assign n14004 = ( ~n12752 & n12948 ) | ( ~n12752 & n14003 ) | ( n12948 & n14003 ) ;
  assign n14005 = n14002 & ~n14004 ;
  assign n14006 = ( n10379 & ~n13103 ) | ( n10379 & n13265 ) | ( ~n13103 & n13265 ) ;
  assign n14007 = ( ~n10379 & n13266 ) | ( ~n10379 & n14006 ) | ( n13266 & n14006 ) ;
  assign n14008 = ~n14005 & n14007 ;
  assign n14009 = n14000 | n14008 ;
  assign n14010 = ~n13998 & n14009 ;
  assign n14011 = n13996 & ~n14010 ;
  assign n14012 = n13992 & n14011 ;
  assign n14013 = ( n10394 & ~n12588 ) | ( n10394 & n12751 ) | ( ~n12588 & n12751 ) ;
  assign n14014 = ( ~n10394 & n12752 ) | ( ~n10394 & n14013 ) | ( n12752 & n14013 ) ;
  assign n14015 = ~n14004 & n14014 ;
  assign n14016 = ~n14002 & n14015 ;
  assign n14017 = ( ~n14002 & n14004 ) | ( ~n14002 & n14016 ) | ( n14004 & n14016 ) ;
  assign n14018 = n14007 | n14017 ;
  assign n14019 = n14000 & n14018 ;
  assign n14020 = n13998 & ~n14019 ;
  assign n14021 = n13996 | n14020 ;
  assign n14022 = ( n13992 & ~n14011 ) | ( n13992 & n14021 ) | ( ~n14011 & n14021 ) ;
  assign n14023 = n13992 & n14021 ;
  assign n14024 = ( n14012 & n14022 ) | ( n14012 & ~n14023 ) | ( n14022 & ~n14023 ) ;
  assign n14025 = n8721 & n13996 ;
  assign n14026 = n8340 & n13998 ;
  assign n14027 = n14025 | n14026 ;
  assign n14028 = n8341 | n14027 ;
  assign n14029 = ( n14024 & n14027 ) | ( n14024 & n14028 ) | ( n14027 & n14028 ) ;
  assign n14030 = x5 & ~n14029 ;
  assign n14031 = ( ~x5 & n13993 ) | ( ~x5 & n14029 ) | ( n13993 & n14029 ) ;
  assign n14032 = ( ~n13994 & n14030 ) | ( ~n13994 & n14031 ) | ( n14030 & n14031 ) ;
  assign n14033 = n40 & ~n14000 ;
  assign n14034 = n8721 & ~n14007 ;
  assign n14035 = n8340 & n14002 ;
  assign n14036 = n14034 | n14035 ;
  assign n14037 = n14033 | n14036 ;
  assign n14038 = x5 & n14037 ;
  assign n14039 = ~n14009 & n14018 ;
  assign n14040 = n14005 & n14007 ;
  assign n14041 = ( ~n14007 & n14019 ) | ( ~n14007 & n14040 ) | ( n14019 & n14040 ) ;
  assign n14042 = ( n14000 & n14039 ) | ( n14000 & ~n14041 ) | ( n14039 & ~n14041 ) ;
  assign n14043 = n8341 & ~n14042 ;
  assign n14044 = ( ~x5 & n14037 ) | ( ~x5 & n14043 ) | ( n14037 & n14043 ) ;
  assign n14045 = x5 & ~n14043 ;
  assign n14046 = ( ~n14038 & n14044 ) | ( ~n14038 & n14045 ) | ( n14044 & n14045 ) ;
  assign n14047 = ( n7644 & n8768 ) | ( n7644 & n14004 ) | ( n8768 & n14004 ) ;
  assign n14048 = ~n14014 & n14047 ;
  assign n14049 = n7342 & n14015 ;
  assign n14050 = n14048 | n14049 ;
  assign n14051 = n7345 & ~n14004 ;
  assign n14052 = n14050 | n14051 ;
  assign n14053 = n7342 & ~n14014 ;
  assign n14054 = x8 & n14053 ;
  assign n14055 = ~n14052 & n14054 ;
  assign n14056 = n14052 & ~n14054 ;
  assign n14057 = n14055 | n14056 ;
  assign n14058 = n40 & ~n14007 ;
  assign n14059 = n8721 & n14002 ;
  assign n14060 = n8340 & ~n14004 ;
  assign n14061 = n14059 | n14060 ;
  assign n14062 = n14058 | n14061 ;
  assign n14063 = x5 & n14062 ;
  assign n14064 = n14007 & ~n14017 ;
  assign n14065 = ( n14005 & ~n14007 ) | ( n14005 & n14017 ) | ( ~n14007 & n14017 ) ;
  assign n14066 = ( ~n14040 & n14064 ) | ( ~n14040 & n14065 ) | ( n14064 & n14065 ) ;
  assign n14067 = n8341 & n14066 ;
  assign n14068 = ( ~x5 & n14062 ) | ( ~x5 & n14067 ) | ( n14062 & n14067 ) ;
  assign n14069 = x5 & ~n14067 ;
  assign n14070 = ( ~n14063 & n14068 ) | ( ~n14063 & n14069 ) | ( n14068 & n14069 ) ;
  assign n14071 = n14002 & ~n14015 ;
  assign n14072 = n14016 | n14071 ;
  assign n14073 = n8341 & n14072 ;
  assign n14074 = n40 & n14002 ;
  assign n14075 = n8721 & ~n14004 ;
  assign n14076 = n8340 & ~n14014 ;
  assign n14077 = n14075 | n14076 ;
  assign n14078 = n14074 | n14077 ;
  assign n14079 = n14073 | n14078 ;
  assign n14080 = ( n8721 & n11802 ) | ( n8721 & n14004 ) | ( n11802 & n14004 ) ;
  assign n14081 = ~n14014 & n14080 ;
  assign n14082 = ( n36 & n40 ) | ( n36 & n14014 ) | ( n40 & n14014 ) ;
  assign n14083 = ~n14004 & n14082 ;
  assign n14084 = n14081 | n14083 ;
  assign n14085 = n11808 & ~n14014 ;
  assign n14086 = ( x5 & n14084 ) | ( x5 & n14085 ) | ( n14084 & n14085 ) ;
  assign n14087 = n14079 | n14086 ;
  assign n14088 = x5 & ~n14087 ;
  assign n14089 = ( n14053 & n14070 ) | ( n14053 & ~n14088 ) | ( n14070 & ~n14088 ) ;
  assign n14090 = n14053 & ~n14088 ;
  assign n14091 = ( n14053 & ~n14070 ) | ( n14053 & n14088 ) | ( ~n14070 & n14088 ) ;
  assign n14092 = ( n14089 & ~n14090 ) | ( n14089 & n14091 ) | ( ~n14090 & n14091 ) ;
  assign n14093 = ( n14053 & n14070 ) | ( n14053 & ~n14092 ) | ( n14070 & ~n14092 ) ;
  assign n14094 = ( n14046 & n14057 ) | ( n14046 & n14093 ) | ( n14057 & n14093 ) ;
  assign n14095 = n7644 & ~n14004 ;
  assign n14096 = n7341 & ~n14014 ;
  assign n14097 = n14095 | n14096 ;
  assign n14098 = n7346 | n14097 ;
  assign n14099 = ( n14072 & n14097 ) | ( n14072 & n14098 ) | ( n14097 & n14098 ) ;
  assign n14100 = n7345 & n14002 ;
  assign n14101 = n14099 | n14100 ;
  assign n14102 = ~x8 & n14101 ;
  assign n14103 = n14052 | n14053 ;
  assign n14104 = ( x8 & n14101 ) | ( x8 & n14103 ) | ( n14101 & n14103 ) ;
  assign n14105 = n14101 & n14103 ;
  assign n14106 = ( n14102 & n14104 ) | ( n14102 & ~n14105 ) | ( n14104 & ~n14105 ) ;
  assign n14107 = n40 & n13998 ;
  assign n14108 = n8721 & ~n14000 ;
  assign n14109 = n8340 & ~n14007 ;
  assign n14110 = n14108 | n14109 ;
  assign n14111 = n14107 | n14110 ;
  assign n14112 = x5 & n14111 ;
  assign n14113 = n13998 & ~n14009 ;
  assign n14114 = ( n13998 & n14009 ) | ( n13998 & ~n14019 ) | ( n14009 & ~n14019 ) ;
  assign n14115 = ( ~n14020 & n14113 ) | ( ~n14020 & n14114 ) | ( n14113 & n14114 ) ;
  assign n14116 = n8341 & n14115 ;
  assign n14117 = ( ~x5 & n14111 ) | ( ~x5 & n14116 ) | ( n14111 & n14116 ) ;
  assign n14118 = x5 & ~n14116 ;
  assign n14119 = ( ~n14112 & n14117 ) | ( ~n14112 & n14118 ) | ( n14117 & n14118 ) ;
  assign n14120 = ( n14094 & n14106 ) | ( n14094 & n14119 ) | ( n14106 & n14119 ) ;
  assign n14121 = n40 & n13996 ;
  assign n14122 = n8721 & n13998 ;
  assign n14123 = n8340 & ~n14000 ;
  assign n14124 = n14122 | n14123 ;
  assign n14125 = n14121 | n14124 ;
  assign n14126 = x5 & n14125 ;
  assign n14127 = ( ~n13996 & n14010 ) | ( ~n13996 & n14020 ) | ( n14010 & n14020 ) ;
  assign n14128 = n13996 & ~n14020 ;
  assign n14129 = ( n13996 & n14010 ) | ( n13996 & n14020 ) | ( n14010 & n14020 ) ;
  assign n14130 = ( n14127 & n14128 ) | ( n14127 & ~n14129 ) | ( n14128 & ~n14129 ) ;
  assign n14131 = n8341 & ~n14130 ;
  assign n14132 = ( ~x5 & n14125 ) | ( ~x5 & n14131 ) | ( n14125 & n14131 ) ;
  assign n14133 = x5 & ~n14131 ;
  assign n14134 = ( ~n14126 & n14132 ) | ( ~n14126 & n14133 ) | ( n14132 & n14133 ) ;
  assign n14135 = x8 & ~n14103 ;
  assign n14136 = ~n14101 & n14135 ;
  assign n14137 = n6568 & ~n14014 ;
  assign n14138 = n7644 & n14002 ;
  assign n14139 = x8 & n14138 ;
  assign n14140 = n7341 & ~n14004 ;
  assign n14141 = n7345 | n14140 ;
  assign n14142 = ( ~n14007 & n14140 ) | ( ~n14007 & n14141 ) | ( n14140 & n14141 ) ;
  assign n14143 = n7346 | n14142 ;
  assign n14144 = ( n14066 & n14142 ) | ( n14066 & n14143 ) | ( n14142 & n14143 ) ;
  assign n14145 = x8 & ~n14144 ;
  assign n14146 = ( ~x8 & n14138 ) | ( ~x8 & n14144 ) | ( n14138 & n14144 ) ;
  assign n14147 = ( ~n14139 & n14145 ) | ( ~n14139 & n14146 ) | ( n14145 & n14146 ) ;
  assign n14148 = ( n14136 & ~n14137 ) | ( n14136 & n14147 ) | ( ~n14137 & n14147 ) ;
  assign n14149 = n14136 & ~n14137 ;
  assign n14150 = ( n14136 & n14137 ) | ( n14136 & ~n14147 ) | ( n14137 & ~n14147 ) ;
  assign n14151 = ( n14148 & ~n14149 ) | ( n14148 & n14150 ) | ( ~n14149 & n14150 ) ;
  assign n14152 = ( n14120 & n14134 ) | ( n14120 & n14151 ) | ( n14134 & n14151 ) ;
  assign n14153 = n7644 & ~n14007 ;
  assign n14154 = x8 & n14153 ;
  assign n14155 = n7341 & n14002 ;
  assign n14156 = n7345 | n14155 ;
  assign n14157 = ( ~n14000 & n14155 ) | ( ~n14000 & n14156 ) | ( n14155 & n14156 ) ;
  assign n14158 = n7346 | n14157 ;
  assign n14159 = ( ~n14042 & n14157 ) | ( ~n14042 & n14158 ) | ( n14157 & n14158 ) ;
  assign n14160 = x8 & ~n14159 ;
  assign n14161 = ( ~x8 & n14153 ) | ( ~x8 & n14159 ) | ( n14153 & n14159 ) ;
  assign n14162 = ( ~n14154 & n14160 ) | ( ~n14154 & n14161 ) | ( n14160 & n14161 ) ;
  assign n14163 = n6571 & n14004 ;
  assign n14164 = n6796 & ~n14014 ;
  assign n14165 = ( ~n14014 & n14163 ) | ( ~n14014 & n14164 ) | ( n14163 & n14164 ) ;
  assign n14166 = ( n6568 & n6570 ) | ( n6568 & n14014 ) | ( n6570 & n14014 ) ;
  assign n14167 = ~n14004 & n14166 ;
  assign n14168 = n14165 | n14167 ;
  assign n14169 = x11 & n14137 ;
  assign n14170 = ~n14168 & n14169 ;
  assign n14171 = n14168 & ~n14169 ;
  assign n14172 = n14170 | n14171 ;
  assign n14173 = ( n14137 & n14147 ) | ( n14137 & ~n14151 ) | ( n14147 & ~n14151 ) ;
  assign n14174 = ( n14162 & n14172 ) | ( n14162 & n14173 ) | ( n14172 & n14173 ) ;
  assign n14175 = ( ~n14162 & n14172 ) | ( ~n14162 & n14173 ) | ( n14172 & n14173 ) ;
  assign n14176 = ( n14162 & ~n14174 ) | ( n14162 & n14175 ) | ( ~n14174 & n14175 ) ;
  assign n14177 = ( n14032 & n14152 ) | ( n14032 & n14176 ) | ( n14152 & n14176 ) ;
  assign n14178 = n7644 & ~n14000 ;
  assign n14179 = x8 & n14178 ;
  assign n14180 = n7341 & ~n14007 ;
  assign n14181 = n7345 | n14180 ;
  assign n14182 = ( n13998 & n14180 ) | ( n13998 & n14181 ) | ( n14180 & n14181 ) ;
  assign n14183 = n7346 | n14182 ;
  assign n14184 = ( n14115 & n14182 ) | ( n14115 & n14183 ) | ( n14182 & n14183 ) ;
  assign n14185 = x8 & ~n14184 ;
  assign n14186 = ( ~x8 & n14178 ) | ( ~x8 & n14184 ) | ( n14178 & n14184 ) ;
  assign n14187 = ( ~n14179 & n14185 ) | ( ~n14179 & n14186 ) | ( n14185 & n14186 ) ;
  assign n14188 = x11 & ~n14137 ;
  assign n14189 = ~n14168 & n14188 ;
  assign n14190 = x11 & ~n14189 ;
  assign n14191 = n6796 & ~n14004 ;
  assign n14192 = n6567 & ~n14014 ;
  assign n14193 = n14191 | n14192 ;
  assign n14194 = n6571 | n14193 ;
  assign n14195 = ( n14072 & n14193 ) | ( n14072 & n14194 ) | ( n14193 & n14194 ) ;
  assign n14196 = n6570 & n14002 ;
  assign n14197 = n14195 | n14196 ;
  assign n14198 = n14190 & ~n14197 ;
  assign n14199 = ~n14190 & n14197 ;
  assign n14200 = n14198 | n14199 ;
  assign n14201 = ( n14174 & ~n14187 ) | ( n14174 & n14200 ) | ( ~n14187 & n14200 ) ;
  assign n14202 = ( n14174 & n14187 ) | ( n14174 & n14200 ) | ( n14187 & n14200 ) ;
  assign n14203 = ( n14187 & n14201 ) | ( n14187 & ~n14202 ) | ( n14201 & ~n14202 ) ;
  assign n14204 = n9600 | n13983 ;
  assign n14205 = ( ~n13475 & n13983 ) | ( ~n13475 & n14204 ) | ( n13983 & n14204 ) ;
  assign n14206 = n40 & ~n13473 ;
  assign n14207 = n8340 & ~n10235 ;
  assign n14208 = n14206 | n14207 ;
  assign n14209 = n8721 & ~n13280 ;
  assign n14210 = n14208 | n14209 ;
  assign n14211 = n8341 | n14210 ;
  assign n14212 = ( ~n13480 & n14210 ) | ( ~n13480 & n14211 ) | ( n14210 & n14211 ) ;
  assign n14213 = x5 & ~n14212 ;
  assign n14214 = ~x5 & n14212 ;
  assign n14215 = n14213 | n14214 ;
  assign n14216 = n7644 & ~n10237 ;
  assign n14217 = x8 & n14216 ;
  assign n14218 = n7341 & ~n10332 ;
  assign n14219 = n7345 | n14218 ;
  assign n14220 = ( n10214 & n14218 ) | ( n10214 & n14219 ) | ( n14218 & n14219 ) ;
  assign n14221 = n7346 | n14220 ;
  assign n14222 = ( n12953 & n14220 ) | ( n12953 & n14221 ) | ( n14220 & n14221 ) ;
  assign n14223 = x8 & ~n14222 ;
  assign n14224 = ( ~x8 & n14216 ) | ( ~x8 & n14222 ) | ( n14216 & n14222 ) ;
  assign n14225 = ( ~n14217 & n14223 ) | ( ~n14217 & n14224 ) | ( n14223 & n14224 ) ;
  assign n14226 = n6571 & n10397 ;
  assign n14227 = x11 & n14226 ;
  assign n14228 = n6567 & n10239 ;
  assign n14229 = n6570 | n14228 ;
  assign n14230 = ( n10329 & n14228 ) | ( n10329 & n14229 ) | ( n14228 & n14229 ) ;
  assign n14231 = n6796 & n10326 ;
  assign n14232 = n14230 | n14231 ;
  assign n14233 = x11 & ~n14232 ;
  assign n14234 = ( ~x11 & n14226 ) | ( ~x11 & n14232 ) | ( n14226 & n14232 ) ;
  assign n14235 = ( ~n14227 & n14233 ) | ( ~n14227 & n14234 ) | ( n14233 & n14234 ) ;
  assign n14236 = n6332 & n10243 ;
  assign n14237 = x14 & n14236 ;
  assign n14238 = n5909 & ~n10320 ;
  assign n14239 = n5914 | n14238 ;
  assign n14240 = ( n10241 & n14238 ) | ( n10241 & n14239 ) | ( n14238 & n14239 ) ;
  assign n14241 = n5915 | n14240 ;
  assign n14242 = ( n12105 & n14240 ) | ( n12105 & n14241 ) | ( n14240 & n14241 ) ;
  assign n14243 = x14 & ~n14242 ;
  assign n14244 = ( ~x14 & n14236 ) | ( ~x14 & n14242 ) | ( n14236 & n14242 ) ;
  assign n14245 = ( ~n14237 & n14243 ) | ( ~n14237 & n14244 ) | ( n14243 & n14244 ) ;
  assign n14246 = n5584 & ~n10316 ;
  assign n14247 = x17 & n14246 ;
  assign n14248 = n5413 & n10247 ;
  assign n14249 = n5417 | n14248 ;
  assign n14250 = ( n10245 & n14248 ) | ( n10245 & n14249 ) | ( n14248 & n14249 ) ;
  assign n14251 = n5418 | n14250 ;
  assign n14252 = ( ~n11676 & n14250 ) | ( ~n11676 & n14251 ) | ( n14250 & n14251 ) ;
  assign n14253 = x17 & ~n14252 ;
  assign n14254 = ( ~x17 & n14246 ) | ( ~x17 & n14252 ) | ( n14246 & n14252 ) ;
  assign n14255 = ( ~n14247 & n14253 ) | ( ~n14247 & n14254 ) | ( n14253 & n14254 ) ;
  assign n14256 = n4878 & n10312 ;
  assign n14257 = n5232 & ~n10249 ;
  assign n14258 = n4874 & n10251 ;
  assign n14259 = n14257 | n14258 ;
  assign n14260 = n14256 | n14259 ;
  assign n14261 = x20 & n14260 ;
  assign n14262 = n4879 & ~n11486 ;
  assign n14263 = x20 & ~n14262 ;
  assign n14264 = ( ~x20 & n14260 ) | ( ~x20 & n14262 ) | ( n14260 & n14262 ) ;
  assign n14265 = ( ~n14261 & n14263 ) | ( ~n14261 & n14264 ) | ( n14263 & n14264 ) ;
  assign n14266 = n4637 & n10255 ;
  assign n14267 = x23 & n14266 ;
  assign n14268 = n4584 & n10257 ;
  assign n14269 = n4649 | n14268 ;
  assign n14270 = ( ~n10253 & n14268 ) | ( ~n10253 & n14269 ) | ( n14268 & n14269 ) ;
  assign n14271 = n4591 | n14270 ;
  assign n14272 = ( ~n11297 & n14270 ) | ( ~n11297 & n14271 ) | ( n14270 & n14271 ) ;
  assign n14273 = x23 & ~n14272 ;
  assign n14274 = ( ~x23 & n14266 ) | ( ~x23 & n14272 ) | ( n14266 & n14272 ) ;
  assign n14275 = ( ~n14267 & n14273 ) | ( ~n14267 & n14274 ) | ( n14273 & n14274 ) ;
  assign n14276 = n3541 & n10804 ;
  assign n14277 = x29 & n14276 ;
  assign n14278 = n3536 & ~n10269 ;
  assign n14279 = n4039 | n14278 ;
  assign n14280 = ( n10265 & n14278 ) | ( n10265 & n14279 ) | ( n14278 & n14279 ) ;
  assign n14281 = n3501 & n10267 ;
  assign n14282 = n14280 | n14281 ;
  assign n14283 = x29 & ~n14282 ;
  assign n14284 = ( ~x29 & n14276 ) | ( ~x29 & n14282 ) | ( n14276 & n14282 ) ;
  assign n14285 = ( ~n14277 & n14283 ) | ( ~n14277 & n14284 ) | ( n14283 & n14284 ) ;
  assign n14286 = n3273 & n10273 ;
  assign n14287 = n3270 | n14286 ;
  assign n14288 = ( n10271 & n14286 ) | ( n10271 & n14287 ) | ( n14286 & n14287 ) ;
  assign n14289 = n390 | n14288 ;
  assign n14290 = ( ~n10656 & n14288 ) | ( ~n10656 & n14289 ) | ( n14288 & n14289 ) ;
  assign n14291 = n3274 & ~n10297 ;
  assign n14292 = n14290 | n14291 ;
  assign n14293 = n2831 | n5674 ;
  assign n14294 = n87 | n150 ;
  assign n14295 = n1012 | n14294 ;
  assign n14296 = n131 | n378 ;
  assign n14297 = n265 | n374 ;
  assign n14298 = n14296 | n14297 ;
  assign n14299 = n450 | n1780 ;
  assign n14300 = n14298 | n14299 ;
  assign n14301 = n14295 | n14300 ;
  assign n14302 = n3000 | n3992 ;
  assign n14303 = n635 | n1126 ;
  assign n14304 = n14302 | n14303 ;
  assign n14305 = n14301 | n14304 ;
  assign n14306 = n14293 | n14305 ;
  assign n14307 = n3653 | n14306 ;
  assign n14308 = n1315 | n1625 ;
  assign n14309 = n14307 | n14308 ;
  assign n14310 = ( n13940 & n14292 ) | ( n13940 & n14309 ) | ( n14292 & n14309 ) ;
  assign n14311 = ( ~n13940 & n14292 ) | ( ~n13940 & n14309 ) | ( n14292 & n14309 ) ;
  assign n14312 = ( n13940 & ~n14310 ) | ( n13940 & n14311 ) | ( ~n14310 & n14311 ) ;
  assign n14313 = ( ~n13944 & n14285 ) | ( ~n13944 & n14312 ) | ( n14285 & n14312 ) ;
  assign n14314 = ( n13944 & n14285 ) | ( n13944 & n14312 ) | ( n14285 & n14312 ) ;
  assign n14315 = ( n13944 & n14313 ) | ( n13944 & ~n14314 ) | ( n14313 & ~n14314 ) ;
  assign n14316 = n4215 & n10259 ;
  assign n14317 = n4200 & n10261 ;
  assign n14318 = n2083 & n10263 ;
  assign n14319 = n14317 | n14318 ;
  assign n14320 = n14316 | n14319 ;
  assign n14321 = x26 & n14320 ;
  assign n14322 = n4203 & n10859 ;
  assign n14323 = ( ~x26 & n14320 ) | ( ~x26 & n14322 ) | ( n14320 & n14322 ) ;
  assign n14324 = x26 & ~n14322 ;
  assign n14325 = ( ~n14321 & n14323 ) | ( ~n14321 & n14324 ) | ( n14323 & n14324 ) ;
  assign n14326 = ( ~n13957 & n14315 ) | ( ~n13957 & n14325 ) | ( n14315 & n14325 ) ;
  assign n14327 = ( n13957 & n14315 ) | ( n13957 & n14325 ) | ( n14315 & n14325 ) ;
  assign n14328 = ( n13957 & n14326 ) | ( n13957 & ~n14327 ) | ( n14326 & ~n14327 ) ;
  assign n14329 = ( ~n13960 & n14275 ) | ( ~n13960 & n14328 ) | ( n14275 & n14328 ) ;
  assign n14330 = ( n13960 & n14275 ) | ( n13960 & n14328 ) | ( n14275 & n14328 ) ;
  assign n14331 = ( n13960 & n14329 ) | ( n13960 & ~n14330 ) | ( n14329 & ~n14330 ) ;
  assign n14332 = ( ~n13963 & n14265 ) | ( ~n13963 & n14331 ) | ( n14265 & n14331 ) ;
  assign n14333 = ( n13963 & n14265 ) | ( n13963 & n14331 ) | ( n14265 & n14331 ) ;
  assign n14334 = ( n13963 & n14332 ) | ( n13963 & ~n14333 ) | ( n14332 & ~n14333 ) ;
  assign n14335 = ( ~n13966 & n14255 ) | ( ~n13966 & n14334 ) | ( n14255 & n14334 ) ;
  assign n14336 = ( n13966 & n14255 ) | ( n13966 & n14334 ) | ( n14255 & n14334 ) ;
  assign n14337 = ( n13966 & n14335 ) | ( n13966 & ~n14336 ) | ( n14335 & ~n14336 ) ;
  assign n14338 = ( ~n13968 & n14245 ) | ( ~n13968 & n14337 ) | ( n14245 & n14337 ) ;
  assign n14339 = ( n13968 & n14245 ) | ( n13968 & n14337 ) | ( n14245 & n14337 ) ;
  assign n14340 = ( n13968 & n14338 ) | ( n13968 & ~n14339 ) | ( n14338 & ~n14339 ) ;
  assign n14341 = ( ~n13972 & n14235 ) | ( ~n13972 & n14340 ) | ( n14235 & n14340 ) ;
  assign n14342 = ( n13972 & n14235 ) | ( n13972 & n14340 ) | ( n14235 & n14340 ) ;
  assign n14343 = ( n13972 & n14341 ) | ( n13972 & ~n14342 ) | ( n14341 & ~n14342 ) ;
  assign n14344 = ( n13975 & ~n14225 ) | ( n13975 & n14343 ) | ( ~n14225 & n14343 ) ;
  assign n14345 = ( n13975 & n14225 ) | ( n13975 & n14343 ) | ( n14225 & n14343 ) ;
  assign n14346 = ( n14225 & n14344 ) | ( n14225 & ~n14345 ) | ( n14344 & ~n14345 ) ;
  assign n14347 = ( ~n13978 & n14215 ) | ( ~n13978 & n14346 ) | ( n14215 & n14346 ) ;
  assign n14348 = ( n13978 & n14215 ) | ( n13978 & n14346 ) | ( n14215 & n14346 ) ;
  assign n14349 = ( n13978 & n14347 ) | ( n13978 & ~n14348 ) | ( n14347 & ~n14348 ) ;
  assign n14350 = ( ~n13991 & n14205 ) | ( ~n13991 & n14349 ) | ( n14205 & n14349 ) ;
  assign n14351 = ( n13991 & n14205 ) | ( n13991 & n14349 ) | ( n14205 & n14349 ) ;
  assign n14352 = ( n13991 & n14350 ) | ( n13991 & ~n14351 ) | ( n14350 & ~n14351 ) ;
  assign n14353 = n40 & n14352 ;
  assign n14354 = n8721 & n13992 ;
  assign n14355 = n8340 & n13996 ;
  assign n14356 = n14354 | n14355 ;
  assign n14357 = n14353 | n14356 ;
  assign n14358 = x5 & n14357 ;
  assign n14359 = n13992 | n14011 ;
  assign n14360 = n14352 | n14359 ;
  assign n14361 = ( n14023 & n14352 ) | ( n14023 & ~n14359 ) | ( n14352 & ~n14359 ) ;
  assign n14362 = n14023 | n14352 ;
  assign n14363 = ( n14360 & n14361 ) | ( n14360 & ~n14362 ) | ( n14361 & ~n14362 ) ;
  assign n14364 = n8341 & n14363 ;
  assign n14365 = ( ~x5 & n14357 ) | ( ~x5 & n14364 ) | ( n14357 & n14364 ) ;
  assign n14366 = x5 & ~n14364 ;
  assign n14367 = ( ~n14358 & n14365 ) | ( ~n14358 & n14366 ) | ( n14365 & n14366 ) ;
  assign n14368 = ( n14177 & n14203 ) | ( n14177 & n14367 ) | ( n14203 & n14367 ) ;
  assign n14369 = n8721 & ~n13473 ;
  assign n14370 = n40 | n14369 ;
  assign n14371 = ( n13475 & n14369 ) | ( n13475 & n14370 ) | ( n14369 & n14370 ) ;
  assign n14372 = n8340 & ~n13280 ;
  assign n14373 = n14371 | n14372 ;
  assign n14374 = x5 & n14373 ;
  assign n14375 = n8341 & n13671 ;
  assign n14376 = ( ~x5 & n14373 ) | ( ~x5 & n14375 ) | ( n14373 & n14375 ) ;
  assign n14377 = x5 & ~n14375 ;
  assign n14378 = ( ~n14374 & n14376 ) | ( ~n14374 & n14377 ) | ( n14376 & n14377 ) ;
  assign n14379 = n7644 & n10214 ;
  assign n14380 = x8 & n14379 ;
  assign n14381 = n7341 & ~n10237 ;
  assign n14382 = n7345 | n14381 ;
  assign n14383 = ( ~n10235 & n14381 ) | ( ~n10235 & n14382 ) | ( n14381 & n14382 ) ;
  assign n14384 = n7346 | n14383 ;
  assign n14385 = ( n10371 & n14383 ) | ( n10371 & n14384 ) | ( n14383 & n14384 ) ;
  assign n14386 = x8 & ~n14385 ;
  assign n14387 = ( ~x8 & n14379 ) | ( ~x8 & n14385 ) | ( n14379 & n14385 ) ;
  assign n14388 = ( ~n14380 & n14386 ) | ( ~n14380 & n14387 ) | ( n14386 & n14387 ) ;
  assign n14389 = n5915 & n12575 ;
  assign n14390 = x14 & n14389 ;
  assign n14391 = n5909 & n10243 ;
  assign n14392 = n5914 | n14391 ;
  assign n14393 = ( n10239 & n14391 ) | ( n10239 & n14392 ) | ( n14391 & n14392 ) ;
  assign n14394 = n6332 & n10241 ;
  assign n14395 = n14393 | n14394 ;
  assign n14396 = x14 & ~n14395 ;
  assign n14397 = ( ~x14 & n14389 ) | ( ~x14 & n14395 ) | ( n14389 & n14395 ) ;
  assign n14398 = ( ~n14390 & n14396 ) | ( ~n14390 & n14397 ) | ( n14396 & n14397 ) ;
  assign n14399 = n5417 & ~n10320 ;
  assign n14400 = x17 & n14399 ;
  assign n14401 = n5584 & n10245 ;
  assign n14402 = n5413 & ~n10316 ;
  assign n14403 = n14401 | n14402 ;
  assign n14404 = n5418 | n14403 ;
  assign n14405 = ( ~n10414 & n14403 ) | ( ~n10414 & n14404 ) | ( n14403 & n14404 ) ;
  assign n14406 = x17 & ~n14405 ;
  assign n14407 = ( ~x17 & n14399 ) | ( ~x17 & n14405 ) | ( n14399 & n14405 ) ;
  assign n14408 = ( ~n14400 & n14406 ) | ( ~n14400 & n14407 ) | ( n14406 & n14407 ) ;
  assign n14409 = n5232 & n10312 ;
  assign n14410 = x20 & n14409 ;
  assign n14411 = n4874 & ~n10249 ;
  assign n14412 = n4878 | n14411 ;
  assign n14413 = ( n10247 & n14411 ) | ( n10247 & n14412 ) | ( n14411 & n14412 ) ;
  assign n14414 = n4879 | n14413 ;
  assign n14415 = ( n10428 & n14413 ) | ( n10428 & n14414 ) | ( n14413 & n14414 ) ;
  assign n14416 = x20 & ~n14415 ;
  assign n14417 = ( ~x20 & n14409 ) | ( ~x20 & n14415 ) | ( n14409 & n14415 ) ;
  assign n14418 = ( ~n14410 & n14416 ) | ( ~n14410 & n14417 ) | ( n14416 & n14417 ) ;
  assign n14419 = n4591 & ~n11309 ;
  assign n14420 = x23 & n14419 ;
  assign n14421 = n4584 & n10255 ;
  assign n14422 = n4649 | n14421 ;
  assign n14423 = ( n10251 & n14421 ) | ( n10251 & n14422 ) | ( n14421 & n14422 ) ;
  assign n14424 = n4637 & ~n10253 ;
  assign n14425 = n14423 | n14424 ;
  assign n14426 = x23 & ~n14425 ;
  assign n14427 = ( ~x23 & n14419 ) | ( ~x23 & n14425 ) | ( n14419 & n14425 ) ;
  assign n14428 = ( ~n14420 & n14426 ) | ( ~n14420 & n14427 ) | ( n14426 & n14427 ) ;
  assign n14429 = n3541 & n10874 ;
  assign n14430 = x29 & n14429 ;
  assign n14431 = n3536 & n10267 ;
  assign n14432 = n4039 | n14431 ;
  assign n14433 = ( n10263 & n14431 ) | ( n10263 & n14432 ) | ( n14431 & n14432 ) ;
  assign n14434 = n3501 & n10265 ;
  assign n14435 = n14433 | n14434 ;
  assign n14436 = x29 & ~n14435 ;
  assign n14437 = ( ~x29 & n14429 ) | ( ~x29 & n14435 ) | ( n14429 & n14435 ) ;
  assign n14438 = ( ~n14430 & n14436 ) | ( ~n14430 & n14437 ) | ( n14436 & n14437 ) ;
  assign n14439 = n3273 & ~n10297 ;
  assign n14440 = n3270 | n14439 ;
  assign n14441 = ( ~n10269 & n14439 ) | ( ~n10269 & n14440 ) | ( n14439 & n14440 ) ;
  assign n14442 = n390 | n14441 ;
  assign n14443 = ( ~n10698 & n14441 ) | ( ~n10698 & n14442 ) | ( n14441 & n14442 ) ;
  assign n14444 = n3274 & n10271 ;
  assign n14445 = n14443 | n14444 ;
  assign n14446 = n358 | n1107 ;
  assign n14447 = n975 | n14446 ;
  assign n14448 = n2727 | n14447 ;
  assign n14449 = n2988 | n3167 ;
  assign n14450 = n1056 | n14449 ;
  assign n14451 = n14448 | n14450 ;
  assign n14452 = n593 | n1094 ;
  assign n14453 = n863 | n14452 ;
  assign n14454 = n684 | n1375 ;
  assign n14455 = n14453 | n14454 ;
  assign n14456 = n614 | n3328 ;
  assign n14457 = n191 | n308 ;
  assign n14458 = n751 | n989 ;
  assign n14459 = n14457 | n14458 ;
  assign n14460 = n14456 | n14459 ;
  assign n14461 = n14455 | n14460 ;
  assign n14462 = n14451 | n14461 ;
  assign n14463 = n3186 | n5053 ;
  assign n14464 = n3907 | n14463 ;
  assign n14465 = n14462 | n14464 ;
  assign n14466 = n1369 | n4802 ;
  assign n14467 = n14465 | n14466 ;
  assign n14468 = ( n14310 & n14445 ) | ( n14310 & n14467 ) | ( n14445 & n14467 ) ;
  assign n14469 = ( ~n14310 & n14445 ) | ( ~n14310 & n14467 ) | ( n14445 & n14467 ) ;
  assign n14470 = ( n14310 & ~n14468 ) | ( n14310 & n14469 ) | ( ~n14468 & n14469 ) ;
  assign n14471 = ( n14314 & n14438 ) | ( n14314 & n14470 ) | ( n14438 & n14470 ) ;
  assign n14472 = ( ~n14314 & n14438 ) | ( ~n14314 & n14470 ) | ( n14438 & n14470 ) ;
  assign n14473 = ( n14314 & ~n14471 ) | ( n14314 & n14472 ) | ( ~n14471 & n14472 ) ;
  assign n14474 = n4215 & n10257 ;
  assign n14475 = n4200 & n10259 ;
  assign n14476 = n2083 & n10261 ;
  assign n14477 = n14475 | n14476 ;
  assign n14478 = n14474 | n14477 ;
  assign n14479 = x26 & n14478 ;
  assign n14480 = n4203 & n11065 ;
  assign n14481 = ( ~x26 & n14478 ) | ( ~x26 & n14480 ) | ( n14478 & n14480 ) ;
  assign n14482 = x26 & ~n14480 ;
  assign n14483 = ( ~n14479 & n14481 ) | ( ~n14479 & n14482 ) | ( n14481 & n14482 ) ;
  assign n14484 = ( n14327 & n14473 ) | ( n14327 & n14483 ) | ( n14473 & n14483 ) ;
  assign n14485 = ( ~n14327 & n14473 ) | ( ~n14327 & n14483 ) | ( n14473 & n14483 ) ;
  assign n14486 = ( n14327 & ~n14484 ) | ( n14327 & n14485 ) | ( ~n14484 & n14485 ) ;
  assign n14487 = ( ~n14330 & n14428 ) | ( ~n14330 & n14486 ) | ( n14428 & n14486 ) ;
  assign n14488 = ( n14330 & n14428 ) | ( n14330 & n14486 ) | ( n14428 & n14486 ) ;
  assign n14489 = ( n14330 & n14487 ) | ( n14330 & ~n14488 ) | ( n14487 & ~n14488 ) ;
  assign n14490 = ( n14333 & n14418 ) | ( n14333 & n14489 ) | ( n14418 & n14489 ) ;
  assign n14491 = ( ~n14333 & n14418 ) | ( ~n14333 & n14489 ) | ( n14418 & n14489 ) ;
  assign n14492 = ( n14333 & ~n14490 ) | ( n14333 & n14491 ) | ( ~n14490 & n14491 ) ;
  assign n14493 = ( ~n14336 & n14408 ) | ( ~n14336 & n14492 ) | ( n14408 & n14492 ) ;
  assign n14494 = ( n14336 & n14408 ) | ( n14336 & n14492 ) | ( n14408 & n14492 ) ;
  assign n14495 = ( n14336 & n14493 ) | ( n14336 & ~n14494 ) | ( n14493 & ~n14494 ) ;
  assign n14496 = ( ~n14339 & n14398 ) | ( ~n14339 & n14495 ) | ( n14398 & n14495 ) ;
  assign n14497 = ( n14339 & n14398 ) | ( n14339 & n14495 ) | ( n14398 & n14495 ) ;
  assign n14498 = ( n14339 & n14496 ) | ( n14339 & ~n14497 ) | ( n14496 & ~n14497 ) ;
  assign n14499 = n6796 & n10329 ;
  assign n14500 = x11 & n14499 ;
  assign n14501 = n6567 & n10326 ;
  assign n14502 = n6570 | n14501 ;
  assign n14503 = ( ~n10332 & n14501 ) | ( ~n10332 & n14502 ) | ( n14501 & n14502 ) ;
  assign n14504 = n6571 | n14503 ;
  assign n14505 = ( ~n10383 & n14503 ) | ( ~n10383 & n14504 ) | ( n14503 & n14504 ) ;
  assign n14506 = x11 & ~n14505 ;
  assign n14507 = ( ~x11 & n14499 ) | ( ~x11 & n14505 ) | ( n14499 & n14505 ) ;
  assign n14508 = ( ~n14500 & n14506 ) | ( ~n14500 & n14507 ) | ( n14506 & n14507 ) ;
  assign n14509 = ( ~n14342 & n14498 ) | ( ~n14342 & n14508 ) | ( n14498 & n14508 ) ;
  assign n14510 = ( n14342 & n14498 ) | ( n14342 & n14508 ) | ( n14498 & n14508 ) ;
  assign n14511 = ( n14342 & n14509 ) | ( n14342 & ~n14510 ) | ( n14509 & ~n14510 ) ;
  assign n14512 = ( n14345 & ~n14388 ) | ( n14345 & n14511 ) | ( ~n14388 & n14511 ) ;
  assign n14513 = ( n14345 & n14388 ) | ( n14345 & n14511 ) | ( n14388 & n14511 ) ;
  assign n14514 = ( n14388 & n14512 ) | ( n14388 & ~n14513 ) | ( n14512 & ~n14513 ) ;
  assign n14515 = ( ~n13983 & n14378 ) | ( ~n13983 & n14514 ) | ( n14378 & n14514 ) ;
  assign n14516 = ( n13983 & n14378 ) | ( n13983 & n14514 ) | ( n14378 & n14514 ) ;
  assign n14517 = ( n13983 & n14515 ) | ( n13983 & ~n14516 ) | ( n14515 & ~n14516 ) ;
  assign n14518 = ( n14348 & ~n14351 ) | ( n14348 & n14517 ) | ( ~n14351 & n14517 ) ;
  assign n14519 = ( n14348 & n14351 ) | ( n14348 & n14517 ) | ( n14351 & n14517 ) ;
  assign n14520 = ( n14351 & n14518 ) | ( n14351 & ~n14519 ) | ( n14518 & ~n14519 ) ;
  assign n14521 = n40 & n14520 ;
  assign n14522 = n8721 & n14352 ;
  assign n14523 = n8340 & n13992 ;
  assign n14524 = n14522 | n14523 ;
  assign n14525 = n14521 | n14524 ;
  assign n14526 = x5 & n14525 ;
  assign n14527 = n14352 & n14359 ;
  assign n14528 = n14520 & n14527 ;
  assign n14529 = n14362 & n14520 ;
  assign n14530 = ( n14362 & n14520 ) | ( n14362 & ~n14527 ) | ( n14520 & ~n14527 ) ;
  assign n14531 = ( n14528 & ~n14529 ) | ( n14528 & n14530 ) | ( ~n14529 & n14530 ) ;
  assign n14532 = n8341 & n14531 ;
  assign n14533 = ( ~x5 & n14525 ) | ( ~x5 & n14532 ) | ( n14525 & n14532 ) ;
  assign n14534 = x5 & ~n14532 ;
  assign n14535 = ( ~n14526 & n14533 ) | ( ~n14526 & n14534 ) | ( n14533 & n14534 ) ;
  assign n14536 = n7644 & n13998 ;
  assign n14537 = x8 & n14536 ;
  assign n14538 = n7341 & ~n14000 ;
  assign n14539 = n7345 | n14538 ;
  assign n14540 = ( n13996 & n14538 ) | ( n13996 & n14539 ) | ( n14538 & n14539 ) ;
  assign n14541 = n7346 | n14540 ;
  assign n14542 = ( ~n14130 & n14540 ) | ( ~n14130 & n14541 ) | ( n14540 & n14541 ) ;
  assign n14543 = x8 & ~n14542 ;
  assign n14544 = ( ~x8 & n14536 ) | ( ~x8 & n14542 ) | ( n14536 & n14542 ) ;
  assign n14545 = ( ~n14537 & n14543 ) | ( ~n14537 & n14544 ) | ( n14543 & n14544 ) ;
  assign n14546 = n14189 & ~n14197 ;
  assign n14547 = n6796 & n14002 ;
  assign n14548 = x11 & n14547 ;
  assign n14549 = n6567 & ~n14004 ;
  assign n14550 = n6570 | n14549 ;
  assign n14551 = ( ~n14007 & n14549 ) | ( ~n14007 & n14550 ) | ( n14549 & n14550 ) ;
  assign n14552 = n6571 | n14551 ;
  assign n14553 = ( n14066 & n14551 ) | ( n14066 & n14552 ) | ( n14551 & n14552 ) ;
  assign n14554 = x11 & ~n14553 ;
  assign n14555 = ( ~x11 & n14547 ) | ( ~x11 & n14553 ) | ( n14547 & n14553 ) ;
  assign n14556 = ( ~n14548 & n14554 ) | ( ~n14548 & n14555 ) | ( n14554 & n14555 ) ;
  assign n14557 = n5911 & ~n14014 ;
  assign n14558 = n14546 | n14557 ;
  assign n14559 = n14556 & n14558 ;
  assign n14560 = ( ~n14546 & n14556 ) | ( ~n14546 & n14557 ) | ( n14556 & n14557 ) ;
  assign n14561 = ( n14546 & ~n14559 ) | ( n14546 & n14560 ) | ( ~n14559 & n14560 ) ;
  assign n14562 = ( ~n14202 & n14545 ) | ( ~n14202 & n14561 ) | ( n14545 & n14561 ) ;
  assign n14563 = ( n14202 & n14545 ) | ( n14202 & n14561 ) | ( n14545 & n14561 ) ;
  assign n14564 = ( n14202 & n14562 ) | ( n14202 & ~n14563 ) | ( n14562 & ~n14563 ) ;
  assign n14565 = ( n14368 & n14535 ) | ( n14368 & n14564 ) | ( n14535 & n14564 ) ;
  assign n14566 = n36 & n13477 ;
  assign n14567 = x5 & n14566 ;
  assign n14568 = n8721 & n13475 ;
  assign n14569 = n8340 & ~n13473 ;
  assign n14570 = n40 | n14569 ;
  assign n14571 = n14568 | n14570 ;
  assign n14572 = x5 & ~n14571 ;
  assign n14573 = ( ~x5 & n14566 ) | ( ~x5 & n14571 ) | ( n14566 & n14571 ) ;
  assign n14574 = ( ~n14567 & n14572 ) | ( ~n14567 & n14573 ) | ( n14572 & n14573 ) ;
  assign n14575 = n7644 & ~n10235 ;
  assign n14576 = x8 & n14575 ;
  assign n14577 = n7341 & n10214 ;
  assign n14578 = n7345 | n14577 ;
  assign n14579 = ( ~n13280 & n14577 ) | ( ~n13280 & n14578 ) | ( n14577 & n14578 ) ;
  assign n14580 = n7346 | n14579 ;
  assign n14581 = ( ~n13285 & n14579 ) | ( ~n13285 & n14580 ) | ( n14579 & n14580 ) ;
  assign n14582 = x8 & ~n14581 ;
  assign n14583 = ( ~x8 & n14575 ) | ( ~x8 & n14581 ) | ( n14575 & n14581 ) ;
  assign n14584 = ( ~n14576 & n14582 ) | ( ~n14576 & n14583 ) | ( n14582 & n14583 ) ;
  assign n14585 = n6571 & n12756 ;
  assign n14586 = x11 & n14585 ;
  assign n14587 = n6567 & n10329 ;
  assign n14588 = n6570 | n14587 ;
  assign n14589 = ( ~n10237 & n14587 ) | ( ~n10237 & n14588 ) | ( n14587 & n14588 ) ;
  assign n14590 = n6796 & ~n10332 ;
  assign n14591 = n14589 | n14590 ;
  assign n14592 = x11 & ~n14591 ;
  assign n14593 = ( ~x11 & n14585 ) | ( ~x11 & n14591 ) | ( n14585 & n14591 ) ;
  assign n14594 = ( ~n14586 & n14592 ) | ( ~n14586 & n14593 ) | ( n14592 & n14593 ) ;
  assign n14595 = n6332 & n10239 ;
  assign n14596 = x14 & n14595 ;
  assign n14597 = n5909 & n10241 ;
  assign n14598 = n5914 | n14597 ;
  assign n14599 = ( n10326 & n14597 ) | ( n10326 & n14598 ) | ( n14597 & n14598 ) ;
  assign n14600 = n5915 | n14599 ;
  assign n14601 = ( n12222 & n14599 ) | ( n12222 & n14600 ) | ( n14599 & n14600 ) ;
  assign n14602 = x14 & ~n14601 ;
  assign n14603 = ( ~x14 & n14595 ) | ( ~x14 & n14601 ) | ( n14595 & n14601 ) ;
  assign n14604 = ( ~n14596 & n14602 ) | ( ~n14596 & n14603 ) | ( n14602 & n14603 ) ;
  assign n14605 = n5418 & ~n11989 ;
  assign n14606 = x17 & n14605 ;
  assign n14607 = n5417 & n10243 ;
  assign n14608 = n5584 & ~n10320 ;
  assign n14609 = n5413 & n10245 ;
  assign n14610 = n14608 | n14609 ;
  assign n14611 = n14607 | n14610 ;
  assign n14612 = x17 & ~n14611 ;
  assign n14613 = ( ~x17 & n14605 ) | ( ~x17 & n14611 ) | ( n14605 & n14611 ) ;
  assign n14614 = ( ~n14606 & n14612 ) | ( ~n14606 & n14613 ) | ( n14612 & n14613 ) ;
  assign n14615 = n4879 & ~n11691 ;
  assign n14616 = x20 & n14615 ;
  assign n14617 = n4874 & n10312 ;
  assign n14618 = n4878 | n14617 ;
  assign n14619 = ( ~n10316 & n14617 ) | ( ~n10316 & n14618 ) | ( n14617 & n14618 ) ;
  assign n14620 = n5232 & n10247 ;
  assign n14621 = n14619 | n14620 ;
  assign n14622 = x20 & ~n14621 ;
  assign n14623 = ( ~x20 & n14615 ) | ( ~x20 & n14621 ) | ( n14615 & n14621 ) ;
  assign n14624 = ( ~n14616 & n14622 ) | ( ~n14616 & n14623 ) | ( n14622 & n14623 ) ;
  assign n14625 = n4637 & n10251 ;
  assign n14626 = x23 & n14625 ;
  assign n14627 = n4584 & ~n10253 ;
  assign n14628 = n4649 | n14627 ;
  assign n14629 = ( ~n10249 & n14627 ) | ( ~n10249 & n14628 ) | ( n14627 & n14628 ) ;
  assign n14630 = n4591 | n14629 ;
  assign n14631 = ( ~n10441 & n14629 ) | ( ~n10441 & n14630 ) | ( n14629 & n14630 ) ;
  assign n14632 = x23 & ~n14631 ;
  assign n14633 = ( ~x23 & n14625 ) | ( ~x23 & n14631 ) | ( n14625 & n14631 ) ;
  assign n14634 = ( ~n14626 & n14632 ) | ( ~n14626 & n14633 ) | ( n14632 & n14633 ) ;
  assign n14635 = n4215 & n10255 ;
  assign n14636 = n4200 & n10257 ;
  assign n14637 = n2083 & n10259 ;
  assign n14638 = n14636 | n14637 ;
  assign n14639 = n14635 | n14638 ;
  assign n14640 = x26 & n14639 ;
  assign n14641 = n4203 & n11148 ;
  assign n14642 = ( ~x26 & n14639 ) | ( ~x26 & n14641 ) | ( n14639 & n14641 ) ;
  assign n14643 = x26 & ~n14641 ;
  assign n14644 = ( ~n14640 & n14642 ) | ( ~n14640 & n14643 ) | ( n14642 & n14643 ) ;
  assign n14645 = n3541 & n11049 ;
  assign n14646 = x29 & n14645 ;
  assign n14647 = n3536 & n10265 ;
  assign n14648 = n4039 | n14647 ;
  assign n14649 = ( n10261 & n14647 ) | ( n10261 & n14648 ) | ( n14647 & n14648 ) ;
  assign n14650 = n3501 & n10263 ;
  assign n14651 = n14649 | n14650 ;
  assign n14652 = x29 & ~n14651 ;
  assign n14653 = ( ~x29 & n14645 ) | ( ~x29 & n14651 ) | ( n14645 & n14651 ) ;
  assign n14654 = ( ~n14646 & n14652 ) | ( ~n14646 & n14653 ) | ( n14652 & n14653 ) ;
  assign n14655 = n1100 | n2332 ;
  assign n14656 = n74 | n674 ;
  assign n14657 = n14655 | n14656 ;
  assign n14658 = n356 | n2481 ;
  assign n14659 = n14657 | n14658 ;
  assign n14660 = n442 | n471 ;
  assign n14661 = n379 | n14660 ;
  assign n14662 = n3032 | n14661 ;
  assign n14663 = n1471 | n14662 ;
  assign n14664 = n14659 | n14663 ;
  assign n14665 = n141 | n616 ;
  assign n14666 = n1720 | n14665 ;
  assign n14667 = n914 | n14666 ;
  assign n14668 = n2419 | n14667 ;
  assign n14669 = n14664 | n14668 ;
  assign n14670 = n623 | n704 ;
  assign n14671 = n1254 | n14670 ;
  assign n14672 = n357 | n362 ;
  assign n14673 = n185 | n14672 ;
  assign n14674 = n14671 | n14673 ;
  assign n14675 = n83 | n212 ;
  assign n14676 = n14674 | n14675 ;
  assign n14677 = n3160 & ~n4949 ;
  assign n14678 = ~n12846 & n14677 ;
  assign n14679 = ~n14676 & n14678 ;
  assign n14680 = n2245 | n12868 ;
  assign n14681 = n14679 & ~n14680 ;
  assign n14682 = ~n14669 & n14681 ;
  assign n14683 = ~n13927 & n14682 ;
  assign n14684 = n3273 & n10271 ;
  assign n14685 = n3270 | n14684 ;
  assign n14686 = ( n10267 & n14684 ) | ( n10267 & n14685 ) | ( n14684 & n14685 ) ;
  assign n14687 = n390 | n14686 ;
  assign n14688 = ( ~n10787 & n14686 ) | ( ~n10787 & n14687 ) | ( n14686 & n14687 ) ;
  assign n14689 = n3274 & ~n10269 ;
  assign n14690 = n14688 | n14689 ;
  assign n14691 = ( n13983 & n14683 ) | ( n13983 & ~n14690 ) | ( n14683 & ~n14690 ) ;
  assign n14692 = ( ~n13983 & n14683 ) | ( ~n13983 & n14690 ) | ( n14683 & n14690 ) ;
  assign n14693 = ( ~n14683 & n14691 ) | ( ~n14683 & n14692 ) | ( n14691 & n14692 ) ;
  assign n14694 = ( n14468 & n14654 ) | ( n14468 & ~n14693 ) | ( n14654 & ~n14693 ) ;
  assign n14695 = ( ~n14468 & n14654 ) | ( ~n14468 & n14693 ) | ( n14654 & n14693 ) ;
  assign n14696 = ( ~n14654 & n14694 ) | ( ~n14654 & n14695 ) | ( n14694 & n14695 ) ;
  assign n14697 = ( ~n14471 & n14644 ) | ( ~n14471 & n14696 ) | ( n14644 & n14696 ) ;
  assign n14698 = ( n14471 & n14644 ) | ( n14471 & ~n14696 ) | ( n14644 & ~n14696 ) ;
  assign n14699 = ( ~n14644 & n14697 ) | ( ~n14644 & n14698 ) | ( n14697 & n14698 ) ;
  assign n14700 = ( ~n14484 & n14634 ) | ( ~n14484 & n14699 ) | ( n14634 & n14699 ) ;
  assign n14701 = ( n14484 & n14634 ) | ( n14484 & ~n14699 ) | ( n14634 & ~n14699 ) ;
  assign n14702 = ( ~n14634 & n14700 ) | ( ~n14634 & n14701 ) | ( n14700 & n14701 ) ;
  assign n14703 = ( ~n14488 & n14624 ) | ( ~n14488 & n14702 ) | ( n14624 & n14702 ) ;
  assign n14704 = ( n14488 & n14624 ) | ( n14488 & ~n14702 ) | ( n14624 & ~n14702 ) ;
  assign n14705 = ( ~n14624 & n14703 ) | ( ~n14624 & n14704 ) | ( n14703 & n14704 ) ;
  assign n14706 = ( ~n14490 & n14614 ) | ( ~n14490 & n14705 ) | ( n14614 & n14705 ) ;
  assign n14707 = ( n14490 & n14614 ) | ( n14490 & ~n14705 ) | ( n14614 & ~n14705 ) ;
  assign n14708 = ( ~n14614 & n14706 ) | ( ~n14614 & n14707 ) | ( n14706 & n14707 ) ;
  assign n14709 = ( n14494 & n14604 ) | ( n14494 & ~n14708 ) | ( n14604 & ~n14708 ) ;
  assign n14710 = ( ~n14494 & n14604 ) | ( ~n14494 & n14708 ) | ( n14604 & n14708 ) ;
  assign n14711 = ( ~n14604 & n14709 ) | ( ~n14604 & n14710 ) | ( n14709 & n14710 ) ;
  assign n14712 = ( ~n14497 & n14594 ) | ( ~n14497 & n14711 ) | ( n14594 & n14711 ) ;
  assign n14713 = ( n14497 & n14594 ) | ( n14497 & ~n14711 ) | ( n14594 & ~n14711 ) ;
  assign n14714 = ( ~n14594 & n14712 ) | ( ~n14594 & n14713 ) | ( n14712 & n14713 ) ;
  assign n14715 = ( ~n14510 & n14584 ) | ( ~n14510 & n14714 ) | ( n14584 & n14714 ) ;
  assign n14716 = ( n14510 & n14584 ) | ( n14510 & ~n14714 ) | ( n14584 & ~n14714 ) ;
  assign n14717 = ( ~n14584 & n14715 ) | ( ~n14584 & n14716 ) | ( n14715 & n14716 ) ;
  assign n14718 = ( n14513 & ~n14574 ) | ( n14513 & n14717 ) | ( ~n14574 & n14717 ) ;
  assign n14719 = ( n14513 & n14574 ) | ( n14513 & ~n14717 ) | ( n14574 & ~n14717 ) ;
  assign n14720 = ( ~n14513 & n14718 ) | ( ~n14513 & n14719 ) | ( n14718 & n14719 ) ;
  assign n14721 = ( ~n14516 & n14519 ) | ( ~n14516 & n14720 ) | ( n14519 & n14720 ) ;
  assign n14722 = ( n14516 & n14519 ) | ( n14516 & ~n14720 ) | ( n14519 & ~n14720 ) ;
  assign n14723 = ( ~n14519 & n14721 ) | ( ~n14519 & n14722 ) | ( n14721 & n14722 ) ;
  assign n14724 = n40 & ~n14723 ;
  assign n14725 = n8721 & n14520 ;
  assign n14726 = n8340 & n14352 ;
  assign n14727 = n14725 | n14726 ;
  assign n14728 = n14724 | n14727 ;
  assign n14729 = x5 & n14728 ;
  assign n14730 = n14520 | n14527 ;
  assign n14731 = n14723 & ~n14730 ;
  assign n14732 = ~n14529 & n14723 ;
  assign n14733 = ( ~n14529 & n14723 ) | ( ~n14529 & n14730 ) | ( n14723 & n14730 ) ;
  assign n14734 = ( n14731 & ~n14732 ) | ( n14731 & n14733 ) | ( ~n14732 & n14733 ) ;
  assign n14735 = n8341 & ~n14734 ;
  assign n14736 = ( ~x5 & n14728 ) | ( ~x5 & n14735 ) | ( n14728 & n14735 ) ;
  assign n14737 = x5 & ~n14735 ;
  assign n14738 = ( ~n14729 & n14736 ) | ( ~n14729 & n14737 ) | ( n14736 & n14737 ) ;
  assign n14739 = n7345 & n13992 ;
  assign n14740 = n7644 & n13996 ;
  assign n14741 = n7341 & n13998 ;
  assign n14742 = n14740 | n14741 ;
  assign n14743 = n14739 | n14742 ;
  assign n14744 = x8 & n14743 ;
  assign n14745 = n7346 & n14024 ;
  assign n14746 = x8 & ~n14745 ;
  assign n14747 = ( ~x8 & n14743 ) | ( ~x8 & n14745 ) | ( n14743 & n14745 ) ;
  assign n14748 = ( ~n14744 & n14746 ) | ( ~n14744 & n14747 ) | ( n14746 & n14747 ) ;
  assign n14749 = n6796 & ~n14007 ;
  assign n14750 = x11 & n14749 ;
  assign n14751 = n6567 & n14002 ;
  assign n14752 = n6570 | n14751 ;
  assign n14753 = ( ~n14000 & n14751 ) | ( ~n14000 & n14752 ) | ( n14751 & n14752 ) ;
  assign n14754 = n6571 | n14753 ;
  assign n14755 = ( ~n14042 & n14753 ) | ( ~n14042 & n14754 ) | ( n14753 & n14754 ) ;
  assign n14756 = x11 & ~n14755 ;
  assign n14757 = ( ~x11 & n14749 ) | ( ~x11 & n14755 ) | ( n14749 & n14755 ) ;
  assign n14758 = ( ~n14750 & n14756 ) | ( ~n14750 & n14757 ) | ( n14756 & n14757 ) ;
  assign n14759 = n5915 & n14004 ;
  assign n14760 = n6332 & ~n14014 ;
  assign n14761 = ( ~n14014 & n14759 ) | ( ~n14014 & n14760 ) | ( n14759 & n14760 ) ;
  assign n14762 = ( n5911 & n5914 ) | ( n5911 & n14014 ) | ( n5914 & n14014 ) ;
  assign n14763 = ~n14004 & n14762 ;
  assign n14764 = n14761 | n14763 ;
  assign n14765 = x14 & n14557 ;
  assign n14766 = ~n14764 & n14765 ;
  assign n14767 = n14764 & ~n14765 ;
  assign n14768 = n14766 | n14767 ;
  assign n14769 = ( n14559 & n14758 ) | ( n14559 & n14768 ) | ( n14758 & n14768 ) ;
  assign n14770 = ( n14559 & ~n14758 ) | ( n14559 & n14768 ) | ( ~n14758 & n14768 ) ;
  assign n14771 = ( n14758 & ~n14769 ) | ( n14758 & n14770 ) | ( ~n14769 & n14770 ) ;
  assign n14772 = ( ~n14563 & n14748 ) | ( ~n14563 & n14771 ) | ( n14748 & n14771 ) ;
  assign n14773 = ( n14563 & n14748 ) | ( n14563 & n14771 ) | ( n14748 & n14771 ) ;
  assign n14774 = ( n14563 & n14772 ) | ( n14563 & ~n14773 ) | ( n14772 & ~n14773 ) ;
  assign n14775 = ( n14565 & n14738 ) | ( n14565 & n14774 ) | ( n14738 & n14774 ) ;
  assign n14776 = n7644 & ~n13280 ;
  assign n14777 = x8 & n14776 ;
  assign n14778 = n7345 & ~n13473 ;
  assign n14779 = n7341 & ~n10235 ;
  assign n14780 = n14778 | n14779 ;
  assign n14781 = n7346 | n14780 ;
  assign n14782 = ( ~n13480 & n14780 ) | ( ~n13480 & n14781 ) | ( n14780 & n14781 ) ;
  assign n14783 = x8 & ~n14782 ;
  assign n14784 = ( ~x8 & n14776 ) | ( ~x8 & n14782 ) | ( n14776 & n14782 ) ;
  assign n14785 = ( ~n14777 & n14783 ) | ( ~n14777 & n14784 ) | ( n14783 & n14784 ) ;
  assign n14786 = n6796 & ~n10237 ;
  assign n14787 = x11 & n14786 ;
  assign n14788 = n6567 & ~n10332 ;
  assign n14789 = n6570 | n14788 ;
  assign n14790 = ( n10214 & n14788 ) | ( n10214 & n14789 ) | ( n14788 & n14789 ) ;
  assign n14791 = n6571 | n14790 ;
  assign n14792 = ( n12953 & n14790 ) | ( n12953 & n14791 ) | ( n14790 & n14791 ) ;
  assign n14793 = x11 & ~n14792 ;
  assign n14794 = ( ~x11 & n14786 ) | ( ~x11 & n14792 ) | ( n14786 & n14792 ) ;
  assign n14795 = ( ~n14787 & n14793 ) | ( ~n14787 & n14794 ) | ( n14793 & n14794 ) ;
  assign n14796 = n6332 & n10326 ;
  assign n14797 = x14 & n14796 ;
  assign n14798 = n5909 & n10239 ;
  assign n14799 = n5914 | n14798 ;
  assign n14800 = ( n10329 & n14798 ) | ( n10329 & n14799 ) | ( n14798 & n14799 ) ;
  assign n14801 = n5915 | n14800 ;
  assign n14802 = ( n10397 & n14800 ) | ( n10397 & n14801 ) | ( n14800 & n14801 ) ;
  assign n14803 = x14 & ~n14802 ;
  assign n14804 = ( ~x14 & n14796 ) | ( ~x14 & n14802 ) | ( n14796 & n14802 ) ;
  assign n14805 = ( ~n14797 & n14803 ) | ( ~n14797 & n14804 ) | ( n14803 & n14804 ) ;
  assign n14806 = n5584 & n10243 ;
  assign n14807 = x17 & n14806 ;
  assign n14808 = n5413 & ~n10320 ;
  assign n14809 = n5417 | n14808 ;
  assign n14810 = ( n10241 & n14808 ) | ( n10241 & n14809 ) | ( n14808 & n14809 ) ;
  assign n14811 = n5418 | n14810 ;
  assign n14812 = ( n12105 & n14810 ) | ( n12105 & n14811 ) | ( n14810 & n14811 ) ;
  assign n14813 = x17 & ~n14812 ;
  assign n14814 = ( ~x17 & n14806 ) | ( ~x17 & n14812 ) | ( n14806 & n14812 ) ;
  assign n14815 = ( ~n14807 & n14813 ) | ( ~n14807 & n14814 ) | ( n14813 & n14814 ) ;
  assign n14816 = n4879 & ~n11676 ;
  assign n14817 = x20 & n14816 ;
  assign n14818 = n4874 & n10247 ;
  assign n14819 = n4878 | n14818 ;
  assign n14820 = ( n10245 & n14818 ) | ( n10245 & n14819 ) | ( n14818 & n14819 ) ;
  assign n14821 = n5232 & ~n10316 ;
  assign n14822 = n14820 | n14821 ;
  assign n14823 = x20 & ~n14822 ;
  assign n14824 = ( ~x20 & n14816 ) | ( ~x20 & n14822 ) | ( n14816 & n14822 ) ;
  assign n14825 = ( ~n14817 & n14823 ) | ( ~n14817 & n14824 ) | ( n14823 & n14824 ) ;
  assign n14826 = n4649 & n10312 ;
  assign n14827 = x23 & n14826 ;
  assign n14828 = n4637 & ~n10249 ;
  assign n14829 = n4584 & n10251 ;
  assign n14830 = n14828 | n14829 ;
  assign n14831 = n4591 | n14830 ;
  assign n14832 = ( ~n11486 & n14830 ) | ( ~n11486 & n14831 ) | ( n14830 & n14831 ) ;
  assign n14833 = x23 & ~n14832 ;
  assign n14834 = ( ~x23 & n14826 ) | ( ~x23 & n14832 ) | ( n14826 & n14832 ) ;
  assign n14835 = ( ~n14827 & n14833 ) | ( ~n14827 & n14834 ) | ( n14833 & n14834 ) ;
  assign n14836 = n4203 & ~n11297 ;
  assign n14837 = n4215 & ~n10253 ;
  assign n14838 = n4200 & n10255 ;
  assign n14839 = n2083 & n10257 ;
  assign n14840 = n14838 | n14839 ;
  assign n14841 = n14837 | n14840 ;
  assign n14842 = n14836 | n14841 ;
  assign n14843 = n2693 | n3931 ;
  assign n14844 = n209 | n1439 ;
  assign n14845 = n14843 | n14844 ;
  assign n14846 = n3096 | n14845 ;
  assign n14847 = n12847 | n14303 ;
  assign n14848 = n14846 | n14847 ;
  assign n14849 = n296 | n688 ;
  assign n14850 = n863 | n14849 ;
  assign n14851 = n13404 | n14850 ;
  assign n14852 = n3294 | n14851 ;
  assign n14853 = n4491 | n14852 ;
  assign n14854 = n14848 | n14853 ;
  assign n14855 = n151 | n338 ;
  assign n14856 = n178 | n777 ;
  assign n14857 = n14855 | n14856 ;
  assign n14858 = n906 | n14857 ;
  assign n14859 = n524 | n1014 ;
  assign n14860 = n202 | n14859 ;
  assign n14861 = n14858 | n14860 ;
  assign n14862 = n839 | n14861 ;
  assign n14863 = n1786 | n2264 ;
  assign n14864 = n3344 | n14863 ;
  assign n14865 = n14862 | n14864 ;
  assign n14866 = n14854 | n14865 ;
  assign n14867 = n1184 | n2432 ;
  assign n14868 = n2420 | n14867 ;
  assign n14869 = n1507 | n14868 ;
  assign n14870 = n368 | n782 ;
  assign n14871 = n268 | n363 ;
  assign n14872 = n14870 | n14871 ;
  assign n14873 = n1231 | n14872 ;
  assign n14874 = n14869 | n14873 ;
  assign n14875 = n163 | n392 ;
  assign n14876 = n700 | n14875 ;
  assign n14877 = n3571 | n14876 ;
  assign n14878 = n629 | n756 ;
  assign n14879 = n14877 | n14878 ;
  assign n14880 = n2222 | n2475 ;
  assign n14881 = n4253 | n14880 ;
  assign n14882 = n70 | n659 ;
  assign n14883 = n1005 | n14882 ;
  assign n14884 = n14881 | n14883 ;
  assign n14885 = n14879 | n14884 ;
  assign n14886 = n14874 | n14885 ;
  assign n14887 = n14866 | n14886 ;
  assign n14888 = ( n14683 & ~n14692 ) | ( n14683 & n14887 ) | ( ~n14692 & n14887 ) ;
  assign n14889 = ( n14683 & n14692 ) | ( n14683 & ~n14887 ) | ( n14692 & ~n14887 ) ;
  assign n14890 = ( ~n14683 & n14888 ) | ( ~n14683 & n14889 ) | ( n14888 & n14889 ) ;
  assign n14891 = n3273 & ~n10269 ;
  assign n14892 = n3270 | n14891 ;
  assign n14893 = ( n10265 & n14891 ) | ( n10265 & n14892 ) | ( n14891 & n14892 ) ;
  assign n14894 = n390 | n14893 ;
  assign n14895 = ( n10804 & n14893 ) | ( n10804 & n14894 ) | ( n14893 & n14894 ) ;
  assign n14896 = n3274 & n10267 ;
  assign n14897 = n14895 | n14896 ;
  assign n14898 = ( ~n14694 & n14890 ) | ( ~n14694 & n14897 ) | ( n14890 & n14897 ) ;
  assign n14899 = ( n14694 & n14890 ) | ( n14694 & n14897 ) | ( n14890 & n14897 ) ;
  assign n14900 = ( n14694 & n14898 ) | ( n14694 & ~n14899 ) | ( n14898 & ~n14899 ) ;
  assign n14901 = n3541 & n10859 ;
  assign n14902 = n4039 & n10259 ;
  assign n14903 = n3501 & n10261 ;
  assign n14904 = n3536 & n10263 ;
  assign n14905 = n14903 | n14904 ;
  assign n14906 = n14902 | n14905 ;
  assign n14907 = n14901 | n14906 ;
  assign n14908 = n6269 & ~n14907 ;
  assign n14909 = ~n6269 & n14907 ;
  assign n14910 = n14908 | n14909 ;
  assign n14911 = ( n14842 & ~n14900 ) | ( n14842 & n14910 ) | ( ~n14900 & n14910 ) ;
  assign n14912 = ( n14842 & n14900 ) | ( n14842 & ~n14910 ) | ( n14900 & ~n14910 ) ;
  assign n14913 = ( ~n14842 & n14911 ) | ( ~n14842 & n14912 ) | ( n14911 & n14912 ) ;
  assign n14914 = ( n14698 & ~n14835 ) | ( n14698 & n14913 ) | ( ~n14835 & n14913 ) ;
  assign n14915 = ( n14698 & n14835 ) | ( n14698 & n14913 ) | ( n14835 & n14913 ) ;
  assign n14916 = ( n14835 & n14914 ) | ( n14835 & ~n14915 ) | ( n14914 & ~n14915 ) ;
  assign n14917 = ( n14701 & ~n14825 ) | ( n14701 & n14916 ) | ( ~n14825 & n14916 ) ;
  assign n14918 = ( n14701 & n14825 ) | ( n14701 & n14916 ) | ( n14825 & n14916 ) ;
  assign n14919 = ( n14825 & n14917 ) | ( n14825 & ~n14918 ) | ( n14917 & ~n14918 ) ;
  assign n14920 = ( n14704 & ~n14815 ) | ( n14704 & n14919 ) | ( ~n14815 & n14919 ) ;
  assign n14921 = ( n14704 & n14815 ) | ( n14704 & n14919 ) | ( n14815 & n14919 ) ;
  assign n14922 = ( n14815 & n14920 ) | ( n14815 & ~n14921 ) | ( n14920 & ~n14921 ) ;
  assign n14923 = ( n14707 & ~n14805 ) | ( n14707 & n14922 ) | ( ~n14805 & n14922 ) ;
  assign n14924 = ( n14707 & n14805 ) | ( n14707 & n14922 ) | ( n14805 & n14922 ) ;
  assign n14925 = ( n14805 & n14923 ) | ( n14805 & ~n14924 ) | ( n14923 & ~n14924 ) ;
  assign n14926 = ( n14709 & ~n14795 ) | ( n14709 & n14925 ) | ( ~n14795 & n14925 ) ;
  assign n14927 = ( n14709 & n14795 ) | ( n14709 & n14925 ) | ( n14795 & n14925 ) ;
  assign n14928 = ( n14795 & n14926 ) | ( n14795 & ~n14927 ) | ( n14926 & ~n14927 ) ;
  assign n14929 = ( n14713 & ~n14785 ) | ( n14713 & n14928 ) | ( ~n14785 & n14928 ) ;
  assign n14930 = ( n14713 & n14785 ) | ( n14713 & n14928 ) | ( n14785 & n14928 ) ;
  assign n14931 = ( n14785 & n14929 ) | ( n14785 & ~n14930 ) | ( n14929 & ~n14930 ) ;
  assign n14932 = ( x2 & ~x3 ) | ( x2 & x4 ) | ( ~x3 & x4 ) ;
  assign n14933 = ( x3 & ~x5 ) | ( x3 & n14932 ) | ( ~x5 & n14932 ) ;
  assign n14934 = n13475 & ~n14933 ;
  assign n14935 = ( n8339 & n13475 ) | ( n8339 & n14933 ) | ( n13475 & n14933 ) ;
  assign n14936 = ( n9196 & ~n14934 ) | ( n9196 & n14935 ) | ( ~n14934 & n14935 ) ;
  assign n14937 = ( n14716 & n14931 ) | ( n14716 & n14936 ) | ( n14931 & n14936 ) ;
  assign n14938 = ( n14716 & ~n14931 ) | ( n14716 & n14936 ) | ( ~n14931 & n14936 ) ;
  assign n14939 = ( n14931 & ~n14937 ) | ( n14931 & n14938 ) | ( ~n14937 & n14938 ) ;
  assign n14940 = ( ~n14719 & n14722 ) | ( ~n14719 & n14939 ) | ( n14722 & n14939 ) ;
  assign n14941 = ( n14719 & n14722 ) | ( n14719 & n14939 ) | ( n14722 & n14939 ) ;
  assign n14942 = ( n14719 & n14940 ) | ( n14719 & ~n14941 ) | ( n14940 & ~n14941 ) ;
  assign n14943 = n40 & n14942 ;
  assign n14944 = n8721 & ~n14723 ;
  assign n14945 = n8340 & n14520 ;
  assign n14946 = n14944 | n14945 ;
  assign n14947 = n14943 | n14946 ;
  assign n14948 = x5 & n14947 ;
  assign n14949 = ~n14723 & n14730 ;
  assign n14950 = n14942 & n14949 ;
  assign n14951 = ~n14732 & n14942 ;
  assign n14952 = ( n14732 & ~n14942 ) | ( n14732 & n14949 ) | ( ~n14942 & n14949 ) ;
  assign n14953 = ( ~n14950 & n14951 ) | ( ~n14950 & n14952 ) | ( n14951 & n14952 ) ;
  assign n14954 = n8341 & ~n14953 ;
  assign n14955 = ( ~x5 & n14947 ) | ( ~x5 & n14954 ) | ( n14947 & n14954 ) ;
  assign n14956 = x5 & ~n14954 ;
  assign n14957 = ( ~n14948 & n14955 ) | ( ~n14948 & n14956 ) | ( n14955 & n14956 ) ;
  assign n14958 = n7644 & n13992 ;
  assign n14959 = x8 & n14958 ;
  assign n14960 = n7341 & n13996 ;
  assign n14961 = n7345 | n14960 ;
  assign n14962 = ( n14352 & n14960 ) | ( n14352 & n14961 ) | ( n14960 & n14961 ) ;
  assign n14963 = n7346 | n14962 ;
  assign n14964 = ( n14363 & n14962 ) | ( n14363 & n14963 ) | ( n14962 & n14963 ) ;
  assign n14965 = x8 & ~n14964 ;
  assign n14966 = ( ~x8 & n14958 ) | ( ~x8 & n14964 ) | ( n14958 & n14964 ) ;
  assign n14967 = ( ~n14959 & n14965 ) | ( ~n14959 & n14966 ) | ( n14965 & n14966 ) ;
  assign n14968 = n6796 & ~n14000 ;
  assign n14969 = x11 & n14968 ;
  assign n14970 = n6567 & ~n14007 ;
  assign n14971 = n6570 | n14970 ;
  assign n14972 = ( n13998 & n14970 ) | ( n13998 & n14971 ) | ( n14970 & n14971 ) ;
  assign n14973 = n6571 | n14972 ;
  assign n14974 = ( n14115 & n14972 ) | ( n14115 & n14973 ) | ( n14972 & n14973 ) ;
  assign n14975 = x11 & ~n14974 ;
  assign n14976 = ( ~x11 & n14968 ) | ( ~x11 & n14974 ) | ( n14968 & n14974 ) ;
  assign n14977 = ( ~n14969 & n14975 ) | ( ~n14969 & n14976 ) | ( n14975 & n14976 ) ;
  assign n14978 = x14 & ~n14557 ;
  assign n14979 = ~n14764 & n14978 ;
  assign n14980 = x14 & ~n14979 ;
  assign n14981 = n6332 & ~n14004 ;
  assign n14982 = n5909 & ~n14014 ;
  assign n14983 = n14981 | n14982 ;
  assign n14984 = n5915 | n14983 ;
  assign n14985 = ( n14072 & n14983 ) | ( n14072 & n14984 ) | ( n14983 & n14984 ) ;
  assign n14986 = n5914 & n14002 ;
  assign n14987 = n14985 | n14986 ;
  assign n14988 = n14980 & ~n14987 ;
  assign n14989 = ~n14980 & n14987 ;
  assign n14990 = n14988 | n14989 ;
  assign n14991 = ( n14769 & ~n14977 ) | ( n14769 & n14990 ) | ( ~n14977 & n14990 ) ;
  assign n14992 = ( n14769 & n14977 ) | ( n14769 & n14990 ) | ( n14977 & n14990 ) ;
  assign n14993 = ( n14977 & n14991 ) | ( n14977 & ~n14992 ) | ( n14991 & ~n14992 ) ;
  assign n14994 = ( n14773 & ~n14967 ) | ( n14773 & n14993 ) | ( ~n14967 & n14993 ) ;
  assign n14995 = ( n14773 & n14967 ) | ( n14773 & n14993 ) | ( n14967 & n14993 ) ;
  assign n14996 = ( n14967 & n14994 ) | ( n14967 & ~n14995 ) | ( n14994 & ~n14995 ) ;
  assign n14997 = ( n14775 & n14957 ) | ( n14775 & n14996 ) | ( n14957 & n14996 ) ;
  assign n14998 = n7345 & n14520 ;
  assign n14999 = n7346 | n14998 ;
  assign n15000 = ( n14531 & n14998 ) | ( n14531 & n14999 ) | ( n14998 & n14999 ) ;
  assign n15001 = n7341 & n13992 ;
  assign n15002 = ( ~x8 & n15000 ) | ( ~x8 & n15001 ) | ( n15000 & n15001 ) ;
  assign n15003 = n7644 & n14352 ;
  assign n15004 = x8 & ~n15001 ;
  assign n15005 = n15003 | n15004 ;
  assign n15006 = ( n15000 & n15003 ) | ( n15000 & n15004 ) | ( n15003 & n15004 ) ;
  assign n15007 = ( n15002 & n15005 ) | ( n15002 & ~n15006 ) | ( n15005 & ~n15006 ) ;
  assign n15008 = n6571 & ~n14130 ;
  assign n15009 = x11 & n15008 ;
  assign n15010 = n6567 & ~n14000 ;
  assign n15011 = n6570 | n15010 ;
  assign n15012 = ( n13996 & n15010 ) | ( n13996 & n15011 ) | ( n15010 & n15011 ) ;
  assign n15013 = n6796 & n13998 ;
  assign n15014 = n15012 | n15013 ;
  assign n15015 = x11 & ~n15014 ;
  assign n15016 = ( ~x11 & n15008 ) | ( ~x11 & n15014 ) | ( n15008 & n15014 ) ;
  assign n15017 = ( ~n15009 & n15015 ) | ( ~n15009 & n15016 ) | ( n15015 & n15016 ) ;
  assign n15018 = n14979 & ~n14987 ;
  assign n15019 = n6332 & n14002 ;
  assign n15020 = x14 & n15019 ;
  assign n15021 = n5909 & ~n14004 ;
  assign n15022 = n5914 | n15021 ;
  assign n15023 = ( ~n14007 & n15021 ) | ( ~n14007 & n15022 ) | ( n15021 & n15022 ) ;
  assign n15024 = n5915 | n15023 ;
  assign n15025 = ( n14066 & n15023 ) | ( n14066 & n15024 ) | ( n15023 & n15024 ) ;
  assign n15026 = x14 & ~n15025 ;
  assign n15027 = ( ~x14 & n15019 ) | ( ~x14 & n15025 ) | ( n15019 & n15025 ) ;
  assign n15028 = ( ~n15020 & n15026 ) | ( ~n15020 & n15027 ) | ( n15026 & n15027 ) ;
  assign n15029 = n5414 & ~n14014 ;
  assign n15030 = n15018 | n15029 ;
  assign n15031 = n15028 & n15030 ;
  assign n15032 = ( ~n15018 & n15028 ) | ( ~n15018 & n15029 ) | ( n15028 & n15029 ) ;
  assign n15033 = ( n15018 & ~n15031 ) | ( n15018 & n15032 ) | ( ~n15031 & n15032 ) ;
  assign n15034 = ( ~n14992 & n15017 ) | ( ~n14992 & n15033 ) | ( n15017 & n15033 ) ;
  assign n15035 = ( n14992 & n15017 ) | ( n14992 & n15033 ) | ( n15017 & n15033 ) ;
  assign n15036 = ( n14992 & n15034 ) | ( n14992 & ~n15035 ) | ( n15034 & ~n15035 ) ;
  assign n15037 = ( n14995 & ~n15007 ) | ( n14995 & n15036 ) | ( ~n15007 & n15036 ) ;
  assign n15038 = ( n14995 & n15007 ) | ( n14995 & n15036 ) | ( n15007 & n15036 ) ;
  assign n15039 = ( n15007 & n15037 ) | ( n15007 & ~n15038 ) | ( n15037 & ~n15038 ) ;
  assign n15040 = n7341 & ~n13280 ;
  assign n15041 = n7345 | n15040 ;
  assign n15042 = ( n13475 & n15040 ) | ( n13475 & n15041 ) | ( n15040 & n15041 ) ;
  assign n15043 = n7644 & ~n13473 ;
  assign n15044 = n15042 | n15043 ;
  assign n15045 = x8 & n15044 ;
  assign n15046 = n7346 & n13671 ;
  assign n15047 = ( ~x8 & n15044 ) | ( ~x8 & n15046 ) | ( n15044 & n15046 ) ;
  assign n15048 = x8 & ~n15046 ;
  assign n15049 = ( ~n15045 & n15047 ) | ( ~n15045 & n15048 ) | ( n15047 & n15048 ) ;
  assign n15050 = n6796 & n10214 ;
  assign n15051 = x11 & n15050 ;
  assign n15052 = n6567 & ~n10237 ;
  assign n15053 = n6570 | n15052 ;
  assign n15054 = ( ~n10235 & n15052 ) | ( ~n10235 & n15053 ) | ( n15052 & n15053 ) ;
  assign n15055 = n6571 | n15054 ;
  assign n15056 = ( n10371 & n15054 ) | ( n10371 & n15055 ) | ( n15054 & n15055 ) ;
  assign n15057 = x11 & ~n15056 ;
  assign n15058 = ( ~x11 & n15050 ) | ( ~x11 & n15056 ) | ( n15050 & n15056 ) ;
  assign n15059 = ( ~n15051 & n15057 ) | ( ~n15051 & n15058 ) | ( n15057 & n15058 ) ;
  assign n15060 = n5909 & n10326 ;
  assign n15061 = n5914 | n15060 ;
  assign n15062 = ( ~n10332 & n15060 ) | ( ~n10332 & n15061 ) | ( n15060 & n15061 ) ;
  assign n15063 = n6332 & n10329 ;
  assign n15064 = n15062 | n15063 ;
  assign n15065 = x14 & n15064 ;
  assign n15066 = n5915 & ~n10383 ;
  assign n15067 = x14 & ~n15066 ;
  assign n15068 = ( ~x14 & n15064 ) | ( ~x14 & n15066 ) | ( n15064 & n15066 ) ;
  assign n15069 = ( ~n15065 & n15067 ) | ( ~n15065 & n15068 ) | ( n15067 & n15068 ) ;
  assign n15070 = n5584 & n10241 ;
  assign n15071 = x17 & n15070 ;
  assign n15072 = n5413 & n10243 ;
  assign n15073 = n5417 | n15072 ;
  assign n15074 = ( n10239 & n15072 ) | ( n10239 & n15073 ) | ( n15072 & n15073 ) ;
  assign n15075 = n5418 | n15074 ;
  assign n15076 = ( n12575 & n15074 ) | ( n12575 & n15075 ) | ( n15074 & n15075 ) ;
  assign n15077 = x17 & ~n15076 ;
  assign n15078 = ( ~x17 & n15070 ) | ( ~x17 & n15076 ) | ( n15070 & n15076 ) ;
  assign n15079 = ( ~n15071 & n15077 ) | ( ~n15071 & n15078 ) | ( n15077 & n15078 ) ;
  assign n15080 = n4878 & ~n10320 ;
  assign n15081 = n5232 & n10245 ;
  assign n15082 = n4874 & ~n10316 ;
  assign n15083 = n15081 | n15082 ;
  assign n15084 = n15080 | n15083 ;
  assign n15085 = x20 & n15084 ;
  assign n15086 = n4879 & ~n10414 ;
  assign n15087 = x20 & ~n15086 ;
  assign n15088 = ( ~x20 & n15084 ) | ( ~x20 & n15086 ) | ( n15084 & n15086 ) ;
  assign n15089 = ( ~n15085 & n15087 ) | ( ~n15085 & n15088 ) | ( n15087 & n15088 ) ;
  assign n15090 = n4637 & n10312 ;
  assign n15091 = x23 & n15090 ;
  assign n15092 = n4584 & ~n10249 ;
  assign n15093 = n4649 | n15092 ;
  assign n15094 = ( n10247 & n15092 ) | ( n10247 & n15093 ) | ( n15092 & n15093 ) ;
  assign n15095 = n4591 | n15094 ;
  assign n15096 = ( n10428 & n15094 ) | ( n10428 & n15095 ) | ( n15094 & n15095 ) ;
  assign n15097 = x23 & ~n15096 ;
  assign n15098 = ( ~x23 & n15090 ) | ( ~x23 & n15096 ) | ( n15090 & n15096 ) ;
  assign n15099 = ( ~n15091 & n15097 ) | ( ~n15091 & n15098 ) | ( n15097 & n15098 ) ;
  assign n15100 = x26 & ~n14842 ;
  assign n15101 = ~x26 & n14842 ;
  assign n15102 = n15100 | n15101 ;
  assign n15103 = x29 & ~n14907 ;
  assign n15104 = ~x29 & n14907 ;
  assign n15105 = n15103 | n15104 ;
  assign n15106 = ( n14900 & n15102 ) | ( n14900 & n15105 ) | ( n15102 & n15105 ) ;
  assign n15107 = n4215 & n10251 ;
  assign n15108 = n4200 & ~n10253 ;
  assign n15109 = n2083 & n10255 ;
  assign n15110 = n15108 | n15109 ;
  assign n15111 = n15107 | n15110 ;
  assign n15112 = x26 & n15111 ;
  assign n15113 = n4203 & ~n11309 ;
  assign n15114 = ( ~x26 & n15111 ) | ( ~x26 & n15113 ) | ( n15111 & n15113 ) ;
  assign n15115 = x26 & ~n15113 ;
  assign n15116 = ( ~n15112 & n15114 ) | ( ~n15112 & n15115 ) | ( n15114 & n15115 ) ;
  assign n15117 = n13983 & ~n14887 ;
  assign n15118 = ( ~n14683 & n14690 ) | ( ~n14683 & n15117 ) | ( n14690 & n15117 ) ;
  assign n15119 = n1816 | n2758 ;
  assign n15120 = n2123 | n2381 ;
  assign n15121 = n15119 | n15120 ;
  assign n15122 = n1796 | n15121 ;
  assign n15123 = n185 | n253 ;
  assign n15124 = n3054 | n15123 ;
  assign n15125 = n279 | n715 ;
  assign n15126 = ~n567 & n618 ;
  assign n15127 = ~n15125 & n15126 ;
  assign n15128 = ~n15124 & n15127 ;
  assign n15129 = ~n3193 & n15128 ;
  assign n15130 = ~n15122 & n15129 ;
  assign n15131 = n169 | n461 ;
  assign n15132 = n15130 & ~n15131 ;
  assign n15133 = ~n3723 & n15132 ;
  assign n15134 = ( n13983 & ~n14887 ) | ( n13983 & n15118 ) | ( ~n14887 & n15118 ) ;
  assign n15135 = ( n15118 & n15133 ) | ( n15118 & ~n15134 ) | ( n15133 & ~n15134 ) ;
  assign n15136 = ( n15118 & ~n15133 ) | ( n15118 & n15134 ) | ( ~n15133 & n15134 ) ;
  assign n15137 = ( ~n15118 & n15135 ) | ( ~n15118 & n15136 ) | ( n15135 & n15136 ) ;
  assign n15138 = n3273 & n10267 ;
  assign n15139 = n3270 | n15138 ;
  assign n15140 = ( n10263 & n15138 ) | ( n10263 & n15139 ) | ( n15138 & n15139 ) ;
  assign n15141 = n390 | n15140 ;
  assign n15142 = ( n10874 & n15140 ) | ( n10874 & n15141 ) | ( n15140 & n15141 ) ;
  assign n15143 = n3274 & n10265 ;
  assign n15144 = n15142 | n15143 ;
  assign n15145 = ( n14899 & ~n15137 ) | ( n14899 & n15144 ) | ( ~n15137 & n15144 ) ;
  assign n15146 = ( n14899 & n15137 ) | ( n14899 & ~n15144 ) | ( n15137 & ~n15144 ) ;
  assign n15147 = ( ~n14899 & n15145 ) | ( ~n14899 & n15146 ) | ( n15145 & n15146 ) ;
  assign n15148 = n3541 & n11065 ;
  assign n15149 = x29 & n15148 ;
  assign n15150 = n3536 & n10261 ;
  assign n15151 = n4039 | n15150 ;
  assign n15152 = ( n10257 & n15150 ) | ( n10257 & n15151 ) | ( n15150 & n15151 ) ;
  assign n15153 = n3501 & n10259 ;
  assign n15154 = n15152 | n15153 ;
  assign n15155 = x29 & ~n15154 ;
  assign n15156 = ( ~x29 & n15148 ) | ( ~x29 & n15154 ) | ( n15148 & n15154 ) ;
  assign n15157 = ( ~n15149 & n15155 ) | ( ~n15149 & n15156 ) | ( n15155 & n15156 ) ;
  assign n15158 = ( n15116 & ~n15147 ) | ( n15116 & n15157 ) | ( ~n15147 & n15157 ) ;
  assign n15159 = ( n15116 & n15147 ) | ( n15116 & ~n15157 ) | ( n15147 & ~n15157 ) ;
  assign n15160 = ( ~n15116 & n15158 ) | ( ~n15116 & n15159 ) | ( n15158 & n15159 ) ;
  assign n15161 = ( n15099 & ~n15106 ) | ( n15099 & n15160 ) | ( ~n15106 & n15160 ) ;
  assign n15162 = ( n15099 & n15106 ) | ( n15099 & ~n15160 ) | ( n15106 & ~n15160 ) ;
  assign n15163 = ( ~n15099 & n15161 ) | ( ~n15099 & n15162 ) | ( n15161 & n15162 ) ;
  assign n15164 = ( n14915 & n15089 ) | ( n14915 & ~n15163 ) | ( n15089 & ~n15163 ) ;
  assign n15165 = ( ~n14915 & n15089 ) | ( ~n14915 & n15163 ) | ( n15089 & n15163 ) ;
  assign n15166 = ( ~n15089 & n15164 ) | ( ~n15089 & n15165 ) | ( n15164 & n15165 ) ;
  assign n15167 = ( ~n14918 & n15079 ) | ( ~n14918 & n15166 ) | ( n15079 & n15166 ) ;
  assign n15168 = ( n14918 & n15079 ) | ( n14918 & ~n15166 ) | ( n15079 & ~n15166 ) ;
  assign n15169 = ( ~n15079 & n15167 ) | ( ~n15079 & n15168 ) | ( n15167 & n15168 ) ;
  assign n15170 = ( ~n14921 & n15069 ) | ( ~n14921 & n15169 ) | ( n15069 & n15169 ) ;
  assign n15171 = ( n14921 & n15069 ) | ( n14921 & ~n15169 ) | ( n15069 & ~n15169 ) ;
  assign n15172 = ( ~n15069 & n15170 ) | ( ~n15069 & n15171 ) | ( n15170 & n15171 ) ;
  assign n15173 = ( n14924 & n15059 ) | ( n14924 & ~n15172 ) | ( n15059 & ~n15172 ) ;
  assign n15174 = ( ~n14924 & n15059 ) | ( ~n14924 & n15172 ) | ( n15059 & n15172 ) ;
  assign n15175 = ( ~n15059 & n15173 ) | ( ~n15059 & n15174 ) | ( n15173 & n15174 ) ;
  assign n15176 = ( n14927 & n15049 ) | ( n14927 & ~n15175 ) | ( n15049 & ~n15175 ) ;
  assign n15177 = ( ~n14927 & n15049 ) | ( ~n14927 & n15175 ) | ( n15049 & n15175 ) ;
  assign n15178 = ( ~n15049 & n15176 ) | ( ~n15049 & n15177 ) | ( n15176 & n15177 ) ;
  assign n15179 = ( n14930 & n14933 ) | ( n14930 & ~n15178 ) | ( n14933 & ~n15178 ) ;
  assign n15180 = ( n14930 & ~n14933 ) | ( n14930 & n15178 ) | ( ~n14933 & n15178 ) ;
  assign n15181 = ( ~n14930 & n15179 ) | ( ~n14930 & n15180 ) | ( n15179 & n15180 ) ;
  assign n15182 = ( ~n14937 & n14941 ) | ( ~n14937 & n15181 ) | ( n14941 & n15181 ) ;
  assign n15183 = ( n14937 & n14941 ) | ( n14937 & ~n15181 ) | ( n14941 & ~n15181 ) ;
  assign n15184 = ( ~n14941 & n15182 ) | ( ~n14941 & n15183 ) | ( n15182 & n15183 ) ;
  assign n15185 = n40 & ~n15184 ;
  assign n15186 = n8721 & n14942 ;
  assign n15187 = n8340 & ~n14723 ;
  assign n15188 = n15186 | n15187 ;
  assign n15189 = n15185 | n15188 ;
  assign n15190 = x5 & n15189 ;
  assign n15191 = n14942 | n14949 ;
  assign n15192 = n15184 & ~n15191 ;
  assign n15193 = ~n14951 & n15184 ;
  assign n15194 = ( ~n14951 & n15184 ) | ( ~n14951 & n15191 ) | ( n15184 & n15191 ) ;
  assign n15195 = ( n15192 & ~n15193 ) | ( n15192 & n15194 ) | ( ~n15193 & n15194 ) ;
  assign n15196 = n8341 & ~n15195 ;
  assign n15197 = ( ~x5 & n15189 ) | ( ~x5 & n15196 ) | ( n15189 & n15196 ) ;
  assign n15198 = x5 & ~n15196 ;
  assign n15199 = ( ~n15190 & n15197 ) | ( ~n15190 & n15198 ) | ( n15197 & n15198 ) ;
  assign n15200 = ( n14997 & n15039 ) | ( n14997 & n15199 ) | ( n15039 & n15199 ) ;
  assign n15201 = n7346 & ~n14734 ;
  assign n15202 = x8 & n15201 ;
  assign n15203 = n7341 & n14352 ;
  assign n15204 = n7345 | n15203 ;
  assign n15205 = ( ~n14723 & n15203 ) | ( ~n14723 & n15204 ) | ( n15203 & n15204 ) ;
  assign n15206 = n7644 & n14520 ;
  assign n15207 = n15205 | n15206 ;
  assign n15208 = x8 & ~n15207 ;
  assign n15209 = ( ~x8 & n15201 ) | ( ~x8 & n15207 ) | ( n15201 & n15207 ) ;
  assign n15210 = ( ~n15202 & n15208 ) | ( ~n15202 & n15209 ) | ( n15208 & n15209 ) ;
  assign n15211 = n6570 & n13992 ;
  assign n15212 = x11 & n15211 ;
  assign n15213 = n6796 & n13996 ;
  assign n15214 = n6567 & n13998 ;
  assign n15215 = n15213 | n15214 ;
  assign n15216 = n6571 | n15215 ;
  assign n15217 = ( n14024 & n15215 ) | ( n14024 & n15216 ) | ( n15215 & n15216 ) ;
  assign n15218 = x11 & ~n15217 ;
  assign n15219 = ( ~x11 & n15211 ) | ( ~x11 & n15217 ) | ( n15211 & n15217 ) ;
  assign n15220 = ( ~n15212 & n15218 ) | ( ~n15212 & n15219 ) | ( n15218 & n15219 ) ;
  assign n15221 = n6332 & ~n14007 ;
  assign n15222 = x14 & n15221 ;
  assign n15223 = n5909 & n14002 ;
  assign n15224 = n5914 | n15223 ;
  assign n15225 = ( ~n14000 & n15223 ) | ( ~n14000 & n15224 ) | ( n15223 & n15224 ) ;
  assign n15226 = n5915 | n15225 ;
  assign n15227 = ( ~n14042 & n15225 ) | ( ~n14042 & n15226 ) | ( n15225 & n15226 ) ;
  assign n15228 = x14 & ~n15227 ;
  assign n15229 = ( ~x14 & n15221 ) | ( ~x14 & n15227 ) | ( n15221 & n15227 ) ;
  assign n15230 = ( ~n15222 & n15228 ) | ( ~n15222 & n15229 ) | ( n15228 & n15229 ) ;
  assign n15231 = n5418 & n14004 ;
  assign n15232 = n5584 & ~n14014 ;
  assign n15233 = ( ~n14014 & n15231 ) | ( ~n14014 & n15232 ) | ( n15231 & n15232 ) ;
  assign n15234 = ( n5414 & n5417 ) | ( n5414 & n14014 ) | ( n5417 & n14014 ) ;
  assign n15235 = ~n14004 & n15234 ;
  assign n15236 = n15233 | n15235 ;
  assign n15237 = x17 & n15029 ;
  assign n15238 = ~n15236 & n15237 ;
  assign n15239 = n15236 & ~n15237 ;
  assign n15240 = n15238 | n15239 ;
  assign n15241 = ( n15031 & n15230 ) | ( n15031 & n15240 ) | ( n15230 & n15240 ) ;
  assign n15242 = ( n15031 & ~n15230 ) | ( n15031 & n15240 ) | ( ~n15230 & n15240 ) ;
  assign n15243 = ( n15230 & ~n15241 ) | ( n15230 & n15242 ) | ( ~n15241 & n15242 ) ;
  assign n15244 = ( ~n15035 & n15220 ) | ( ~n15035 & n15243 ) | ( n15220 & n15243 ) ;
  assign n15245 = ( n15035 & n15220 ) | ( n15035 & n15243 ) | ( n15220 & n15243 ) ;
  assign n15246 = ( n15035 & n15244 ) | ( n15035 & ~n15245 ) | ( n15244 & ~n15245 ) ;
  assign n15247 = ( n15038 & n15210 ) | ( n15038 & n15246 ) | ( n15210 & n15246 ) ;
  assign n15248 = ( ~n15038 & n15210 ) | ( ~n15038 & n15246 ) | ( n15210 & n15246 ) ;
  assign n15249 = ( n15038 & ~n15247 ) | ( n15038 & n15248 ) | ( ~n15247 & n15248 ) ;
  assign n15250 = n7341 | n7345 ;
  assign n15251 = ( n7345 & ~n13473 ) | ( n7345 & n15250 ) | ( ~n13473 & n15250 ) ;
  assign n15252 = n7644 | n15251 ;
  assign n15253 = ( n13475 & n15251 ) | ( n13475 & n15252 ) | ( n15251 & n15252 ) ;
  assign n15254 = x8 & n15253 ;
  assign n15255 = n7342 & n13477 ;
  assign n15256 = x8 & ~n15255 ;
  assign n15257 = ( ~x8 & n15253 ) | ( ~x8 & n15255 ) | ( n15253 & n15255 ) ;
  assign n15258 = ( ~n15254 & n15256 ) | ( ~n15254 & n15257 ) | ( n15256 & n15257 ) ;
  assign n15259 = n6571 & ~n13285 ;
  assign n15260 = x11 & n15259 ;
  assign n15261 = n6567 & n10214 ;
  assign n15262 = n6570 | n15261 ;
  assign n15263 = ( ~n13280 & n15261 ) | ( ~n13280 & n15262 ) | ( n15261 & n15262 ) ;
  assign n15264 = n6796 & ~n10235 ;
  assign n15265 = n15263 | n15264 ;
  assign n15266 = x11 & ~n15265 ;
  assign n15267 = ( ~x11 & n15259 ) | ( ~x11 & n15265 ) | ( n15259 & n15265 ) ;
  assign n15268 = ( ~n15260 & n15266 ) | ( ~n15260 & n15267 ) | ( n15266 & n15267 ) ;
  assign n15269 = n5915 & n12756 ;
  assign n15270 = x14 & n15269 ;
  assign n15271 = n5914 & ~n10237 ;
  assign n15272 = n6332 & ~n10332 ;
  assign n15273 = n5909 & n10329 ;
  assign n15274 = n15272 | n15273 ;
  assign n15275 = n15271 | n15274 ;
  assign n15276 = x14 & ~n15275 ;
  assign n15277 = ( ~x14 & n15269 ) | ( ~x14 & n15275 ) | ( n15269 & n15275 ) ;
  assign n15278 = ( ~n15270 & n15276 ) | ( ~n15270 & n15277 ) | ( n15276 & n15277 ) ;
  assign n15279 = n5413 & n10241 ;
  assign n15280 = n5417 | n15279 ;
  assign n15281 = ( n10326 & n15279 ) | ( n10326 & n15280 ) | ( n15279 & n15280 ) ;
  assign n15282 = n5584 & n10239 ;
  assign n15283 = n15281 | n15282 ;
  assign n15284 = x17 & n15283 ;
  assign n15285 = n5418 & n12222 ;
  assign n15286 = x17 & ~n15285 ;
  assign n15287 = ( ~x17 & n15283 ) | ( ~x17 & n15285 ) | ( n15283 & n15285 ) ;
  assign n15288 = ( ~n15284 & n15286 ) | ( ~n15284 & n15287 ) | ( n15286 & n15287 ) ;
  assign n15289 = n4879 & ~n11989 ;
  assign n15290 = x20 & n15289 ;
  assign n15291 = n4878 & n10243 ;
  assign n15292 = n5232 & ~n10320 ;
  assign n15293 = n4874 & n10245 ;
  assign n15294 = n15292 | n15293 ;
  assign n15295 = n15291 | n15294 ;
  assign n15296 = x20 & ~n15295 ;
  assign n15297 = ( ~x20 & n15289 ) | ( ~x20 & n15295 ) | ( n15289 & n15295 ) ;
  assign n15298 = ( ~n15290 & n15296 ) | ( ~n15290 & n15297 ) | ( n15296 & n15297 ) ;
  assign n15299 = n4591 & ~n11691 ;
  assign n15300 = x23 & n15299 ;
  assign n15301 = n4584 & n10312 ;
  assign n15302 = n4649 | n15301 ;
  assign n15303 = ( ~n10316 & n15301 ) | ( ~n10316 & n15302 ) | ( n15301 & n15302 ) ;
  assign n15304 = n4637 & n10247 ;
  assign n15305 = n15303 | n15304 ;
  assign n15306 = x23 & ~n15305 ;
  assign n15307 = ( ~x23 & n15299 ) | ( ~x23 & n15305 ) | ( n15299 & n15305 ) ;
  assign n15308 = ( ~n15300 & n15306 ) | ( ~n15300 & n15307 ) | ( n15306 & n15307 ) ;
  assign n15309 = n4215 & ~n10249 ;
  assign n15310 = n4200 & n10251 ;
  assign n15311 = n2083 & ~n10253 ;
  assign n15312 = n15310 | n15311 ;
  assign n15313 = n15309 | n15312 ;
  assign n15314 = x26 & n15313 ;
  assign n15315 = n4203 & ~n10441 ;
  assign n15316 = ( ~x26 & n15313 ) | ( ~x26 & n15315 ) | ( n15313 & n15315 ) ;
  assign n15317 = x26 & ~n15315 ;
  assign n15318 = ( ~n15314 & n15316 ) | ( ~n15314 & n15317 ) | ( n15316 & n15317 ) ;
  assign n15319 = n3541 & n11148 ;
  assign n15320 = x29 & n15319 ;
  assign n15321 = n3536 & n10259 ;
  assign n15322 = n4039 | n15321 ;
  assign n15323 = ( n10255 & n15321 ) | ( n10255 & n15322 ) | ( n15321 & n15322 ) ;
  assign n15324 = n3501 & n10257 ;
  assign n15325 = n15323 | n15324 ;
  assign n15326 = x29 & ~n15325 ;
  assign n15327 = ( ~x29 & n15319 ) | ( ~x29 & n15325 ) | ( n15319 & n15325 ) ;
  assign n15328 = ( ~n15320 & n15326 ) | ( ~n15320 & n15327 ) | ( n15326 & n15327 ) ;
  assign n15329 = n3273 & n10265 ;
  assign n15330 = n3270 | n15329 ;
  assign n15331 = ( n10261 & n15329 ) | ( n10261 & n15330 ) | ( n15329 & n15330 ) ;
  assign n15332 = n390 | n15331 ;
  assign n15333 = ( n11049 & n15331 ) | ( n11049 & n15332 ) | ( n15331 & n15332 ) ;
  assign n15334 = n3274 & n10263 ;
  assign n15335 = n15333 | n15334 ;
  assign n15336 = n14683 & ~n14887 ;
  assign n15337 = n13983 & ~n15133 ;
  assign n15338 = ( n13983 & ~n15336 ) | ( n13983 & n15337 ) | ( ~n15336 & n15337 ) ;
  assign n15339 = ~n14683 & n14887 ;
  assign n15340 = ~n13983 & n15133 ;
  assign n15341 = ( n13983 & n15339 ) | ( n13983 & ~n15340 ) | ( n15339 & ~n15340 ) ;
  assign n15342 = ( n14690 & n15338 ) | ( n14690 & n15341 ) | ( n15338 & n15341 ) ;
  assign n15343 = n3928 | n5661 ;
  assign n15344 = n287 | n362 ;
  assign n15345 = n15343 | n15344 ;
  assign n15346 = n5615 | n15345 ;
  assign n15347 = n3816 | n15346 ;
  assign n15348 = n680 | n3686 ;
  assign n15349 = n1144 | n15348 ;
  assign n15350 = n280 | n15349 ;
  assign n15351 = n5950 | n15350 ;
  assign n15352 = n15347 | n15351 ;
  assign n15353 = n1855 | n3021 ;
  assign n15354 = ~n2164 & n15126 ;
  assign n15355 = ~n15353 & n15354 ;
  assign n15356 = n289 | n455 ;
  assign n15357 = n226 | n15356 ;
  assign n15358 = n2653 | n15357 ;
  assign n15359 = n15355 & ~n15358 ;
  assign n15360 = ~n15352 & n15359 ;
  assign n15361 = ~n14866 & n15360 ;
  assign n15362 = ( ~n13983 & n14933 ) | ( ~n13983 & n15361 ) | ( n14933 & n15361 ) ;
  assign n15363 = ( n13983 & n14933 ) | ( n13983 & n15361 ) | ( n14933 & n15361 ) ;
  assign n15364 = ( n13983 & n15362 ) | ( n13983 & ~n15363 ) | ( n15362 & ~n15363 ) ;
  assign n15365 = ( n15335 & n15342 ) | ( n15335 & ~n15364 ) | ( n15342 & ~n15364 ) ;
  assign n15366 = ( n15335 & ~n15342 ) | ( n15335 & n15364 ) | ( ~n15342 & n15364 ) ;
  assign n15367 = ( ~n15335 & n15365 ) | ( ~n15335 & n15366 ) | ( n15365 & n15366 ) ;
  assign n15368 = ( n15145 & n15328 ) | ( n15145 & ~n15367 ) | ( n15328 & ~n15367 ) ;
  assign n15369 = ( n15145 & ~n15328 ) | ( n15145 & n15367 ) | ( ~n15328 & n15367 ) ;
  assign n15370 = ( ~n15145 & n15368 ) | ( ~n15145 & n15369 ) | ( n15368 & n15369 ) ;
  assign n15371 = ( ~n15158 & n15318 ) | ( ~n15158 & n15370 ) | ( n15318 & n15370 ) ;
  assign n15372 = ( n15158 & n15318 ) | ( n15158 & ~n15370 ) | ( n15318 & ~n15370 ) ;
  assign n15373 = ( ~n15318 & n15371 ) | ( ~n15318 & n15372 ) | ( n15371 & n15372 ) ;
  assign n15374 = ( n15162 & n15308 ) | ( n15162 & ~n15373 ) | ( n15308 & ~n15373 ) ;
  assign n15375 = ( n15162 & ~n15308 ) | ( n15162 & n15373 ) | ( ~n15308 & n15373 ) ;
  assign n15376 = ( ~n15162 & n15374 ) | ( ~n15162 & n15375 ) | ( n15374 & n15375 ) ;
  assign n15377 = ( n15164 & n15298 ) | ( n15164 & ~n15376 ) | ( n15298 & ~n15376 ) ;
  assign n15378 = ( n15164 & ~n15298 ) | ( n15164 & n15376 ) | ( ~n15298 & n15376 ) ;
  assign n15379 = ( ~n15164 & n15377 ) | ( ~n15164 & n15378 ) | ( n15377 & n15378 ) ;
  assign n15380 = ( ~n15168 & n15288 ) | ( ~n15168 & n15379 ) | ( n15288 & n15379 ) ;
  assign n15381 = ( n15168 & n15288 ) | ( n15168 & ~n15379 ) | ( n15288 & ~n15379 ) ;
  assign n15382 = ( ~n15288 & n15380 ) | ( ~n15288 & n15381 ) | ( n15380 & n15381 ) ;
  assign n15383 = ( n15171 & n15278 ) | ( n15171 & ~n15382 ) | ( n15278 & ~n15382 ) ;
  assign n15384 = ( n15171 & ~n15278 ) | ( n15171 & n15382 ) | ( ~n15278 & n15382 ) ;
  assign n15385 = ( ~n15171 & n15383 ) | ( ~n15171 & n15384 ) | ( n15383 & n15384 ) ;
  assign n15386 = ( n15173 & n15268 ) | ( n15173 & ~n15385 ) | ( n15268 & ~n15385 ) ;
  assign n15387 = ( n15173 & ~n15268 ) | ( n15173 & n15385 ) | ( ~n15268 & n15385 ) ;
  assign n15388 = ( ~n15173 & n15386 ) | ( ~n15173 & n15387 ) | ( n15386 & n15387 ) ;
  assign n15389 = ( n15176 & ~n15258 ) | ( n15176 & n15388 ) | ( ~n15258 & n15388 ) ;
  assign n15390 = ( n15176 & n15258 ) | ( n15176 & ~n15388 ) | ( n15258 & ~n15388 ) ;
  assign n15391 = ( ~n15176 & n15389 ) | ( ~n15176 & n15390 ) | ( n15389 & n15390 ) ;
  assign n15392 = ( ~n15179 & n15183 ) | ( ~n15179 & n15391 ) | ( n15183 & n15391 ) ;
  assign n15393 = ( n15179 & n15183 ) | ( n15179 & ~n15391 ) | ( n15183 & ~n15391 ) ;
  assign n15394 = ( ~n15183 & n15392 ) | ( ~n15183 & n15393 ) | ( n15392 & n15393 ) ;
  assign n15395 = n40 & ~n15394 ;
  assign n15396 = n8721 & ~n15184 ;
  assign n15397 = n8340 & n14942 ;
  assign n15398 = n15396 | n15397 ;
  assign n15399 = n15395 | n15398 ;
  assign n15400 = x5 & n15399 ;
  assign n15401 = ~n15184 & n15191 ;
  assign n15402 = n15394 & n15401 ;
  assign n15403 = ~n15193 & n15394 ;
  assign n15404 = ( n15193 & ~n15394 ) | ( n15193 & n15401 ) | ( ~n15394 & n15401 ) ;
  assign n15405 = ( ~n15402 & n15403 ) | ( ~n15402 & n15404 ) | ( n15403 & n15404 ) ;
  assign n15406 = n8341 & n15405 ;
  assign n15407 = ( ~x5 & n15399 ) | ( ~x5 & n15406 ) | ( n15399 & n15406 ) ;
  assign n15408 = x5 & ~n15406 ;
  assign n15409 = ( ~n15400 & n15407 ) | ( ~n15400 & n15408 ) | ( n15407 & n15408 ) ;
  assign n15410 = ( n15200 & n15249 ) | ( n15200 & n15409 ) | ( n15249 & n15409 ) ;
  assign n15411 = n6570 & ~n13473 ;
  assign n15412 = n6567 & ~n10235 ;
  assign n15413 = n15411 | n15412 ;
  assign n15414 = n6796 & ~n13280 ;
  assign n15415 = n15413 | n15414 ;
  assign n15416 = n6571 | n15415 ;
  assign n15417 = ( ~n13480 & n15415 ) | ( ~n13480 & n15416 ) | ( n15415 & n15416 ) ;
  assign n15418 = x11 & ~n15417 ;
  assign n15419 = ~x11 & n15417 ;
  assign n15420 = n15418 | n15419 ;
  assign n15421 = n5915 & n12953 ;
  assign n15422 = x14 & n15421 ;
  assign n15423 = n5909 & ~n10332 ;
  assign n15424 = n5914 | n15423 ;
  assign n15425 = ( n10214 & n15423 ) | ( n10214 & n15424 ) | ( n15423 & n15424 ) ;
  assign n15426 = n6332 & ~n10237 ;
  assign n15427 = n15425 | n15426 ;
  assign n15428 = x14 & ~n15427 ;
  assign n15429 = ( ~x14 & n15421 ) | ( ~x14 & n15427 ) | ( n15421 & n15427 ) ;
  assign n15430 = ( ~n15422 & n15428 ) | ( ~n15422 & n15429 ) | ( n15428 & n15429 ) ;
  assign n15431 = n5418 & n10397 ;
  assign n15432 = x17 & n15431 ;
  assign n15433 = n5413 & n10239 ;
  assign n15434 = n5417 | n15433 ;
  assign n15435 = ( n10329 & n15433 ) | ( n10329 & n15434 ) | ( n15433 & n15434 ) ;
  assign n15436 = n5584 & n10326 ;
  assign n15437 = n15435 | n15436 ;
  assign n15438 = x17 & ~n15437 ;
  assign n15439 = ( ~x17 & n15431 ) | ( ~x17 & n15437 ) | ( n15431 & n15437 ) ;
  assign n15440 = ( ~n15432 & n15438 ) | ( ~n15432 & n15439 ) | ( n15438 & n15439 ) ;
  assign n15441 = n5232 & n10243 ;
  assign n15442 = x20 & n15441 ;
  assign n15443 = n4874 & ~n10320 ;
  assign n15444 = n4878 | n15443 ;
  assign n15445 = ( n10241 & n15443 ) | ( n10241 & n15444 ) | ( n15443 & n15444 ) ;
  assign n15446 = n4879 | n15445 ;
  assign n15447 = ( n12105 & n15445 ) | ( n12105 & n15446 ) | ( n15445 & n15446 ) ;
  assign n15448 = x20 & ~n15447 ;
  assign n15449 = ( ~x20 & n15441 ) | ( ~x20 & n15447 ) | ( n15441 & n15447 ) ;
  assign n15450 = ( ~n15442 & n15448 ) | ( ~n15442 & n15449 ) | ( n15448 & n15449 ) ;
  assign n15451 = n4637 & ~n10316 ;
  assign n15452 = x23 & n15451 ;
  assign n15453 = n4584 & n10247 ;
  assign n15454 = n4649 | n15453 ;
  assign n15455 = ( n10245 & n15453 ) | ( n10245 & n15454 ) | ( n15453 & n15454 ) ;
  assign n15456 = n4591 | n15455 ;
  assign n15457 = ( ~n11676 & n15455 ) | ( ~n11676 & n15456 ) | ( n15455 & n15456 ) ;
  assign n15458 = x23 & ~n15457 ;
  assign n15459 = ( ~x23 & n15451 ) | ( ~x23 & n15457 ) | ( n15451 & n15457 ) ;
  assign n15460 = ( ~n15452 & n15458 ) | ( ~n15452 & n15459 ) | ( n15458 & n15459 ) ;
  assign n15461 = n4215 & n10312 ;
  assign n15462 = x26 & n15461 ;
  assign n15463 = n4200 & ~n10249 ;
  assign n15464 = n2083 & n10251 ;
  assign n15465 = n15463 | n15464 ;
  assign n15466 = n4203 | n15465 ;
  assign n15467 = ( ~n11486 & n15465 ) | ( ~n11486 & n15466 ) | ( n15465 & n15466 ) ;
  assign n15468 = x26 & ~n15467 ;
  assign n15469 = ( ~x26 & n15461 ) | ( ~x26 & n15467 ) | ( n15461 & n15467 ) ;
  assign n15470 = ( ~n15462 & n15468 ) | ( ~n15462 & n15469 ) | ( n15468 & n15469 ) ;
  assign n15471 = n3501 & n10255 ;
  assign n15472 = x29 & n15471 ;
  assign n15473 = n3536 & n10257 ;
  assign n15474 = n4039 | n15473 ;
  assign n15475 = ( ~n10253 & n15473 ) | ( ~n10253 & n15474 ) | ( n15473 & n15474 ) ;
  assign n15476 = n3541 | n15475 ;
  assign n15477 = ( ~n11297 & n15475 ) | ( ~n11297 & n15476 ) | ( n15475 & n15476 ) ;
  assign n15478 = x29 & ~n15477 ;
  assign n15479 = ( ~x29 & n15471 ) | ( ~x29 & n15477 ) | ( n15471 & n15477 ) ;
  assign n15480 = ( ~n15472 & n15478 ) | ( ~n15472 & n15479 ) | ( n15478 & n15479 ) ;
  assign n15481 = n3273 & n10263 ;
  assign n15482 = n3270 | n15481 ;
  assign n15483 = ( n10259 & n15481 ) | ( n10259 & n15482 ) | ( n15481 & n15482 ) ;
  assign n15484 = n390 | n15483 ;
  assign n15485 = ( n10859 & n15483 ) | ( n10859 & n15484 ) | ( n15483 & n15484 ) ;
  assign n15486 = n3274 & n10261 ;
  assign n15487 = n15485 | n15486 ;
  assign n15488 = n1148 | n1816 ;
  assign n15489 = n2470 | n15488 ;
  assign n15490 = n701 | n850 ;
  assign n15491 = n408 | n15490 ;
  assign n15492 = n15489 | n15491 ;
  assign n15493 = n2851 | n3868 ;
  assign n15494 = n15492 | n15493 ;
  assign n15495 = n902 | n1022 ;
  assign n15496 = n361 | n15495 ;
  assign n15497 = n15494 | n15496 ;
  assign n15498 = n185 | n215 ;
  assign n15499 = n844 | n15498 ;
  assign n15500 = n1167 | n15499 ;
  assign n15501 = n46 & n102 ;
  assign n15502 = n589 | n15501 ;
  assign n15503 = n662 | n15502 ;
  assign n15504 = n5612 | n15503 ;
  assign n15505 = n570 | n1786 ;
  assign n15506 = n15504 | n15505 ;
  assign n15507 = n15500 | n15506 ;
  assign n15508 = n15497 | n15507 ;
  assign n15509 = n2819 | n15508 ;
  assign n15510 = n956 | n4271 ;
  assign n15511 = n808 | n2074 ;
  assign n15512 = n15510 | n15511 ;
  assign n15513 = n704 | n13615 ;
  assign n15514 = n15512 | n15513 ;
  assign n15515 = n1887 | n2263 ;
  assign n15516 = n1226 | n15515 ;
  assign n15517 = n191 | n268 ;
  assign n15518 = n1365 | n15517 ;
  assign n15519 = n15516 | n15518 ;
  assign n15520 = n381 | n3116 ;
  assign n15521 = n4276 | n15520 ;
  assign n15522 = n4959 | n15521 ;
  assign n15523 = n15519 | n15522 ;
  assign n15524 = n15514 | n15523 ;
  assign n15525 = n15509 | n15524 ;
  assign n15526 = ( n15363 & ~n15487 ) | ( n15363 & n15525 ) | ( ~n15487 & n15525 ) ;
  assign n15527 = ( n15363 & n15487 ) | ( n15363 & n15525 ) | ( n15487 & n15525 ) ;
  assign n15528 = ( n15487 & n15526 ) | ( n15487 & ~n15527 ) | ( n15526 & ~n15527 ) ;
  assign n15529 = ( n15365 & ~n15480 ) | ( n15365 & n15528 ) | ( ~n15480 & n15528 ) ;
  assign n15530 = ( n15365 & n15480 ) | ( n15365 & n15528 ) | ( n15480 & n15528 ) ;
  assign n15531 = ( n15480 & n15529 ) | ( n15480 & ~n15530 ) | ( n15529 & ~n15530 ) ;
  assign n15532 = ( n15368 & ~n15470 ) | ( n15368 & n15531 ) | ( ~n15470 & n15531 ) ;
  assign n15533 = ( n15368 & n15470 ) | ( n15368 & n15531 ) | ( n15470 & n15531 ) ;
  assign n15534 = ( n15470 & n15532 ) | ( n15470 & ~n15533 ) | ( n15532 & ~n15533 ) ;
  assign n15535 = ( n15372 & n15460 ) | ( n15372 & n15534 ) | ( n15460 & n15534 ) ;
  assign n15536 = ( n15372 & ~n15460 ) | ( n15372 & n15534 ) | ( ~n15460 & n15534 ) ;
  assign n15537 = ( n15460 & ~n15535 ) | ( n15460 & n15536 ) | ( ~n15535 & n15536 ) ;
  assign n15538 = ( n15374 & ~n15450 ) | ( n15374 & n15537 ) | ( ~n15450 & n15537 ) ;
  assign n15539 = ( n15374 & n15450 ) | ( n15374 & n15537 ) | ( n15450 & n15537 ) ;
  assign n15540 = ( n15450 & n15538 ) | ( n15450 & ~n15539 ) | ( n15538 & ~n15539 ) ;
  assign n15541 = ( n15377 & n15440 ) | ( n15377 & n15540 ) | ( n15440 & n15540 ) ;
  assign n15542 = ( n15377 & ~n15440 ) | ( n15377 & n15540 ) | ( ~n15440 & n15540 ) ;
  assign n15543 = ( n15440 & ~n15541 ) | ( n15440 & n15542 ) | ( ~n15541 & n15542 ) ;
  assign n15544 = ( ~n15381 & n15430 ) | ( ~n15381 & n15543 ) | ( n15430 & n15543 ) ;
  assign n15545 = ( n15381 & n15430 ) | ( n15381 & n15543 ) | ( n15430 & n15543 ) ;
  assign n15546 = ( n15381 & n15544 ) | ( n15381 & ~n15545 ) | ( n15544 & ~n15545 ) ;
  assign n15547 = ( n15383 & ~n15420 ) | ( n15383 & n15546 ) | ( ~n15420 & n15546 ) ;
  assign n15548 = ( n15383 & n15420 ) | ( n15383 & n15546 ) | ( n15420 & n15546 ) ;
  assign n15549 = ( n15420 & n15547 ) | ( n15420 & ~n15548 ) | ( n15547 & ~n15548 ) ;
  assign n15550 = ( x5 & ~x6 ) | ( x5 & x7 ) | ( ~x6 & x7 ) ;
  assign n15551 = ( x6 & ~x8 ) | ( x6 & n15550 ) | ( ~x8 & n15550 ) ;
  assign n15552 = ~n7340 & n15551 ;
  assign n15553 = ( n13475 & n15551 ) | ( n13475 & n15552 ) | ( n15551 & n15552 ) ;
  assign n15554 = n7337 & ~n13475 ;
  assign n15555 = n15553 | n15554 ;
  assign n15556 = ( n15386 & n15549 ) | ( n15386 & n15555 ) | ( n15549 & n15555 ) ;
  assign n15557 = ( n15386 & ~n15549 ) | ( n15386 & n15555 ) | ( ~n15549 & n15555 ) ;
  assign n15558 = ( n15549 & ~n15556 ) | ( n15549 & n15557 ) | ( ~n15556 & n15557 ) ;
  assign n15559 = ( n15390 & ~n15393 ) | ( n15390 & n15558 ) | ( ~n15393 & n15558 ) ;
  assign n15560 = ( n15390 & n15393 ) | ( n15390 & n15558 ) | ( n15393 & n15558 ) ;
  assign n15561 = ( n15393 & n15559 ) | ( n15393 & ~n15560 ) | ( n15559 & ~n15560 ) ;
  assign n15562 = n40 & n15561 ;
  assign n15563 = n8721 & ~n15394 ;
  assign n15564 = n8340 & ~n15184 ;
  assign n15565 = n15563 | n15564 ;
  assign n15566 = n15562 | n15565 ;
  assign n15567 = x5 & n15566 ;
  assign n15568 = n15193 | n15394 ;
  assign n15569 = n15561 & ~n15568 ;
  assign n15570 = n15394 & ~n15401 ;
  assign n15571 = ( n15561 & n15568 ) | ( n15561 & ~n15570 ) | ( n15568 & ~n15570 ) ;
  assign n15572 = n15561 & ~n15570 ;
  assign n15573 = ( n15569 & n15571 ) | ( n15569 & ~n15572 ) | ( n15571 & ~n15572 ) ;
  assign n15574 = n8341 & n15573 ;
  assign n15575 = ( ~x5 & n15566 ) | ( ~x5 & n15574 ) | ( n15566 & n15574 ) ;
  assign n15576 = x5 & ~n15574 ;
  assign n15577 = ( ~n15567 & n15575 ) | ( ~n15567 & n15576 ) | ( n15575 & n15576 ) ;
  assign n15578 = n7644 & ~n14723 ;
  assign n15579 = x8 & n15578 ;
  assign n15580 = n7341 & n14520 ;
  assign n15581 = n7345 | n15580 ;
  assign n15582 = ( n14942 & n15580 ) | ( n14942 & n15581 ) | ( n15580 & n15581 ) ;
  assign n15583 = n7346 | n15582 ;
  assign n15584 = ( ~n14953 & n15582 ) | ( ~n14953 & n15583 ) | ( n15582 & n15583 ) ;
  assign n15585 = x8 & ~n15584 ;
  assign n15586 = ( ~x8 & n15578 ) | ( ~x8 & n15584 ) | ( n15578 & n15584 ) ;
  assign n15587 = ( ~n15579 & n15585 ) | ( ~n15579 & n15586 ) | ( n15585 & n15586 ) ;
  assign n15588 = n6796 & n13992 ;
  assign n15589 = x11 & n15588 ;
  assign n15590 = n6567 & n13996 ;
  assign n15591 = n6570 | n15590 ;
  assign n15592 = ( n14352 & n15590 ) | ( n14352 & n15591 ) | ( n15590 & n15591 ) ;
  assign n15593 = n6571 | n15592 ;
  assign n15594 = ( n14363 & n15592 ) | ( n14363 & n15593 ) | ( n15592 & n15593 ) ;
  assign n15595 = x11 & ~n15594 ;
  assign n15596 = ( ~x11 & n15588 ) | ( ~x11 & n15594 ) | ( n15588 & n15594 ) ;
  assign n15597 = ( ~n15589 & n15595 ) | ( ~n15589 & n15596 ) | ( n15595 & n15596 ) ;
  assign n15598 = n6332 & ~n14000 ;
  assign n15599 = x14 & n15598 ;
  assign n15600 = n5909 & ~n14007 ;
  assign n15601 = n5914 | n15600 ;
  assign n15602 = ( n13998 & n15600 ) | ( n13998 & n15601 ) | ( n15600 & n15601 ) ;
  assign n15603 = n5915 | n15602 ;
  assign n15604 = ( n14115 & n15602 ) | ( n14115 & n15603 ) | ( n15602 & n15603 ) ;
  assign n15605 = x14 & ~n15604 ;
  assign n15606 = ( ~x14 & n15598 ) | ( ~x14 & n15604 ) | ( n15598 & n15604 ) ;
  assign n15607 = ( ~n15599 & n15605 ) | ( ~n15599 & n15606 ) | ( n15605 & n15606 ) ;
  assign n15608 = x17 & ~n15029 ;
  assign n15609 = ~n15236 & n15608 ;
  assign n15610 = x17 & ~n15609 ;
  assign n15611 = n5584 & ~n14004 ;
  assign n15612 = n5413 & ~n14014 ;
  assign n15613 = n15611 | n15612 ;
  assign n15614 = n5418 | n15613 ;
  assign n15615 = ( n14072 & n15613 ) | ( n14072 & n15614 ) | ( n15613 & n15614 ) ;
  assign n15616 = n5417 & n14002 ;
  assign n15617 = n15615 | n15616 ;
  assign n15618 = n15610 & ~n15617 ;
  assign n15619 = ~n15610 & n15617 ;
  assign n15620 = n15618 | n15619 ;
  assign n15621 = ( ~n15241 & n15607 ) | ( ~n15241 & n15620 ) | ( n15607 & n15620 ) ;
  assign n15622 = ( n15241 & n15607 ) | ( n15241 & n15620 ) | ( n15607 & n15620 ) ;
  assign n15623 = ( n15241 & n15621 ) | ( n15241 & ~n15622 ) | ( n15621 & ~n15622 ) ;
  assign n15624 = ( ~n15245 & n15597 ) | ( ~n15245 & n15623 ) | ( n15597 & n15623 ) ;
  assign n15625 = ( n15245 & n15597 ) | ( n15245 & n15623 ) | ( n15597 & n15623 ) ;
  assign n15626 = ( n15245 & n15624 ) | ( n15245 & ~n15625 ) | ( n15624 & ~n15625 ) ;
  assign n15627 = ( ~n15247 & n15587 ) | ( ~n15247 & n15626 ) | ( n15587 & n15626 ) ;
  assign n15628 = ( n15247 & n15587 ) | ( n15247 & n15626 ) | ( n15587 & n15626 ) ;
  assign n15629 = ( n15247 & n15627 ) | ( n15247 & ~n15628 ) | ( n15627 & ~n15628 ) ;
  assign n15630 = ( n15410 & n15577 ) | ( n15410 & n15629 ) | ( n15577 & n15629 ) ;
  assign n15631 = n7644 & n14942 ;
  assign n15632 = x8 & n15631 ;
  assign n15633 = n7341 & ~n14723 ;
  assign n15634 = n7345 | n15633 ;
  assign n15635 = ( ~n15184 & n15633 ) | ( ~n15184 & n15634 ) | ( n15633 & n15634 ) ;
  assign n15636 = n7346 | n15635 ;
  assign n15637 = ( ~n15195 & n15635 ) | ( ~n15195 & n15636 ) | ( n15635 & n15636 ) ;
  assign n15638 = x8 & ~n15637 ;
  assign n15639 = ( ~x8 & n15631 ) | ( ~x8 & n15637 ) | ( n15631 & n15637 ) ;
  assign n15640 = ( ~n15632 & n15638 ) | ( ~n15632 & n15639 ) | ( n15638 & n15639 ) ;
  assign n15641 = n6570 & n14520 ;
  assign n15642 = n6571 | n15641 ;
  assign n15643 = ( n14531 & n15641 ) | ( n14531 & n15642 ) | ( n15641 & n15642 ) ;
  assign n15644 = n6567 & n13992 ;
  assign n15645 = ( ~x11 & n15643 ) | ( ~x11 & n15644 ) | ( n15643 & n15644 ) ;
  assign n15646 = n6796 & n14352 ;
  assign n15647 = x11 & ~n15644 ;
  assign n15648 = n15646 | n15647 ;
  assign n15649 = ( n15643 & n15646 ) | ( n15643 & n15647 ) | ( n15646 & n15647 ) ;
  assign n15650 = ( n15645 & n15648 ) | ( n15645 & ~n15649 ) | ( n15648 & ~n15649 ) ;
  assign n15651 = n5915 & ~n14130 ;
  assign n15652 = x14 & n15651 ;
  assign n15653 = n5909 & ~n14000 ;
  assign n15654 = n5914 | n15653 ;
  assign n15655 = ( n13996 & n15653 ) | ( n13996 & n15654 ) | ( n15653 & n15654 ) ;
  assign n15656 = n6332 & n13998 ;
  assign n15657 = n15655 | n15656 ;
  assign n15658 = x14 & ~n15657 ;
  assign n15659 = ( ~x14 & n15651 ) | ( ~x14 & n15657 ) | ( n15651 & n15657 ) ;
  assign n15660 = ( ~n15652 & n15658 ) | ( ~n15652 & n15659 ) | ( n15658 & n15659 ) ;
  assign n15661 = n15609 & ~n15617 ;
  assign n15662 = n5584 & n14002 ;
  assign n15663 = x17 & n15662 ;
  assign n15664 = n5413 & ~n14004 ;
  assign n15665 = n5417 | n15664 ;
  assign n15666 = ( ~n14007 & n15664 ) | ( ~n14007 & n15665 ) | ( n15664 & n15665 ) ;
  assign n15667 = n5418 | n15666 ;
  assign n15668 = ( n14066 & n15666 ) | ( n14066 & n15667 ) | ( n15666 & n15667 ) ;
  assign n15669 = x17 & ~n15668 ;
  assign n15670 = ( ~x17 & n15662 ) | ( ~x17 & n15668 ) | ( n15662 & n15668 ) ;
  assign n15671 = ( ~n15663 & n15669 ) | ( ~n15663 & n15670 ) | ( n15669 & n15670 ) ;
  assign n15672 = n4875 & ~n14014 ;
  assign n15673 = n15661 | n15672 ;
  assign n15674 = n15671 & n15673 ;
  assign n15675 = ( ~n15661 & n15671 ) | ( ~n15661 & n15672 ) | ( n15671 & n15672 ) ;
  assign n15676 = ( n15661 & ~n15674 ) | ( n15661 & n15675 ) | ( ~n15674 & n15675 ) ;
  assign n15677 = ( ~n15622 & n15660 ) | ( ~n15622 & n15676 ) | ( n15660 & n15676 ) ;
  assign n15678 = ( n15622 & n15660 ) | ( n15622 & n15676 ) | ( n15660 & n15676 ) ;
  assign n15679 = ( n15622 & n15677 ) | ( n15622 & ~n15678 ) | ( n15677 & ~n15678 ) ;
  assign n15680 = ( n15625 & ~n15650 ) | ( n15625 & n15679 ) | ( ~n15650 & n15679 ) ;
  assign n15681 = ( n15625 & n15650 ) | ( n15625 & n15679 ) | ( n15650 & n15679 ) ;
  assign n15682 = ( n15650 & n15680 ) | ( n15650 & ~n15681 ) | ( n15680 & ~n15681 ) ;
  assign n15683 = ( ~n15628 & n15640 ) | ( ~n15628 & n15682 ) | ( n15640 & n15682 ) ;
  assign n15684 = ( n15628 & n15640 ) | ( n15628 & n15682 ) | ( n15640 & n15682 ) ;
  assign n15685 = ( n15628 & n15683 ) | ( n15628 & ~n15684 ) | ( n15683 & ~n15684 ) ;
  assign n15686 = n6567 & ~n13280 ;
  assign n15687 = n6570 | n15686 ;
  assign n15688 = ( n13475 & n15686 ) | ( n13475 & n15687 ) | ( n15686 & n15687 ) ;
  assign n15689 = n6796 & ~n13473 ;
  assign n15690 = n15688 | n15689 ;
  assign n15691 = x11 & n15690 ;
  assign n15692 = n6571 & n13671 ;
  assign n15693 = ( ~x11 & n15690 ) | ( ~x11 & n15692 ) | ( n15690 & n15692 ) ;
  assign n15694 = x11 & ~n15692 ;
  assign n15695 = ( ~n15691 & n15693 ) | ( ~n15691 & n15694 ) | ( n15693 & n15694 ) ;
  assign n15696 = n5909 & ~n10237 ;
  assign n15697 = n5914 | n15696 ;
  assign n15698 = ( ~n10235 & n15696 ) | ( ~n10235 & n15697 ) | ( n15696 & n15697 ) ;
  assign n15699 = n6332 & n10214 ;
  assign n15700 = n15698 | n15699 ;
  assign n15701 = x14 & n15700 ;
  assign n15702 = n5915 & n10371 ;
  assign n15703 = x14 & ~n15702 ;
  assign n15704 = ( ~x14 & n15700 ) | ( ~x14 & n15702 ) | ( n15700 & n15702 ) ;
  assign n15705 = ( ~n15701 & n15703 ) | ( ~n15701 & n15704 ) | ( n15703 & n15704 ) ;
  assign n15706 = n5584 & n10329 ;
  assign n15707 = x17 & n15706 ;
  assign n15708 = n5413 & n10326 ;
  assign n15709 = n5417 | n15708 ;
  assign n15710 = ( ~n10332 & n15708 ) | ( ~n10332 & n15709 ) | ( n15708 & n15709 ) ;
  assign n15711 = n5418 | n15710 ;
  assign n15712 = ( ~n10383 & n15710 ) | ( ~n10383 & n15711 ) | ( n15710 & n15711 ) ;
  assign n15713 = x17 & ~n15712 ;
  assign n15714 = ( ~x17 & n15706 ) | ( ~x17 & n15712 ) | ( n15706 & n15712 ) ;
  assign n15715 = ( ~n15707 & n15713 ) | ( ~n15707 & n15714 ) | ( n15713 & n15714 ) ;
  assign n15716 = n4879 & n12575 ;
  assign n15717 = x20 & n15716 ;
  assign n15718 = n4874 & n10243 ;
  assign n15719 = n4878 | n15718 ;
  assign n15720 = ( n10239 & n15718 ) | ( n10239 & n15719 ) | ( n15718 & n15719 ) ;
  assign n15721 = n5232 & n10241 ;
  assign n15722 = n15720 | n15721 ;
  assign n15723 = x20 & ~n15722 ;
  assign n15724 = ( ~x20 & n15716 ) | ( ~x20 & n15722 ) | ( n15716 & n15722 ) ;
  assign n15725 = ( ~n15717 & n15723 ) | ( ~n15717 & n15724 ) | ( n15723 & n15724 ) ;
  assign n15726 = n4649 & ~n10320 ;
  assign n15727 = x23 & n15726 ;
  assign n15728 = n4637 & n10245 ;
  assign n15729 = n4584 & ~n10316 ;
  assign n15730 = n15728 | n15729 ;
  assign n15731 = n4591 | n15730 ;
  assign n15732 = ( ~n10414 & n15730 ) | ( ~n10414 & n15731 ) | ( n15730 & n15731 ) ;
  assign n15733 = x23 & ~n15732 ;
  assign n15734 = ( ~x23 & n15726 ) | ( ~x23 & n15732 ) | ( n15726 & n15732 ) ;
  assign n15735 = ( ~n15727 & n15733 ) | ( ~n15727 & n15734 ) | ( n15733 & n15734 ) ;
  assign n15736 = n4203 & n10428 ;
  assign n15737 = n4215 & n10247 ;
  assign n15738 = n4200 & n10312 ;
  assign n15739 = n2083 & ~n10249 ;
  assign n15740 = n15738 | n15739 ;
  assign n15741 = n15737 | n15740 ;
  assign n15742 = n15736 | n15741 ;
  assign n15743 = n4039 & n10251 ;
  assign n15744 = n3541 | n15743 ;
  assign n15745 = ( ~n11309 & n15743 ) | ( ~n11309 & n15744 ) | ( n15743 & n15744 ) ;
  assign n15746 = n3501 & ~n10253 ;
  assign n15747 = n15745 | n15746 ;
  assign n15748 = n3536 & n10255 ;
  assign n15749 = n15747 | n15748 ;
  assign n15750 = ( x26 & ~x29 ) | ( x26 & n15747 ) | ( ~x29 & n15747 ) ;
  assign n15751 = ( ~x26 & x29 ) | ( ~x26 & n15747 ) | ( x29 & n15747 ) ;
  assign n15752 = ( ~n15749 & n15750 ) | ( ~n15749 & n15751 ) | ( n15750 & n15751 ) ;
  assign n15753 = n1139 | n2549 ;
  assign n15754 = n313 | n434 ;
  assign n15755 = n470 | n15754 ;
  assign n15756 = n15753 | n15755 ;
  assign n15757 = n822 | n15756 ;
  assign n15758 = n755 | n15757 ;
  assign n15759 = n44 | n71 ;
  assign n15760 = n84 & n15759 ;
  assign n15761 = n4425 | n15760 ;
  assign n15762 = n2611 | n15761 ;
  assign n15763 = n269 | n432 ;
  assign n15764 = n1745 | n15763 ;
  assign n15765 = n5051 | n15764 ;
  assign n15766 = n15762 | n15765 ;
  assign n15767 = n15758 | n15766 ;
  assign n15768 = n2361 | n15767 ;
  assign n15769 = n2464 & ~n15768 ;
  assign n15770 = ( n15525 & n15526 ) | ( n15525 & n15769 ) | ( n15526 & n15769 ) ;
  assign n15771 = ( ~n15525 & n15526 ) | ( ~n15525 & n15769 ) | ( n15526 & n15769 ) ;
  assign n15772 = ( n15525 & ~n15770 ) | ( n15525 & n15771 ) | ( ~n15770 & n15771 ) ;
  assign n15773 = n3273 & n10261 ;
  assign n15774 = n3270 | n15773 ;
  assign n15775 = ( n10257 & n15773 ) | ( n10257 & n15774 ) | ( n15773 & n15774 ) ;
  assign n15776 = n390 | n15775 ;
  assign n15777 = ( n11065 & n15775 ) | ( n11065 & n15776 ) | ( n15775 & n15776 ) ;
  assign n15778 = n3274 & n10259 ;
  assign n15779 = n15777 | n15778 ;
  assign n15780 = ( n15530 & n15772 ) | ( n15530 & n15779 ) | ( n15772 & n15779 ) ;
  assign n15781 = ( n15530 & ~n15772 ) | ( n15530 & n15779 ) | ( ~n15772 & n15779 ) ;
  assign n15782 = ( n15772 & ~n15780 ) | ( n15772 & n15781 ) | ( ~n15780 & n15781 ) ;
  assign n15783 = ( ~n15742 & n15752 ) | ( ~n15742 & n15782 ) | ( n15752 & n15782 ) ;
  assign n15784 = ( n15742 & n15752 ) | ( n15742 & n15782 ) | ( n15752 & n15782 ) ;
  assign n15785 = ( n15742 & n15783 ) | ( n15742 & ~n15784 ) | ( n15783 & ~n15784 ) ;
  assign n15786 = ( n15533 & n15735 ) | ( n15533 & ~n15785 ) | ( n15735 & ~n15785 ) ;
  assign n15787 = ( ~n15533 & n15735 ) | ( ~n15533 & n15785 ) | ( n15735 & n15785 ) ;
  assign n15788 = ( ~n15735 & n15786 ) | ( ~n15735 & n15787 ) | ( n15786 & n15787 ) ;
  assign n15789 = ( ~n15535 & n15725 ) | ( ~n15535 & n15788 ) | ( n15725 & n15788 ) ;
  assign n15790 = ( n15535 & n15725 ) | ( n15535 & ~n15788 ) | ( n15725 & ~n15788 ) ;
  assign n15791 = ( ~n15725 & n15789 ) | ( ~n15725 & n15790 ) | ( n15789 & n15790 ) ;
  assign n15792 = ( ~n15539 & n15715 ) | ( ~n15539 & n15791 ) | ( n15715 & n15791 ) ;
  assign n15793 = ( n15539 & n15715 ) | ( n15539 & ~n15791 ) | ( n15715 & ~n15791 ) ;
  assign n15794 = ( ~n15715 & n15792 ) | ( ~n15715 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = ( n15541 & n15705 ) | ( n15541 & ~n15794 ) | ( n15705 & ~n15794 ) ;
  assign n15796 = ( ~n15541 & n15705 ) | ( ~n15541 & n15794 ) | ( n15705 & n15794 ) ;
  assign n15797 = ( ~n15705 & n15795 ) | ( ~n15705 & n15796 ) | ( n15795 & n15796 ) ;
  assign n15798 = ( n15545 & n15695 ) | ( n15545 & ~n15797 ) | ( n15695 & ~n15797 ) ;
  assign n15799 = ( ~n15545 & n15695 ) | ( ~n15545 & n15797 ) | ( n15695 & n15797 ) ;
  assign n15800 = ( ~n15695 & n15798 ) | ( ~n15695 & n15799 ) | ( n15798 & n15799 ) ;
  assign n15801 = ( n15548 & n15551 ) | ( n15548 & ~n15800 ) | ( n15551 & ~n15800 ) ;
  assign n15802 = ( n15548 & ~n15551 ) | ( n15548 & n15800 ) | ( ~n15551 & n15800 ) ;
  assign n15803 = ( ~n15548 & n15801 ) | ( ~n15548 & n15802 ) | ( n15801 & n15802 ) ;
  assign n15804 = ( ~n15556 & n15560 ) | ( ~n15556 & n15803 ) | ( n15560 & n15803 ) ;
  assign n15805 = ( n15556 & n15560 ) | ( n15556 & ~n15803 ) | ( n15560 & ~n15803 ) ;
  assign n15806 = ( ~n15560 & n15804 ) | ( ~n15560 & n15805 ) | ( n15804 & n15805 ) ;
  assign n15807 = n40 & ~n15806 ;
  assign n15808 = n8721 & n15561 ;
  assign n15809 = n8340 & ~n15394 ;
  assign n15810 = n15808 | n15809 ;
  assign n15811 = n15807 | n15810 ;
  assign n15812 = x5 & n15811 ;
  assign n15813 = n15572 & ~n15806 ;
  assign n15814 = ~n15561 & n15568 ;
  assign n15815 = n15806 | n15814 ;
  assign n15816 = ( n15572 & n15806 ) | ( n15572 & n15814 ) | ( n15806 & n15814 ) ;
  assign n15817 = ( n15813 & n15815 ) | ( n15813 & ~n15816 ) | ( n15815 & ~n15816 ) ;
  assign n15818 = n8341 & n15817 ;
  assign n15819 = ( ~x5 & n15811 ) | ( ~x5 & n15818 ) | ( n15811 & n15818 ) ;
  assign n15820 = x5 & ~n15818 ;
  assign n15821 = ( ~n15812 & n15819 ) | ( ~n15812 & n15820 ) | ( n15819 & n15820 ) ;
  assign n15822 = ( n15630 & n15685 ) | ( n15630 & n15821 ) | ( n15685 & n15821 ) ;
  assign n15823 = n6332 & ~n10235 ;
  assign n15824 = x14 & n15823 ;
  assign n15825 = n5909 & n10214 ;
  assign n15826 = n5914 | n15825 ;
  assign n15827 = ( ~n13280 & n15825 ) | ( ~n13280 & n15826 ) | ( n15825 & n15826 ) ;
  assign n15828 = n5915 | n15827 ;
  assign n15829 = ( ~n13285 & n15827 ) | ( ~n13285 & n15828 ) | ( n15827 & n15828 ) ;
  assign n15830 = x14 & ~n15829 ;
  assign n15831 = ( ~x14 & n15823 ) | ( ~x14 & n15829 ) | ( n15823 & n15829 ) ;
  assign n15832 = ( ~n15824 & n15830 ) | ( ~n15824 & n15831 ) | ( n15830 & n15831 ) ;
  assign n15833 = n5418 & n12756 ;
  assign n15834 = x17 & n15833 ;
  assign n15835 = n5417 & ~n10237 ;
  assign n15836 = n5584 & ~n10332 ;
  assign n15837 = n5413 & n10329 ;
  assign n15838 = n15836 | n15837 ;
  assign n15839 = n15835 | n15838 ;
  assign n15840 = x17 & ~n15839 ;
  assign n15841 = ( ~x17 & n15833 ) | ( ~x17 & n15839 ) | ( n15833 & n15839 ) ;
  assign n15842 = ( ~n15834 & n15840 ) | ( ~n15834 & n15841 ) | ( n15840 & n15841 ) ;
  assign n15843 = n5232 & n10239 ;
  assign n15844 = x20 & n15843 ;
  assign n15845 = n4874 & n10241 ;
  assign n15846 = n4878 | n15845 ;
  assign n15847 = ( n10326 & n15845 ) | ( n10326 & n15846 ) | ( n15845 & n15846 ) ;
  assign n15848 = n4879 | n15847 ;
  assign n15849 = ( n12222 & n15847 ) | ( n12222 & n15848 ) | ( n15847 & n15848 ) ;
  assign n15850 = x20 & ~n15849 ;
  assign n15851 = ( ~x20 & n15843 ) | ( ~x20 & n15849 ) | ( n15843 & n15849 ) ;
  assign n15852 = ( ~n15844 & n15850 ) | ( ~n15844 & n15851 ) | ( n15850 & n15851 ) ;
  assign n15853 = n4591 & ~n11989 ;
  assign n15854 = x23 & n15853 ;
  assign n15855 = n4649 & n10243 ;
  assign n15856 = n4637 & ~n10320 ;
  assign n15857 = n4584 & n10245 ;
  assign n15858 = n15856 | n15857 ;
  assign n15859 = n15855 | n15858 ;
  assign n15860 = x23 & ~n15859 ;
  assign n15861 = ( ~x23 & n15853 ) | ( ~x23 & n15859 ) | ( n15853 & n15859 ) ;
  assign n15862 = ( ~n15854 & n15860 ) | ( ~n15854 & n15861 ) | ( n15860 & n15861 ) ;
  assign n15863 = n4215 & ~n10316 ;
  assign n15864 = n4200 & n10247 ;
  assign n15865 = n2083 & n10312 ;
  assign n15866 = n15864 | n15865 ;
  assign n15867 = n15863 | n15866 ;
  assign n15868 = x26 & n15867 ;
  assign n15869 = n4203 & ~n11691 ;
  assign n15870 = ( ~x26 & n15867 ) | ( ~x26 & n15869 ) | ( n15867 & n15869 ) ;
  assign n15871 = x26 & ~n15869 ;
  assign n15872 = ( ~n15868 & n15870 ) | ( ~n15868 & n15871 ) | ( n15870 & n15871 ) ;
  assign n15873 = x26 & ~n15742 ;
  assign n15874 = ~x26 & n15742 ;
  assign n15875 = n15873 | n15874 ;
  assign n15876 = x29 & ~n15749 ;
  assign n15877 = ~x29 & n15749 ;
  assign n15878 = n15876 | n15877 ;
  assign n15879 = ( ~n15782 & n15875 ) | ( ~n15782 & n15878 ) | ( n15875 & n15878 ) ;
  assign n15880 = n3501 & n10251 ;
  assign n15881 = x29 & n15880 ;
  assign n15882 = n3536 & ~n10253 ;
  assign n15883 = n4039 | n15882 ;
  assign n15884 = ( ~n10249 & n15882 ) | ( ~n10249 & n15883 ) | ( n15882 & n15883 ) ;
  assign n15885 = n3541 | n15884 ;
  assign n15886 = ( ~n10441 & n15884 ) | ( ~n10441 & n15885 ) | ( n15884 & n15885 ) ;
  assign n15887 = x29 & ~n15886 ;
  assign n15888 = ( ~x29 & n15880 ) | ( ~x29 & n15886 ) | ( n15880 & n15886 ) ;
  assign n15889 = ( ~n15881 & n15887 ) | ( ~n15881 & n15888 ) | ( n15887 & n15888 ) ;
  assign n15890 = n3273 & n10259 ;
  assign n15891 = n3270 | n15890 ;
  assign n15892 = ( n10255 & n15890 ) | ( n10255 & n15891 ) | ( n15890 & n15891 ) ;
  assign n15893 = n390 | n15892 ;
  assign n15894 = ( n11148 & n15892 ) | ( n11148 & n15893 ) | ( n15892 & n15893 ) ;
  assign n15895 = n3274 & n10257 ;
  assign n15896 = n15894 | n15895 ;
  assign n15897 = ~n1790 & n13393 ;
  assign n15898 = n1319 | n2913 ;
  assign n15899 = n4892 | n6137 ;
  assign n15900 = n15898 | n15899 ;
  assign n15901 = n440 | n589 ;
  assign n15902 = n614 | n15901 ;
  assign n15903 = n1711 | n15902 ;
  assign n15904 = n4131 | n15903 ;
  assign n15905 = n2382 | n15904 ;
  assign n15906 = n15900 | n15905 ;
  assign n15907 = n80 | n742 ;
  assign n15908 = n364 | n15907 ;
  assign n15909 = n296 | n617 ;
  assign n15910 = n254 | n15909 ;
  assign n15911 = n223 | n15910 ;
  assign n15912 = n15908 | n15911 ;
  assign n15913 = n15906 | n15912 ;
  assign n15914 = n3398 | n15913 ;
  assign n15915 = n15897 & ~n15914 ;
  assign n15916 = ( n15525 & n15551 ) | ( n15525 & n15915 ) | ( n15551 & n15915 ) ;
  assign n15917 = ( ~n15525 & n15551 ) | ( ~n15525 & n15915 ) | ( n15551 & n15915 ) ;
  assign n15918 = ( n15525 & ~n15916 ) | ( n15525 & n15917 ) | ( ~n15916 & n15917 ) ;
  assign n15919 = ( n15770 & n15896 ) | ( n15770 & ~n15918 ) | ( n15896 & ~n15918 ) ;
  assign n15920 = ( ~n15770 & n15896 ) | ( ~n15770 & n15918 ) | ( n15896 & n15918 ) ;
  assign n15921 = ( ~n15896 & n15919 ) | ( ~n15896 & n15920 ) | ( n15919 & n15920 ) ;
  assign n15922 = ( n15781 & n15889 ) | ( n15781 & ~n15921 ) | ( n15889 & ~n15921 ) ;
  assign n15923 = ( ~n15781 & n15889 ) | ( ~n15781 & n15921 ) | ( n15889 & n15921 ) ;
  assign n15924 = ( ~n15889 & n15922 ) | ( ~n15889 & n15923 ) | ( n15922 & n15923 ) ;
  assign n15925 = ( n15872 & ~n15879 ) | ( n15872 & n15924 ) | ( ~n15879 & n15924 ) ;
  assign n15926 = ( n15872 & n15879 ) | ( n15872 & ~n15924 ) | ( n15879 & ~n15924 ) ;
  assign n15927 = ( ~n15872 & n15925 ) | ( ~n15872 & n15926 ) | ( n15925 & n15926 ) ;
  assign n15928 = ( n15786 & n15862 ) | ( n15786 & ~n15927 ) | ( n15862 & ~n15927 ) ;
  assign n15929 = ( n15786 & ~n15862 ) | ( n15786 & n15927 ) | ( ~n15862 & n15927 ) ;
  assign n15930 = ( ~n15786 & n15928 ) | ( ~n15786 & n15929 ) | ( n15928 & n15929 ) ;
  assign n15931 = ( n15790 & n15852 ) | ( n15790 & ~n15930 ) | ( n15852 & ~n15930 ) ;
  assign n15932 = ( n15790 & ~n15852 ) | ( n15790 & n15930 ) | ( ~n15852 & n15930 ) ;
  assign n15933 = ( ~n15790 & n15931 ) | ( ~n15790 & n15932 ) | ( n15931 & n15932 ) ;
  assign n15934 = ( n15793 & ~n15842 ) | ( n15793 & n15933 ) | ( ~n15842 & n15933 ) ;
  assign n15935 = ( n15793 & n15842 ) | ( n15793 & ~n15933 ) | ( n15842 & ~n15933 ) ;
  assign n15936 = ( ~n15793 & n15934 ) | ( ~n15793 & n15935 ) | ( n15934 & n15935 ) ;
  assign n15937 = ( n15795 & n15832 ) | ( n15795 & ~n15936 ) | ( n15832 & ~n15936 ) ;
  assign n15938 = ( n15795 & ~n15832 ) | ( n15795 & n15936 ) | ( ~n15832 & n15936 ) ;
  assign n15939 = ( ~n15795 & n15937 ) | ( ~n15795 & n15938 ) | ( n15937 & n15938 ) ;
  assign n15940 = n6567 | n6570 ;
  assign n15941 = ( n6570 & ~n13473 ) | ( n6570 & n15940 ) | ( ~n13473 & n15940 ) ;
  assign n15942 = n6796 | n15941 ;
  assign n15943 = ( n13475 & n15941 ) | ( n13475 & n15942 ) | ( n15941 & n15942 ) ;
  assign n15944 = x11 & n15943 ;
  assign n15945 = n6568 & n13477 ;
  assign n15946 = x11 & ~n15945 ;
  assign n15947 = ( ~x11 & n15943 ) | ( ~x11 & n15945 ) | ( n15943 & n15945 ) ;
  assign n15948 = ( ~n15944 & n15946 ) | ( ~n15944 & n15947 ) | ( n15946 & n15947 ) ;
  assign n15949 = ( n15798 & n15939 ) | ( n15798 & n15948 ) | ( n15939 & n15948 ) ;
  assign n15950 = ( n15798 & ~n15939 ) | ( n15798 & n15948 ) | ( ~n15939 & n15948 ) ;
  assign n15951 = ( n15939 & ~n15949 ) | ( n15939 & n15950 ) | ( ~n15949 & n15950 ) ;
  assign n15952 = ( n15801 & n15805 ) | ( n15801 & ~n15951 ) | ( n15805 & ~n15951 ) ;
  assign n15953 = ( ~n15801 & n15805 ) | ( ~n15801 & n15951 ) | ( n15805 & n15951 ) ;
  assign n15954 = ( ~n15805 & n15952 ) | ( ~n15805 & n15953 ) | ( n15952 & n15953 ) ;
  assign n15955 = n40 & ~n15954 ;
  assign n15956 = n8721 & ~n15806 ;
  assign n15957 = n8340 & n15561 ;
  assign n15958 = n15956 | n15957 ;
  assign n15959 = n15955 | n15958 ;
  assign n15960 = x5 & n15959 ;
  assign n15961 = ~n15572 & n15806 ;
  assign n15962 = n15954 & n15961 ;
  assign n15963 = n15815 & n15954 ;
  assign n15964 = ( n15815 & n15954 ) | ( n15815 & ~n15961 ) | ( n15954 & ~n15961 ) ;
  assign n15965 = ( n15962 & ~n15963 ) | ( n15962 & n15964 ) | ( ~n15963 & n15964 ) ;
  assign n15966 = n8341 & ~n15965 ;
  assign n15967 = ( ~x5 & n15959 ) | ( ~x5 & n15966 ) | ( n15959 & n15966 ) ;
  assign n15968 = x5 & ~n15966 ;
  assign n15969 = ( ~n15960 & n15967 ) | ( ~n15960 & n15968 ) | ( n15967 & n15968 ) ;
  assign n15970 = n7644 & ~n15184 ;
  assign n15971 = x8 & n15970 ;
  assign n15972 = n7341 & n14942 ;
  assign n15973 = n7345 | n15972 ;
  assign n15974 = ( ~n15394 & n15972 ) | ( ~n15394 & n15973 ) | ( n15972 & n15973 ) ;
  assign n15975 = n7346 | n15974 ;
  assign n15976 = ( n15405 & n15974 ) | ( n15405 & n15975 ) | ( n15974 & n15975 ) ;
  assign n15977 = x8 & ~n15976 ;
  assign n15978 = ( ~x8 & n15970 ) | ( ~x8 & n15976 ) | ( n15970 & n15976 ) ;
  assign n15979 = ( ~n15971 & n15977 ) | ( ~n15971 & n15978 ) | ( n15977 & n15978 ) ;
  assign n15980 = n6796 & n14520 ;
  assign n15981 = x11 & n15980 ;
  assign n15982 = n6567 & n14352 ;
  assign n15983 = n6570 | n15982 ;
  assign n15984 = ( ~n14723 & n15982 ) | ( ~n14723 & n15983 ) | ( n15982 & n15983 ) ;
  assign n15985 = n6571 | n15984 ;
  assign n15986 = ( ~n14734 & n15984 ) | ( ~n14734 & n15985 ) | ( n15984 & n15985 ) ;
  assign n15987 = x11 & ~n15986 ;
  assign n15988 = ( ~x11 & n15980 ) | ( ~x11 & n15986 ) | ( n15980 & n15986 ) ;
  assign n15989 = ( ~n15981 & n15987 ) | ( ~n15981 & n15988 ) | ( n15987 & n15988 ) ;
  assign n15990 = n5914 & n13992 ;
  assign n15991 = x14 & n15990 ;
  assign n15992 = n6332 & n13996 ;
  assign n15993 = n5909 & n13998 ;
  assign n15994 = n15992 | n15993 ;
  assign n15995 = n5915 | n15994 ;
  assign n15996 = ( n14024 & n15994 ) | ( n14024 & n15995 ) | ( n15994 & n15995 ) ;
  assign n15997 = x14 & ~n15996 ;
  assign n15998 = ( ~x14 & n15990 ) | ( ~x14 & n15996 ) | ( n15990 & n15996 ) ;
  assign n15999 = ( ~n15991 & n15997 ) | ( ~n15991 & n15998 ) | ( n15997 & n15998 ) ;
  assign n16000 = n5584 & ~n14007 ;
  assign n16001 = x17 & n16000 ;
  assign n16002 = n5413 & n14002 ;
  assign n16003 = n5417 | n16002 ;
  assign n16004 = ( ~n14000 & n16002 ) | ( ~n14000 & n16003 ) | ( n16002 & n16003 ) ;
  assign n16005 = n5418 | n16004 ;
  assign n16006 = ( ~n14042 & n16004 ) | ( ~n14042 & n16005 ) | ( n16004 & n16005 ) ;
  assign n16007 = x17 & ~n16006 ;
  assign n16008 = ( ~x17 & n16000 ) | ( ~x17 & n16006 ) | ( n16000 & n16006 ) ;
  assign n16009 = ( ~n16001 & n16007 ) | ( ~n16001 & n16008 ) | ( n16007 & n16008 ) ;
  assign n16010 = ( n5232 & n7364 ) | ( n5232 & n14004 ) | ( n7364 & n14004 ) ;
  assign n16011 = ~n14014 & n16010 ;
  assign n16012 = n4875 & n14015 ;
  assign n16013 = n16011 | n16012 ;
  assign n16014 = n4878 & ~n14004 ;
  assign n16015 = n16013 | n16014 ;
  assign n16016 = x20 & n15672 ;
  assign n16017 = ~n16015 & n16016 ;
  assign n16018 = n16015 & ~n16016 ;
  assign n16019 = n16017 | n16018 ;
  assign n16020 = ( n15674 & n16009 ) | ( n15674 & n16019 ) | ( n16009 & n16019 ) ;
  assign n16021 = ( n15674 & ~n16009 ) | ( n15674 & n16019 ) | ( ~n16009 & n16019 ) ;
  assign n16022 = ( n16009 & ~n16020 ) | ( n16009 & n16021 ) | ( ~n16020 & n16021 ) ;
  assign n16023 = ( ~n15678 & n15999 ) | ( ~n15678 & n16022 ) | ( n15999 & n16022 ) ;
  assign n16024 = ( n15678 & n15999 ) | ( n15678 & n16022 ) | ( n15999 & n16022 ) ;
  assign n16025 = ( n15678 & n16023 ) | ( n15678 & ~n16024 ) | ( n16023 & ~n16024 ) ;
  assign n16026 = ( ~n15681 & n15989 ) | ( ~n15681 & n16025 ) | ( n15989 & n16025 ) ;
  assign n16027 = ( n15681 & n15989 ) | ( n15681 & n16025 ) | ( n15989 & n16025 ) ;
  assign n16028 = ( n15681 & n16026 ) | ( n15681 & ~n16027 ) | ( n16026 & ~n16027 ) ;
  assign n16029 = ( ~n15684 & n15979 ) | ( ~n15684 & n16028 ) | ( n15979 & n16028 ) ;
  assign n16030 = ( n15684 & n15979 ) | ( n15684 & n16028 ) | ( n15979 & n16028 ) ;
  assign n16031 = ( n15684 & n16029 ) | ( n15684 & ~n16030 ) | ( n16029 & ~n16030 ) ;
  assign n16032 = ( n15822 & n15969 ) | ( n15822 & n16031 ) | ( n15969 & n16031 ) ;
  assign n16033 = n5914 & ~n13473 ;
  assign n16034 = n6332 & ~n13280 ;
  assign n16035 = n5909 & ~n10235 ;
  assign n16036 = n16034 | n16035 ;
  assign n16037 = n16033 | n16036 ;
  assign n16038 = n5915 | n16037 ;
  assign n16039 = ( ~n13480 & n16037 ) | ( ~n13480 & n16038 ) | ( n16037 & n16038 ) ;
  assign n16040 = x14 & ~n16039 ;
  assign n16041 = ~x14 & n16039 ;
  assign n16042 = n16040 | n16041 ;
  assign n16043 = n5584 & ~n10237 ;
  assign n16044 = x17 & n16043 ;
  assign n16045 = n5413 & ~n10332 ;
  assign n16046 = n5417 | n16045 ;
  assign n16047 = ( n10214 & n16045 ) | ( n10214 & n16046 ) | ( n16045 & n16046 ) ;
  assign n16048 = n5418 | n16047 ;
  assign n16049 = ( n12953 & n16047 ) | ( n12953 & n16048 ) | ( n16047 & n16048 ) ;
  assign n16050 = x17 & ~n16049 ;
  assign n16051 = ( ~x17 & n16043 ) | ( ~x17 & n16049 ) | ( n16043 & n16049 ) ;
  assign n16052 = ( ~n16044 & n16050 ) | ( ~n16044 & n16051 ) | ( n16050 & n16051 ) ;
  assign n16053 = n4879 & n10397 ;
  assign n16054 = x20 & n16053 ;
  assign n16055 = n4874 & n10239 ;
  assign n16056 = n4878 | n16055 ;
  assign n16057 = ( n10329 & n16055 ) | ( n10329 & n16056 ) | ( n16055 & n16056 ) ;
  assign n16058 = n5232 & n10326 ;
  assign n16059 = n16057 | n16058 ;
  assign n16060 = x20 & ~n16059 ;
  assign n16061 = ( ~x20 & n16053 ) | ( ~x20 & n16059 ) | ( n16053 & n16059 ) ;
  assign n16062 = ( ~n16054 & n16060 ) | ( ~n16054 & n16061 ) | ( n16060 & n16061 ) ;
  assign n16063 = n4637 & n10243 ;
  assign n16064 = x23 & n16063 ;
  assign n16065 = n4584 & ~n10320 ;
  assign n16066 = n4649 | n16065 ;
  assign n16067 = ( n10241 & n16065 ) | ( n10241 & n16066 ) | ( n16065 & n16066 ) ;
  assign n16068 = n4591 | n16067 ;
  assign n16069 = ( n12105 & n16067 ) | ( n12105 & n16068 ) | ( n16067 & n16068 ) ;
  assign n16070 = x23 & ~n16069 ;
  assign n16071 = ( ~x23 & n16063 ) | ( ~x23 & n16069 ) | ( n16063 & n16069 ) ;
  assign n16072 = ( ~n16064 & n16070 ) | ( ~n16064 & n16071 ) | ( n16070 & n16071 ) ;
  assign n16073 = n4215 & n10245 ;
  assign n16074 = n4200 & ~n10316 ;
  assign n16075 = n2083 & n10247 ;
  assign n16076 = n16074 | n16075 ;
  assign n16077 = n16073 | n16076 ;
  assign n16078 = x26 & n16077 ;
  assign n16079 = n4203 & ~n11676 ;
  assign n16080 = ( ~x26 & n16077 ) | ( ~x26 & n16079 ) | ( n16077 & n16079 ) ;
  assign n16081 = x26 & ~n16079 ;
  assign n16082 = ( ~n16078 & n16080 ) | ( ~n16078 & n16081 ) | ( n16080 & n16081 ) ;
  assign n16083 = n4039 & n10312 ;
  assign n16084 = x29 & n16083 ;
  assign n16085 = n3501 & ~n10249 ;
  assign n16086 = n3536 & n10251 ;
  assign n16087 = n16085 | n16086 ;
  assign n16088 = n3541 | n16087 ;
  assign n16089 = ( ~n11486 & n16087 ) | ( ~n11486 & n16088 ) | ( n16087 & n16088 ) ;
  assign n16090 = x29 & ~n16089 ;
  assign n16091 = ( ~x29 & n16083 ) | ( ~x29 & n16089 ) | ( n16083 & n16089 ) ;
  assign n16092 = ( ~n16084 & n16090 ) | ( ~n16084 & n16091 ) | ( n16090 & n16091 ) ;
  assign n16093 = n3273 & n10257 ;
  assign n16094 = n3270 | n16093 ;
  assign n16095 = ( ~n10253 & n16093 ) | ( ~n10253 & n16094 ) | ( n16093 & n16094 ) ;
  assign n16096 = n390 | n16095 ;
  assign n16097 = ( ~n11297 & n16095 ) | ( ~n11297 & n16096 ) | ( n16095 & n16096 ) ;
  assign n16098 = n3274 & n10255 ;
  assign n16099 = n16097 | n16098 ;
  assign n16100 = n900 | n10135 ;
  assign n16101 = n3037 | n16100 ;
  assign n16102 = n200 | n350 ;
  assign n16103 = n322 | n16102 ;
  assign n16104 = n2488 | n16103 ;
  assign n16105 = n16101 | n16104 ;
  assign n16106 = n4287 | n16105 ;
  assign n16107 = n284 | n4381 ;
  assign n16108 = n165 | n238 ;
  assign n16109 = n16107 | n16108 ;
  assign n16110 = n164 | n397 ;
  assign n16111 = n661 | n16110 ;
  assign n16112 = n16109 | n16111 ;
  assign n16113 = n14455 | n16112 ;
  assign n16114 = n15359 & ~n16113 ;
  assign n16115 = ~n16106 & n16114 ;
  assign n16116 = ~n5633 & n16115 ;
  assign n16117 = ~n3231 & n16116 ;
  assign n16118 = ( ~n15917 & n16099 ) | ( ~n15917 & n16117 ) | ( n16099 & n16117 ) ;
  assign n16119 = ( n15917 & n16099 ) | ( n15917 & ~n16117 ) | ( n16099 & ~n16117 ) ;
  assign n16120 = ( ~n16099 & n16118 ) | ( ~n16099 & n16119 ) | ( n16118 & n16119 ) ;
  assign n16121 = ( ~n15920 & n16092 ) | ( ~n15920 & n16120 ) | ( n16092 & n16120 ) ;
  assign n16122 = ( n15920 & n16092 ) | ( n15920 & ~n16120 ) | ( n16092 & ~n16120 ) ;
  assign n16123 = ( ~n16092 & n16121 ) | ( ~n16092 & n16122 ) | ( n16121 & n16122 ) ;
  assign n16124 = ( n15922 & n16082 ) | ( n15922 & ~n16123 ) | ( n16082 & ~n16123 ) ;
  assign n16125 = ( ~n15922 & n16082 ) | ( ~n15922 & n16123 ) | ( n16082 & n16123 ) ;
  assign n16126 = ( ~n16082 & n16124 ) | ( ~n16082 & n16125 ) | ( n16124 & n16125 ) ;
  assign n16127 = ( ~n15926 & n16072 ) | ( ~n15926 & n16126 ) | ( n16072 & n16126 ) ;
  assign n16128 = ( n15926 & n16072 ) | ( n15926 & ~n16126 ) | ( n16072 & ~n16126 ) ;
  assign n16129 = ( ~n16072 & n16127 ) | ( ~n16072 & n16128 ) | ( n16127 & n16128 ) ;
  assign n16130 = ( ~n15928 & n16062 ) | ( ~n15928 & n16129 ) | ( n16062 & n16129 ) ;
  assign n16131 = ( n15928 & n16062 ) | ( n15928 & ~n16129 ) | ( n16062 & ~n16129 ) ;
  assign n16132 = ( ~n16062 & n16130 ) | ( ~n16062 & n16131 ) | ( n16130 & n16131 ) ;
  assign n16133 = ( n15931 & n16052 ) | ( n15931 & ~n16132 ) | ( n16052 & ~n16132 ) ;
  assign n16134 = ( ~n15931 & n16052 ) | ( ~n15931 & n16132 ) | ( n16052 & n16132 ) ;
  assign n16135 = ( ~n16052 & n16133 ) | ( ~n16052 & n16134 ) | ( n16133 & n16134 ) ;
  assign n16136 = ( ~n15935 & n16042 ) | ( ~n15935 & n16135 ) | ( n16042 & n16135 ) ;
  assign n16137 = ( n15935 & n16042 ) | ( n15935 & ~n16135 ) | ( n16042 & ~n16135 ) ;
  assign n16138 = ( ~n16042 & n16136 ) | ( ~n16042 & n16137 ) | ( n16136 & n16137 ) ;
  assign n16139 = ( x8 & ~x9 ) | ( x8 & x10 ) | ( ~x9 & x10 ) ;
  assign n16140 = ( x9 & ~x11 ) | ( x9 & n16139 ) | ( ~x11 & n16139 ) ;
  assign n16141 = x11 & ~n6795 ;
  assign n16142 = n13475 | n16141 ;
  assign n16143 = ( n6795 & ~n13475 ) | ( n6795 & n16141 ) | ( ~n13475 & n16141 ) ;
  assign n16144 = ( n16140 & n16142 ) | ( n16140 & n16143 ) | ( n16142 & n16143 ) ;
  assign n16145 = ( n15937 & ~n16138 ) | ( n15937 & n16144 ) | ( ~n16138 & n16144 ) ;
  assign n16146 = ( n15937 & n16138 ) | ( n15937 & n16144 ) | ( n16138 & n16144 ) ;
  assign n16147 = ( n16138 & n16145 ) | ( n16138 & ~n16146 ) | ( n16145 & ~n16146 ) ;
  assign n16148 = ( n15950 & n15952 ) | ( n15950 & ~n16147 ) | ( n15952 & ~n16147 ) ;
  assign n16149 = ( ~n15950 & n15952 ) | ( ~n15950 & n16147 ) | ( n15952 & n16147 ) ;
  assign n16150 = ( ~n15952 & n16148 ) | ( ~n15952 & n16149 ) | ( n16148 & n16149 ) ;
  assign n16151 = n40 & ~n16150 ;
  assign n16152 = n8721 & ~n15954 ;
  assign n16153 = n8340 & ~n15806 ;
  assign n16154 = n16152 | n16153 ;
  assign n16155 = n16151 | n16154 ;
  assign n16156 = x5 & n16155 ;
  assign n16157 = n15954 | n15961 ;
  assign n16158 = n16150 | n16157 ;
  assign n16159 = n15963 | n16150 ;
  assign n16160 = ( n15963 & n16150 ) | ( n15963 & ~n16157 ) | ( n16150 & ~n16157 ) ;
  assign n16161 = ( n16158 & ~n16159 ) | ( n16158 & n16160 ) | ( ~n16159 & n16160 ) ;
  assign n16162 = n8341 & ~n16161 ;
  assign n16163 = ( ~x5 & n16155 ) | ( ~x5 & n16162 ) | ( n16155 & n16162 ) ;
  assign n16164 = x5 & ~n16162 ;
  assign n16165 = ( ~n16156 & n16163 ) | ( ~n16156 & n16164 ) | ( n16163 & n16164 ) ;
  assign n16166 = n7644 & ~n15394 ;
  assign n16167 = x8 & n16166 ;
  assign n16168 = n7341 & ~n15184 ;
  assign n16169 = n7345 | n16168 ;
  assign n16170 = ( n15561 & n16168 ) | ( n15561 & n16169 ) | ( n16168 & n16169 ) ;
  assign n16171 = n7346 | n16170 ;
  assign n16172 = ( n15573 & n16170 ) | ( n15573 & n16171 ) | ( n16170 & n16171 ) ;
  assign n16173 = x8 & ~n16172 ;
  assign n16174 = ( ~x8 & n16166 ) | ( ~x8 & n16172 ) | ( n16166 & n16172 ) ;
  assign n16175 = ( ~n16167 & n16173 ) | ( ~n16167 & n16174 ) | ( n16173 & n16174 ) ;
  assign n16176 = n6332 & n13992 ;
  assign n16177 = x14 & n16176 ;
  assign n16178 = n5909 & n13996 ;
  assign n16179 = n5914 | n16178 ;
  assign n16180 = ( n14352 & n16178 ) | ( n14352 & n16179 ) | ( n16178 & n16179 ) ;
  assign n16181 = n5915 | n16180 ;
  assign n16182 = ( n14363 & n16180 ) | ( n14363 & n16181 ) | ( n16180 & n16181 ) ;
  assign n16183 = x14 & ~n16182 ;
  assign n16184 = ( ~x14 & n16176 ) | ( ~x14 & n16182 ) | ( n16176 & n16182 ) ;
  assign n16185 = ( ~n16177 & n16183 ) | ( ~n16177 & n16184 ) | ( n16183 & n16184 ) ;
  assign n16186 = n5584 & ~n14000 ;
  assign n16187 = x17 & n16186 ;
  assign n16188 = n5413 & ~n14007 ;
  assign n16189 = n5417 | n16188 ;
  assign n16190 = ( n13998 & n16188 ) | ( n13998 & n16189 ) | ( n16188 & n16189 ) ;
  assign n16191 = n5418 | n16190 ;
  assign n16192 = ( n14115 & n16190 ) | ( n14115 & n16191 ) | ( n16190 & n16191 ) ;
  assign n16193 = x17 & ~n16192 ;
  assign n16194 = ( ~x17 & n16186 ) | ( ~x17 & n16192 ) | ( n16186 & n16192 ) ;
  assign n16195 = ( ~n16187 & n16193 ) | ( ~n16187 & n16194 ) | ( n16193 & n16194 ) ;
  assign n16196 = n5232 & ~n14004 ;
  assign n16197 = n4874 & ~n14014 ;
  assign n16198 = n16196 | n16197 ;
  assign n16199 = n4879 | n16198 ;
  assign n16200 = ( n14072 & n16198 ) | ( n14072 & n16199 ) | ( n16198 & n16199 ) ;
  assign n16201 = n4878 & n14002 ;
  assign n16202 = n16200 | n16201 ;
  assign n16203 = ~x20 & n16202 ;
  assign n16204 = x20 & ~n15672 ;
  assign n16205 = ~n16015 & n16204 ;
  assign n16206 = ( x20 & n16202 ) | ( x20 & ~n16205 ) | ( n16202 & ~n16205 ) ;
  assign n16207 = n16202 & ~n16205 ;
  assign n16208 = ( n16203 & n16206 ) | ( n16203 & ~n16207 ) | ( n16206 & ~n16207 ) ;
  assign n16209 = ( ~n16020 & n16195 ) | ( ~n16020 & n16208 ) | ( n16195 & n16208 ) ;
  assign n16210 = ( n16020 & n16195 ) | ( n16020 & n16208 ) | ( n16195 & n16208 ) ;
  assign n16211 = ( n16020 & n16209 ) | ( n16020 & ~n16210 ) | ( n16209 & ~n16210 ) ;
  assign n16212 = ( ~n16024 & n16185 ) | ( ~n16024 & n16211 ) | ( n16185 & n16211 ) ;
  assign n16213 = ( n16024 & n16185 ) | ( n16024 & n16211 ) | ( n16185 & n16211 ) ;
  assign n16214 = ( n16024 & n16212 ) | ( n16024 & ~n16213 ) | ( n16212 & ~n16213 ) ;
  assign n16215 = n6796 & ~n14723 ;
  assign n16216 = x11 & n16215 ;
  assign n16217 = n6567 & n14520 ;
  assign n16218 = n6570 | n16217 ;
  assign n16219 = ( n14942 & n16217 ) | ( n14942 & n16218 ) | ( n16217 & n16218 ) ;
  assign n16220 = n6571 | n16219 ;
  assign n16221 = ( ~n14953 & n16219 ) | ( ~n14953 & n16220 ) | ( n16219 & n16220 ) ;
  assign n16222 = x11 & ~n16221 ;
  assign n16223 = ( ~x11 & n16215 ) | ( ~x11 & n16221 ) | ( n16215 & n16221 ) ;
  assign n16224 = ( ~n16216 & n16222 ) | ( ~n16216 & n16223 ) | ( n16222 & n16223 ) ;
  assign n16225 = ( ~n16027 & n16214 ) | ( ~n16027 & n16224 ) | ( n16214 & n16224 ) ;
  assign n16226 = ( n16027 & n16214 ) | ( n16027 & n16224 ) | ( n16214 & n16224 ) ;
  assign n16227 = ( n16027 & n16225 ) | ( n16027 & ~n16226 ) | ( n16225 & ~n16226 ) ;
  assign n16228 = ( n16030 & n16175 ) | ( n16030 & n16227 ) | ( n16175 & n16227 ) ;
  assign n16229 = ( ~n16030 & n16175 ) | ( ~n16030 & n16227 ) | ( n16175 & n16227 ) ;
  assign n16230 = ( n16030 & ~n16228 ) | ( n16030 & n16229 ) | ( ~n16228 & n16229 ) ;
  assign n16231 = ( n16032 & n16165 ) | ( n16032 & n16230 ) | ( n16165 & n16230 ) ;
  assign n16232 = n5909 & ~n13280 ;
  assign n16233 = n5914 | n16232 ;
  assign n16234 = ( n13475 & n16232 ) | ( n13475 & n16233 ) | ( n16232 & n16233 ) ;
  assign n16235 = n6332 & ~n13473 ;
  assign n16236 = n16234 | n16235 ;
  assign n16237 = x14 & n16236 ;
  assign n16238 = n5915 & n13671 ;
  assign n16239 = ( ~x14 & n16236 ) | ( ~x14 & n16238 ) | ( n16236 & n16238 ) ;
  assign n16240 = x14 & ~n16238 ;
  assign n16241 = ( ~n16237 & n16239 ) | ( ~n16237 & n16240 ) | ( n16239 & n16240 ) ;
  assign n16242 = n5584 & n10214 ;
  assign n16243 = x17 & n16242 ;
  assign n16244 = n5413 & ~n10237 ;
  assign n16245 = n5417 | n16244 ;
  assign n16246 = ( ~n10235 & n16244 ) | ( ~n10235 & n16245 ) | ( n16244 & n16245 ) ;
  assign n16247 = n5418 | n16246 ;
  assign n16248 = ( n10371 & n16246 ) | ( n10371 & n16247 ) | ( n16246 & n16247 ) ;
  assign n16249 = x17 & ~n16248 ;
  assign n16250 = ( ~x17 & n16242 ) | ( ~x17 & n16248 ) | ( n16242 & n16248 ) ;
  assign n16251 = ( ~n16243 & n16249 ) | ( ~n16243 & n16250 ) | ( n16249 & n16250 ) ;
  assign n16252 = n5232 & n10329 ;
  assign n16253 = x20 & n16252 ;
  assign n16254 = n4874 & n10326 ;
  assign n16255 = n4878 | n16254 ;
  assign n16256 = ( ~n10332 & n16254 ) | ( ~n10332 & n16255 ) | ( n16254 & n16255 ) ;
  assign n16257 = n4879 | n16256 ;
  assign n16258 = ( ~n10383 & n16256 ) | ( ~n10383 & n16257 ) | ( n16256 & n16257 ) ;
  assign n16259 = x20 & ~n16258 ;
  assign n16260 = ( ~x20 & n16252 ) | ( ~x20 & n16258 ) | ( n16252 & n16258 ) ;
  assign n16261 = ( ~n16253 & n16259 ) | ( ~n16253 & n16260 ) | ( n16259 & n16260 ) ;
  assign n16262 = n4637 & n10241 ;
  assign n16263 = x23 & n16262 ;
  assign n16264 = n4584 & n10243 ;
  assign n16265 = n4649 | n16264 ;
  assign n16266 = ( n10239 & n16264 ) | ( n10239 & n16265 ) | ( n16264 & n16265 ) ;
  assign n16267 = n4591 | n16266 ;
  assign n16268 = ( n12575 & n16266 ) | ( n12575 & n16267 ) | ( n16266 & n16267 ) ;
  assign n16269 = x23 & ~n16268 ;
  assign n16270 = ( ~x23 & n16262 ) | ( ~x23 & n16268 ) | ( n16262 & n16268 ) ;
  assign n16271 = ( ~n16263 & n16269 ) | ( ~n16263 & n16270 ) | ( n16269 & n16270 ) ;
  assign n16272 = n4215 & ~n10320 ;
  assign n16273 = x26 & n16272 ;
  assign n16274 = n4200 & n10245 ;
  assign n16275 = n2083 & ~n10316 ;
  assign n16276 = n16274 | n16275 ;
  assign n16277 = n4203 | n16276 ;
  assign n16278 = ( ~n10414 & n16276 ) | ( ~n10414 & n16277 ) | ( n16276 & n16277 ) ;
  assign n16279 = x26 & ~n16278 ;
  assign n16280 = ( ~x26 & n16272 ) | ( ~x26 & n16278 ) | ( n16272 & n16278 ) ;
  assign n16281 = ( ~n16273 & n16279 ) | ( ~n16273 & n16280 ) | ( n16279 & n16280 ) ;
  assign n16282 = n3501 & n10312 ;
  assign n16283 = x29 & n16282 ;
  assign n16284 = n3536 & ~n10249 ;
  assign n16285 = n4039 | n16284 ;
  assign n16286 = ( n10247 & n16284 ) | ( n10247 & n16285 ) | ( n16284 & n16285 ) ;
  assign n16287 = n3541 | n16286 ;
  assign n16288 = ( n10428 & n16286 ) | ( n10428 & n16287 ) | ( n16286 & n16287 ) ;
  assign n16289 = x29 & ~n16288 ;
  assign n16290 = ( ~x29 & n16282 ) | ( ~x29 & n16288 ) | ( n16282 & n16288 ) ;
  assign n16291 = ( ~n16283 & n16289 ) | ( ~n16283 & n16290 ) | ( n16289 & n16290 ) ;
  assign n16292 = n48 | n3561 ;
  assign n16293 = n3743 | n16292 ;
  assign n16294 = n736 | n16293 ;
  assign n16295 = n361 | n1379 ;
  assign n16296 = n16294 | n16295 ;
  assign n16297 = n689 | n3206 ;
  assign n16298 = n663 | n14871 ;
  assign n16299 = n16297 | n16298 ;
  assign n16300 = n2128 | n16299 ;
  assign n16301 = n16296 | n16300 ;
  assign n16302 = n13206 | n16301 ;
  assign n16303 = n4518 | n16302 ;
  assign n16304 = n12857 & ~n16303 ;
  assign n16305 = ( n16117 & n16118 ) | ( n16117 & ~n16304 ) | ( n16118 & ~n16304 ) ;
  assign n16306 = ( n16117 & ~n16118 ) | ( n16117 & n16304 ) | ( ~n16118 & n16304 ) ;
  assign n16307 = ( ~n16117 & n16305 ) | ( ~n16117 & n16306 ) | ( n16305 & n16306 ) ;
  assign n16308 = n3273 & n10255 ;
  assign n16309 = n3270 | n16308 ;
  assign n16310 = ( n10251 & n16308 ) | ( n10251 & n16309 ) | ( n16308 & n16309 ) ;
  assign n16311 = n390 | n16310 ;
  assign n16312 = ( ~n11309 & n16310 ) | ( ~n11309 & n16311 ) | ( n16310 & n16311 ) ;
  assign n16313 = n3274 & ~n10253 ;
  assign n16314 = n16312 | n16313 ;
  assign n16315 = ( n16291 & ~n16307 ) | ( n16291 & n16314 ) | ( ~n16307 & n16314 ) ;
  assign n16316 = ( n16291 & n16307 ) | ( n16291 & ~n16314 ) | ( n16307 & ~n16314 ) ;
  assign n16317 = ( ~n16291 & n16315 ) | ( ~n16291 & n16316 ) | ( n16315 & n16316 ) ;
  assign n16318 = ( n16122 & n16281 ) | ( n16122 & ~n16317 ) | ( n16281 & ~n16317 ) ;
  assign n16319 = ( ~n16122 & n16281 ) | ( ~n16122 & n16317 ) | ( n16281 & n16317 ) ;
  assign n16320 = ( ~n16281 & n16318 ) | ( ~n16281 & n16319 ) | ( n16318 & n16319 ) ;
  assign n16321 = ( ~n16124 & n16271 ) | ( ~n16124 & n16320 ) | ( n16271 & n16320 ) ;
  assign n16322 = ( n16124 & n16271 ) | ( n16124 & ~n16320 ) | ( n16271 & ~n16320 ) ;
  assign n16323 = ( ~n16271 & n16321 ) | ( ~n16271 & n16322 ) | ( n16321 & n16322 ) ;
  assign n16324 = ( n16128 & n16261 ) | ( n16128 & ~n16323 ) | ( n16261 & ~n16323 ) ;
  assign n16325 = ( ~n16128 & n16261 ) | ( ~n16128 & n16323 ) | ( n16261 & n16323 ) ;
  assign n16326 = ( ~n16261 & n16324 ) | ( ~n16261 & n16325 ) | ( n16324 & n16325 ) ;
  assign n16327 = ( ~n16131 & n16251 ) | ( ~n16131 & n16326 ) | ( n16251 & n16326 ) ;
  assign n16328 = ( n16131 & n16251 ) | ( n16131 & ~n16326 ) | ( n16251 & ~n16326 ) ;
  assign n16329 = ( ~n16251 & n16327 ) | ( ~n16251 & n16328 ) | ( n16327 & n16328 ) ;
  assign n16330 = ( n16133 & n16241 ) | ( n16133 & ~n16329 ) | ( n16241 & ~n16329 ) ;
  assign n16331 = ( ~n16133 & n16241 ) | ( ~n16133 & n16329 ) | ( n16241 & n16329 ) ;
  assign n16332 = ( ~n16241 & n16330 ) | ( ~n16241 & n16331 ) | ( n16330 & n16331 ) ;
  assign n16333 = ( n16137 & ~n16140 ) | ( n16137 & n16332 ) | ( ~n16140 & n16332 ) ;
  assign n16334 = ( n16137 & n16140 ) | ( n16137 & ~n16332 ) | ( n16140 & ~n16332 ) ;
  assign n16335 = ( ~n16137 & n16333 ) | ( ~n16137 & n16334 ) | ( n16333 & n16334 ) ;
  assign n16336 = ( n16145 & ~n16148 ) | ( n16145 & n16335 ) | ( ~n16148 & n16335 ) ;
  assign n16337 = ( n16145 & n16148 ) | ( n16145 & ~n16335 ) | ( n16148 & ~n16335 ) ;
  assign n16338 = ( ~n16145 & n16336 ) | ( ~n16145 & n16337 ) | ( n16336 & n16337 ) ;
  assign n16339 = n40 & ~n16338 ;
  assign n16340 = n8721 & ~n16150 ;
  assign n16341 = n8340 & ~n15954 ;
  assign n16342 = n16340 | n16341 ;
  assign n16343 = n16339 | n16342 ;
  assign n16344 = x5 & n16343 ;
  assign n16345 = n16150 & n16157 ;
  assign n16346 = n16338 & n16345 ;
  assign n16347 = n16159 & n16338 ;
  assign n16348 = ( n16159 & n16338 ) | ( n16159 & ~n16345 ) | ( n16338 & ~n16345 ) ;
  assign n16349 = ( n16346 & ~n16347 ) | ( n16346 & n16348 ) | ( ~n16347 & n16348 ) ;
  assign n16350 = n8341 & ~n16349 ;
  assign n16351 = ( ~x5 & n16343 ) | ( ~x5 & n16350 ) | ( n16343 & n16350 ) ;
  assign n16352 = x5 & ~n16350 ;
  assign n16353 = ( ~n16344 & n16351 ) | ( ~n16344 & n16352 ) | ( n16351 & n16352 ) ;
  assign n16354 = n7644 & n15561 ;
  assign n16355 = x8 & n16354 ;
  assign n16356 = n7341 & ~n15394 ;
  assign n16357 = n7345 | n16356 ;
  assign n16358 = ( ~n15806 & n16356 ) | ( ~n15806 & n16357 ) | ( n16356 & n16357 ) ;
  assign n16359 = n7346 | n16358 ;
  assign n16360 = ( n15817 & n16358 ) | ( n15817 & n16359 ) | ( n16358 & n16359 ) ;
  assign n16361 = x8 & ~n16360 ;
  assign n16362 = ( ~x8 & n16354 ) | ( ~x8 & n16360 ) | ( n16354 & n16360 ) ;
  assign n16363 = ( ~n16355 & n16361 ) | ( ~n16355 & n16362 ) | ( n16361 & n16362 ) ;
  assign n16364 = n6796 & n14942 ;
  assign n16365 = x11 & n16364 ;
  assign n16366 = n6567 & ~n14723 ;
  assign n16367 = n6570 | n16366 ;
  assign n16368 = ( ~n15184 & n16366 ) | ( ~n15184 & n16367 ) | ( n16366 & n16367 ) ;
  assign n16369 = n6571 | n16368 ;
  assign n16370 = ( ~n15195 & n16368 ) | ( ~n15195 & n16369 ) | ( n16368 & n16369 ) ;
  assign n16371 = x11 & ~n16370 ;
  assign n16372 = ( ~x11 & n16364 ) | ( ~x11 & n16370 ) | ( n16364 & n16370 ) ;
  assign n16373 = ( ~n16365 & n16371 ) | ( ~n16365 & n16372 ) | ( n16371 & n16372 ) ;
  assign n16374 = n6332 & n14352 ;
  assign n16375 = x14 & n16374 ;
  assign n16376 = n5909 & n13992 ;
  assign n16377 = n5914 | n16376 ;
  assign n16378 = ( n14520 & n16376 ) | ( n14520 & n16377 ) | ( n16376 & n16377 ) ;
  assign n16379 = n5915 | n16378 ;
  assign n16380 = ( n14531 & n16378 ) | ( n14531 & n16379 ) | ( n16378 & n16379 ) ;
  assign n16381 = x14 & ~n16380 ;
  assign n16382 = ( ~x14 & n16374 ) | ( ~x14 & n16380 ) | ( n16374 & n16380 ) ;
  assign n16383 = ( ~n16375 & n16381 ) | ( ~n16375 & n16382 ) | ( n16381 & n16382 ) ;
  assign n16384 = n5584 & n13998 ;
  assign n16385 = x17 & n16384 ;
  assign n16386 = n5413 & ~n14000 ;
  assign n16387 = n5417 | n16386 ;
  assign n16388 = ( n13996 & n16386 ) | ( n13996 & n16387 ) | ( n16386 & n16387 ) ;
  assign n16389 = n5418 | n16388 ;
  assign n16390 = ( ~n14130 & n16388 ) | ( ~n14130 & n16389 ) | ( n16388 & n16389 ) ;
  assign n16391 = x17 & ~n16390 ;
  assign n16392 = ( ~x17 & n16384 ) | ( ~x17 & n16390 ) | ( n16384 & n16390 ) ;
  assign n16393 = ( ~n16385 & n16391 ) | ( ~n16385 & n16392 ) | ( n16391 & n16392 ) ;
  assign n16394 = ~n16202 & n16205 ;
  assign n16395 = n5232 & n14002 ;
  assign n16396 = x20 & n16395 ;
  assign n16397 = n4874 & ~n14004 ;
  assign n16398 = n4878 | n16397 ;
  assign n16399 = ( ~n14007 & n16397 ) | ( ~n14007 & n16398 ) | ( n16397 & n16398 ) ;
  assign n16400 = n4879 | n16399 ;
  assign n16401 = ( n14066 & n16399 ) | ( n14066 & n16400 ) | ( n16399 & n16400 ) ;
  assign n16402 = x20 & ~n16401 ;
  assign n16403 = ( ~x20 & n16395 ) | ( ~x20 & n16401 ) | ( n16395 & n16401 ) ;
  assign n16404 = ( ~n16396 & n16402 ) | ( ~n16396 & n16403 ) | ( n16402 & n16403 ) ;
  assign n16405 = n4590 & ~n14014 ;
  assign n16406 = n16394 | n16405 ;
  assign n16407 = n16404 & n16406 ;
  assign n16408 = ( ~n16394 & n16404 ) | ( ~n16394 & n16405 ) | ( n16404 & n16405 ) ;
  assign n16409 = ( n16394 & ~n16407 ) | ( n16394 & n16408 ) | ( ~n16407 & n16408 ) ;
  assign n16410 = ( ~n16210 & n16393 ) | ( ~n16210 & n16409 ) | ( n16393 & n16409 ) ;
  assign n16411 = ( n16210 & n16393 ) | ( n16210 & n16409 ) | ( n16393 & n16409 ) ;
  assign n16412 = ( n16210 & n16410 ) | ( n16210 & ~n16411 ) | ( n16410 & ~n16411 ) ;
  assign n16413 = ( ~n16213 & n16383 ) | ( ~n16213 & n16412 ) | ( n16383 & n16412 ) ;
  assign n16414 = ( n16213 & n16383 ) | ( n16213 & n16412 ) | ( n16383 & n16412 ) ;
  assign n16415 = ( n16213 & n16413 ) | ( n16213 & ~n16414 ) | ( n16413 & ~n16414 ) ;
  assign n16416 = ( ~n16226 & n16373 ) | ( ~n16226 & n16415 ) | ( n16373 & n16415 ) ;
  assign n16417 = ( n16226 & n16373 ) | ( n16226 & n16415 ) | ( n16373 & n16415 ) ;
  assign n16418 = ( n16226 & n16416 ) | ( n16226 & ~n16417 ) | ( n16416 & ~n16417 ) ;
  assign n16419 = ( ~n16228 & n16363 ) | ( ~n16228 & n16418 ) | ( n16363 & n16418 ) ;
  assign n16420 = ( n16228 & n16363 ) | ( n16228 & n16418 ) | ( n16363 & n16418 ) ;
  assign n16421 = ( n16228 & n16419 ) | ( n16228 & ~n16420 ) | ( n16419 & ~n16420 ) ;
  assign n16422 = ( n16231 & n16353 ) | ( n16231 & n16421 ) | ( n16353 & n16421 ) ;
  assign n16423 = ( n5911 & n5914 ) | ( n5911 & n13477 ) | ( n5914 & n13477 ) ;
  assign n16424 = ~x14 & n16423 ;
  assign n16425 = n5909 & ~n13473 ;
  assign n16426 = n6332 | n16425 ;
  assign n16427 = ( n13475 & n16425 ) | ( n13475 & n16426 ) | ( n16425 & n16426 ) ;
  assign n16428 = ( x14 & n16423 ) | ( x14 & n16427 ) | ( n16423 & n16427 ) ;
  assign n16429 = x14 | n16427 ;
  assign n16430 = ( n16424 & ~n16428 ) | ( n16424 & n16429 ) | ( ~n16428 & n16429 ) ;
  assign n16431 = n4879 & n12756 ;
  assign n16432 = x20 & n16431 ;
  assign n16433 = n4878 & ~n10237 ;
  assign n16434 = n5232 & ~n10332 ;
  assign n16435 = n4874 & n10329 ;
  assign n16436 = n16434 | n16435 ;
  assign n16437 = n16433 | n16436 ;
  assign n16438 = x20 & ~n16437 ;
  assign n16439 = ( ~x20 & n16431 ) | ( ~x20 & n16437 ) | ( n16431 & n16437 ) ;
  assign n16440 = ( ~n16432 & n16438 ) | ( ~n16432 & n16439 ) | ( n16438 & n16439 ) ;
  assign n16441 = n4637 & n10239 ;
  assign n16442 = x23 & n16441 ;
  assign n16443 = n4584 & n10241 ;
  assign n16444 = n4649 | n16443 ;
  assign n16445 = ( n10326 & n16443 ) | ( n10326 & n16444 ) | ( n16443 & n16444 ) ;
  assign n16446 = n4591 | n16445 ;
  assign n16447 = ( n12222 & n16445 ) | ( n12222 & n16446 ) | ( n16445 & n16446 ) ;
  assign n16448 = x23 & ~n16447 ;
  assign n16449 = ( ~x23 & n16441 ) | ( ~x23 & n16447 ) | ( n16441 & n16447 ) ;
  assign n16450 = ( ~n16442 & n16448 ) | ( ~n16442 & n16449 ) | ( n16448 & n16449 ) ;
  assign n16451 = n4215 & n10243 ;
  assign n16452 = n4200 & ~n10320 ;
  assign n16453 = n2083 & n10245 ;
  assign n16454 = n16452 | n16453 ;
  assign n16455 = n16451 | n16454 ;
  assign n16456 = x26 & n16455 ;
  assign n16457 = n4203 & ~n11989 ;
  assign n16458 = ( ~x26 & n16455 ) | ( ~x26 & n16457 ) | ( n16455 & n16457 ) ;
  assign n16459 = x26 & ~n16457 ;
  assign n16460 = ( ~n16456 & n16458 ) | ( ~n16456 & n16459 ) | ( n16458 & n16459 ) ;
  assign n16461 = n3541 & ~n11691 ;
  assign n16462 = x29 & n16461 ;
  assign n16463 = n3536 & n10312 ;
  assign n16464 = n4039 | n16463 ;
  assign n16465 = ( ~n10316 & n16463 ) | ( ~n10316 & n16464 ) | ( n16463 & n16464 ) ;
  assign n16466 = n3501 & n10247 ;
  assign n16467 = n16465 | n16466 ;
  assign n16468 = x29 & ~n16467 ;
  assign n16469 = ( ~x29 & n16461 ) | ( ~x29 & n16467 ) | ( n16461 & n16467 ) ;
  assign n16470 = ( ~n16462 & n16468 ) | ( ~n16462 & n16469 ) | ( n16468 & n16469 ) ;
  assign n16471 = n3273 & ~n10253 ;
  assign n16472 = n3270 | n16471 ;
  assign n16473 = ( ~n10249 & n16471 ) | ( ~n10249 & n16472 ) | ( n16471 & n16472 ) ;
  assign n16474 = n390 | n16473 ;
  assign n16475 = ( ~n10441 & n16473 ) | ( ~n10441 & n16474 ) | ( n16473 & n16474 ) ;
  assign n16476 = n3274 & n10251 ;
  assign n16477 = n16475 | n16476 ;
  assign n16478 = n653 & ~n1142 ;
  assign n16479 = ~n5489 & n16478 ;
  assign n16480 = n1777 | n4382 ;
  assign n16481 = n962 | n16480 ;
  assign n16482 = n151 | n734 ;
  assign n16483 = n695 | n16482 ;
  assign n16484 = n16481 | n16483 ;
  assign n16485 = n1586 | n2753 ;
  assign n16486 = n16484 | n16485 ;
  assign n16487 = n1701 | n16486 ;
  assign n16488 = n1756 | n2912 ;
  assign n16489 = n444 | n16488 ;
  assign n16490 = n2647 | n12851 ;
  assign n16491 = n1746 | n16490 ;
  assign n16492 = n16489 | n16491 ;
  assign n16493 = n16487 | n16492 ;
  assign n16494 = n16479 & ~n16493 ;
  assign n16495 = ( ~n16117 & n16140 ) | ( ~n16117 & n16494 ) | ( n16140 & n16494 ) ;
  assign n16496 = ( n16117 & n16140 ) | ( n16117 & n16494 ) | ( n16140 & n16494 ) ;
  assign n16497 = ( n16117 & n16495 ) | ( n16117 & ~n16496 ) | ( n16495 & ~n16496 ) ;
  assign n16498 = ( n16305 & ~n16477 ) | ( n16305 & n16497 ) | ( ~n16477 & n16497 ) ;
  assign n16499 = ( n16305 & n16477 ) | ( n16305 & n16497 ) | ( n16477 & n16497 ) ;
  assign n16500 = ( n16477 & n16498 ) | ( n16477 & ~n16499 ) | ( n16498 & ~n16499 ) ;
  assign n16501 = ( n16315 & n16470 ) | ( n16315 & ~n16500 ) | ( n16470 & ~n16500 ) ;
  assign n16502 = ( n16315 & ~n16470 ) | ( n16315 & n16500 ) | ( ~n16470 & n16500 ) ;
  assign n16503 = ( ~n16315 & n16501 ) | ( ~n16315 & n16502 ) | ( n16501 & n16502 ) ;
  assign n16504 = ( n16318 & n16460 ) | ( n16318 & ~n16503 ) | ( n16460 & ~n16503 ) ;
  assign n16505 = ( n16318 & ~n16460 ) | ( n16318 & n16503 ) | ( ~n16460 & n16503 ) ;
  assign n16506 = ( ~n16318 & n16504 ) | ( ~n16318 & n16505 ) | ( n16504 & n16505 ) ;
  assign n16507 = ( ~n16322 & n16450 ) | ( ~n16322 & n16506 ) | ( n16450 & n16506 ) ;
  assign n16508 = ( n16322 & n16450 ) | ( n16322 & ~n16506 ) | ( n16450 & ~n16506 ) ;
  assign n16509 = ( ~n16450 & n16507 ) | ( ~n16450 & n16508 ) | ( n16507 & n16508 ) ;
  assign n16510 = ( n16324 & ~n16440 ) | ( n16324 & n16509 ) | ( ~n16440 & n16509 ) ;
  assign n16511 = ( n16324 & n16440 ) | ( n16324 & ~n16509 ) | ( n16440 & ~n16509 ) ;
  assign n16512 = ( ~n16324 & n16510 ) | ( ~n16324 & n16511 ) | ( n16510 & n16511 ) ;
  assign n16513 = n5418 & ~n13285 ;
  assign n16514 = x17 & n16513 ;
  assign n16515 = n5413 & n10214 ;
  assign n16516 = n5417 | n16515 ;
  assign n16517 = ( ~n13280 & n16515 ) | ( ~n13280 & n16516 ) | ( n16515 & n16516 ) ;
  assign n16518 = n5584 & ~n10235 ;
  assign n16519 = n16517 | n16518 ;
  assign n16520 = x17 & ~n16519 ;
  assign n16521 = ( ~x17 & n16513 ) | ( ~x17 & n16519 ) | ( n16513 & n16519 ) ;
  assign n16522 = ( ~n16514 & n16520 ) | ( ~n16514 & n16521 ) | ( n16520 & n16521 ) ;
  assign n16523 = ( n16328 & ~n16512 ) | ( n16328 & n16522 ) | ( ~n16512 & n16522 ) ;
  assign n16524 = ( n16328 & n16512 ) | ( n16328 & ~n16522 ) | ( n16512 & ~n16522 ) ;
  assign n16525 = ( ~n16328 & n16523 ) | ( ~n16328 & n16524 ) | ( n16523 & n16524 ) ;
  assign n16526 = ( n16330 & ~n16430 ) | ( n16330 & n16525 ) | ( ~n16430 & n16525 ) ;
  assign n16527 = ( n16330 & n16430 ) | ( n16330 & ~n16525 ) | ( n16430 & ~n16525 ) ;
  assign n16528 = ( ~n16330 & n16526 ) | ( ~n16330 & n16527 ) | ( n16526 & n16527 ) ;
  assign n16529 = ( n16334 & n16337 ) | ( n16334 & ~n16528 ) | ( n16337 & ~n16528 ) ;
  assign n16530 = ( ~n16334 & n16337 ) | ( ~n16334 & n16528 ) | ( n16337 & n16528 ) ;
  assign n16531 = ( ~n16337 & n16529 ) | ( ~n16337 & n16530 ) | ( n16529 & n16530 ) ;
  assign n16532 = n40 & ~n16531 ;
  assign n16533 = n8721 & ~n16338 ;
  assign n16534 = n8340 & ~n16150 ;
  assign n16535 = n16533 | n16534 ;
  assign n16536 = n16532 | n16535 ;
  assign n16537 = x5 & n16536 ;
  assign n16538 = n16338 | n16345 ;
  assign n16539 = n16531 | n16538 ;
  assign n16540 = n16347 | n16531 ;
  assign n16541 = ( n16347 & n16531 ) | ( n16347 & ~n16538 ) | ( n16531 & ~n16538 ) ;
  assign n16542 = ( n16539 & ~n16540 ) | ( n16539 & n16541 ) | ( ~n16540 & n16541 ) ;
  assign n16543 = n8341 & ~n16542 ;
  assign n16544 = ( ~x5 & n16536 ) | ( ~x5 & n16543 ) | ( n16536 & n16543 ) ;
  assign n16545 = x5 & ~n16543 ;
  assign n16546 = ( ~n16537 & n16544 ) | ( ~n16537 & n16545 ) | ( n16544 & n16545 ) ;
  assign n16547 = n7644 & ~n15806 ;
  assign n16548 = x8 & n16547 ;
  assign n16549 = n7341 & n15561 ;
  assign n16550 = n7345 | n16549 ;
  assign n16551 = ( ~n15954 & n16549 ) | ( ~n15954 & n16550 ) | ( n16549 & n16550 ) ;
  assign n16552 = n7346 | n16551 ;
  assign n16553 = ( ~n15965 & n16551 ) | ( ~n15965 & n16552 ) | ( n16551 & n16552 ) ;
  assign n16554 = x8 & ~n16553 ;
  assign n16555 = ( ~x8 & n16547 ) | ( ~x8 & n16553 ) | ( n16547 & n16553 ) ;
  assign n16556 = ( ~n16548 & n16554 ) | ( ~n16548 & n16555 ) | ( n16554 & n16555 ) ;
  assign n16557 = n6796 & ~n15184 ;
  assign n16558 = x11 & n16557 ;
  assign n16559 = n6567 & n14942 ;
  assign n16560 = n6570 | n16559 ;
  assign n16561 = ( ~n15394 & n16559 ) | ( ~n15394 & n16560 ) | ( n16559 & n16560 ) ;
  assign n16562 = n6571 | n16561 ;
  assign n16563 = ( n15405 & n16561 ) | ( n15405 & n16562 ) | ( n16561 & n16562 ) ;
  assign n16564 = x11 & ~n16563 ;
  assign n16565 = ( ~x11 & n16557 ) | ( ~x11 & n16563 ) | ( n16557 & n16563 ) ;
  assign n16566 = ( ~n16558 & n16564 ) | ( ~n16558 & n16565 ) | ( n16564 & n16565 ) ;
  assign n16567 = n5915 & ~n14734 ;
  assign n16568 = x14 & n16567 ;
  assign n16569 = n5909 & n14352 ;
  assign n16570 = n5914 | n16569 ;
  assign n16571 = ( ~n14723 & n16569 ) | ( ~n14723 & n16570 ) | ( n16569 & n16570 ) ;
  assign n16572 = n6332 & n14520 ;
  assign n16573 = n16571 | n16572 ;
  assign n16574 = x14 & ~n16573 ;
  assign n16575 = ( ~x14 & n16567 ) | ( ~x14 & n16573 ) | ( n16567 & n16573 ) ;
  assign n16576 = ( ~n16568 & n16574 ) | ( ~n16568 & n16575 ) | ( n16574 & n16575 ) ;
  assign n16577 = n5417 & n13992 ;
  assign n16578 = n5584 & n13996 ;
  assign n16579 = n5413 & n13998 ;
  assign n16580 = n16578 | n16579 ;
  assign n16581 = n16577 | n16580 ;
  assign n16582 = x17 & n16581 ;
  assign n16583 = n5418 & n14024 ;
  assign n16584 = x17 & ~n16583 ;
  assign n16585 = ( ~x17 & n16581 ) | ( ~x17 & n16583 ) | ( n16581 & n16583 ) ;
  assign n16586 = ( ~n16582 & n16584 ) | ( ~n16582 & n16585 ) | ( n16584 & n16585 ) ;
  assign n16587 = n5232 & ~n14007 ;
  assign n16588 = x20 & n16587 ;
  assign n16589 = n4874 & n14002 ;
  assign n16590 = n4878 | n16589 ;
  assign n16591 = ( ~n14000 & n16589 ) | ( ~n14000 & n16590 ) | ( n16589 & n16590 ) ;
  assign n16592 = n4879 | n16591 ;
  assign n16593 = ( ~n14042 & n16591 ) | ( ~n14042 & n16592 ) | ( n16591 & n16592 ) ;
  assign n16594 = x20 & ~n16593 ;
  assign n16595 = ( ~x20 & n16587 ) | ( ~x20 & n16593 ) | ( n16587 & n16593 ) ;
  assign n16596 = ( ~n16588 & n16594 ) | ( ~n16588 & n16595 ) | ( n16594 & n16595 ) ;
  assign n16597 = n4591 & n14004 ;
  assign n16598 = n4637 & ~n14014 ;
  assign n16599 = ( ~n14014 & n16597 ) | ( ~n14014 & n16598 ) | ( n16597 & n16598 ) ;
  assign n16600 = ( n4590 & n4649 ) | ( n4590 & n14014 ) | ( n4649 & n14014 ) ;
  assign n16601 = ~n14004 & n16600 ;
  assign n16602 = n16599 | n16601 ;
  assign n16603 = n16405 | n16602 ;
  assign n16604 = ( x23 & n16405 ) | ( x23 & ~n16602 ) | ( n16405 & ~n16602 ) ;
  assign n16605 = x23 & ~n16602 ;
  assign n16606 = ( n16603 & ~n16604 ) | ( n16603 & n16605 ) | ( ~n16604 & n16605 ) ;
  assign n16607 = ( n16407 & n16596 ) | ( n16407 & n16606 ) | ( n16596 & n16606 ) ;
  assign n16608 = ( n16407 & ~n16596 ) | ( n16407 & n16606 ) | ( ~n16596 & n16606 ) ;
  assign n16609 = ( n16596 & ~n16607 ) | ( n16596 & n16608 ) | ( ~n16607 & n16608 ) ;
  assign n16610 = ( ~n16411 & n16586 ) | ( ~n16411 & n16609 ) | ( n16586 & n16609 ) ;
  assign n16611 = ( n16411 & n16586 ) | ( n16411 & n16609 ) | ( n16586 & n16609 ) ;
  assign n16612 = ( n16411 & n16610 ) | ( n16411 & ~n16611 ) | ( n16610 & ~n16611 ) ;
  assign n16613 = ( ~n16414 & n16576 ) | ( ~n16414 & n16612 ) | ( n16576 & n16612 ) ;
  assign n16614 = ( n16414 & n16576 ) | ( n16414 & n16612 ) | ( n16576 & n16612 ) ;
  assign n16615 = ( n16414 & n16613 ) | ( n16414 & ~n16614 ) | ( n16613 & ~n16614 ) ;
  assign n16616 = ( n16417 & n16566 ) | ( n16417 & n16615 ) | ( n16566 & n16615 ) ;
  assign n16617 = ( ~n16417 & n16566 ) | ( ~n16417 & n16615 ) | ( n16566 & n16615 ) ;
  assign n16618 = ( n16417 & ~n16616 ) | ( n16417 & n16617 ) | ( ~n16616 & n16617 ) ;
  assign n16619 = ( ~n16420 & n16556 ) | ( ~n16420 & n16618 ) | ( n16556 & n16618 ) ;
  assign n16620 = ( n16420 & n16556 ) | ( n16420 & n16618 ) | ( n16556 & n16618 ) ;
  assign n16621 = ( n16420 & n16619 ) | ( n16420 & ~n16620 ) | ( n16619 & ~n16620 ) ;
  assign n16622 = ( n16422 & n16546 ) | ( n16422 & n16621 ) | ( n16546 & n16621 ) ;
  assign n16623 = ( x11 & ~x12 ) | ( x11 & x13 ) | ( ~x12 & x13 ) ;
  assign n16624 = ( x12 & ~x14 ) | ( x12 & n16623 ) | ( ~x14 & n16623 ) ;
  assign n16625 = ~n5908 & n16624 ;
  assign n16626 = ( n13475 & n16624 ) | ( n13475 & n16625 ) | ( n16624 & n16625 ) ;
  assign n16627 = n5905 & ~n13475 ;
  assign n16628 = n16626 | n16627 ;
  assign n16629 = n5417 & ~n13473 ;
  assign n16630 = n5413 & ~n10235 ;
  assign n16631 = n16629 | n16630 ;
  assign n16632 = n5584 & ~n13280 ;
  assign n16633 = n16631 | n16632 ;
  assign n16634 = n5418 | n16633 ;
  assign n16635 = ( ~n13480 & n16633 ) | ( ~n13480 & n16634 ) | ( n16633 & n16634 ) ;
  assign n16636 = x17 & ~n16635 ;
  assign n16637 = ~x17 & n16635 ;
  assign n16638 = n16636 | n16637 ;
  assign n16639 = n5232 & ~n10237 ;
  assign n16640 = x20 & n16639 ;
  assign n16641 = n4874 & ~n10332 ;
  assign n16642 = n4878 | n16641 ;
  assign n16643 = ( n10214 & n16641 ) | ( n10214 & n16642 ) | ( n16641 & n16642 ) ;
  assign n16644 = n4879 | n16643 ;
  assign n16645 = ( n12953 & n16643 ) | ( n12953 & n16644 ) | ( n16643 & n16644 ) ;
  assign n16646 = x20 & ~n16645 ;
  assign n16647 = ( ~x20 & n16639 ) | ( ~x20 & n16645 ) | ( n16639 & n16645 ) ;
  assign n16648 = ( ~n16640 & n16646 ) | ( ~n16640 & n16647 ) | ( n16646 & n16647 ) ;
  assign n16649 = n4649 & n10329 ;
  assign n16650 = n4591 | n16649 ;
  assign n16651 = ( n10397 & n16649 ) | ( n10397 & n16650 ) | ( n16649 & n16650 ) ;
  assign n16652 = n4584 & n10239 ;
  assign n16653 = ( ~x23 & n16651 ) | ( ~x23 & n16652 ) | ( n16651 & n16652 ) ;
  assign n16654 = n4637 & n10326 ;
  assign n16655 = x23 & ~n16652 ;
  assign n16656 = n16654 | n16655 ;
  assign n16657 = ( n16651 & n16654 ) | ( n16651 & n16655 ) | ( n16654 & n16655 ) ;
  assign n16658 = ( n16653 & n16656 ) | ( n16653 & ~n16657 ) | ( n16656 & ~n16657 ) ;
  assign n16659 = n4215 & n10241 ;
  assign n16660 = n4200 & n10243 ;
  assign n16661 = n2083 & ~n10320 ;
  assign n16662 = n16660 | n16661 ;
  assign n16663 = n16659 | n16662 ;
  assign n16664 = x26 & n16663 ;
  assign n16665 = n4203 & n12105 ;
  assign n16666 = ( ~x26 & n16663 ) | ( ~x26 & n16665 ) | ( n16663 & n16665 ) ;
  assign n16667 = x26 & ~n16665 ;
  assign n16668 = ( ~n16664 & n16666 ) | ( ~n16664 & n16667 ) | ( n16666 & n16667 ) ;
  assign n16669 = n3501 & ~n10316 ;
  assign n16670 = x29 & n16669 ;
  assign n16671 = n3536 & n10247 ;
  assign n16672 = n4039 | n16671 ;
  assign n16673 = ( n10245 & n16671 ) | ( n10245 & n16672 ) | ( n16671 & n16672 ) ;
  assign n16674 = n3541 | n16673 ;
  assign n16675 = ( ~n11676 & n16673 ) | ( ~n11676 & n16674 ) | ( n16673 & n16674 ) ;
  assign n16676 = x29 & ~n16675 ;
  assign n16677 = ( ~x29 & n16669 ) | ( ~x29 & n16675 ) | ( n16669 & n16675 ) ;
  assign n16678 = ( ~n16670 & n16676 ) | ( ~n16670 & n16677 ) | ( n16676 & n16677 ) ;
  assign n16679 = ( n16305 & n16477 ) | ( n16305 & ~n16497 ) | ( n16477 & ~n16497 ) ;
  assign n16680 = n3274 & ~n10249 ;
  assign n16681 = n3273 & n10251 ;
  assign n16682 = n16680 | n16681 ;
  assign n16683 = n390 | n16682 ;
  assign n16684 = ( ~n11486 & n16682 ) | ( ~n11486 & n16683 ) | ( n16682 & n16683 ) ;
  assign n16685 = n3270 & n10312 ;
  assign n16686 = n16684 | n16685 ;
  assign n16687 = n1804 | n4980 ;
  assign n16688 = n662 | n3453 ;
  assign n16689 = n174 | n567 ;
  assign n16690 = n16688 | n16689 ;
  assign n16691 = n477 | n756 ;
  assign n16692 = n3055 | n16691 ;
  assign n16693 = n16690 | n16692 ;
  assign n16694 = n3006 | n16693 ;
  assign n16695 = n443 | n3355 ;
  assign n16696 = n3347 | n16695 ;
  assign n16697 = n1788 | n16696 ;
  assign n16698 = n16694 | n16697 ;
  assign n16699 = n994 | n16698 ;
  assign n16700 = n16687 | n16699 ;
  assign n16701 = ( n16496 & ~n16686 ) | ( n16496 & n16700 ) | ( ~n16686 & n16700 ) ;
  assign n16702 = ( n16496 & n16686 ) | ( n16496 & n16700 ) | ( n16686 & n16700 ) ;
  assign n16703 = ( n16686 & n16701 ) | ( n16686 & ~n16702 ) | ( n16701 & ~n16702 ) ;
  assign n16704 = ( ~n16678 & n16679 ) | ( ~n16678 & n16703 ) | ( n16679 & n16703 ) ;
  assign n16705 = ( n16678 & n16679 ) | ( n16678 & n16703 ) | ( n16679 & n16703 ) ;
  assign n16706 = ( n16678 & n16704 ) | ( n16678 & ~n16705 ) | ( n16704 & ~n16705 ) ;
  assign n16707 = ( n16501 & n16668 ) | ( n16501 & n16706 ) | ( n16668 & n16706 ) ;
  assign n16708 = ( n16501 & ~n16668 ) | ( n16501 & n16706 ) | ( ~n16668 & n16706 ) ;
  assign n16709 = ( n16668 & ~n16707 ) | ( n16668 & n16708 ) | ( ~n16707 & n16708 ) ;
  assign n16710 = ( ~n16504 & n16658 ) | ( ~n16504 & n16709 ) | ( n16658 & n16709 ) ;
  assign n16711 = ( n16504 & n16658 ) | ( n16504 & n16709 ) | ( n16658 & n16709 ) ;
  assign n16712 = ( n16504 & n16710 ) | ( n16504 & ~n16711 ) | ( n16710 & ~n16711 ) ;
  assign n16713 = ( n16508 & ~n16648 ) | ( n16508 & n16712 ) | ( ~n16648 & n16712 ) ;
  assign n16714 = ( n16508 & n16648 ) | ( n16508 & n16712 ) | ( n16648 & n16712 ) ;
  assign n16715 = ( n16648 & n16713 ) | ( n16648 & ~n16714 ) | ( n16713 & ~n16714 ) ;
  assign n16716 = ( ~n16511 & n16638 ) | ( ~n16511 & n16715 ) | ( n16638 & n16715 ) ;
  assign n16717 = ( n16511 & n16638 ) | ( n16511 & n16715 ) | ( n16638 & n16715 ) ;
  assign n16718 = ( n16511 & n16716 ) | ( n16511 & ~n16717 ) | ( n16716 & ~n16717 ) ;
  assign n16719 = ( ~n16523 & n16628 ) | ( ~n16523 & n16718 ) | ( n16628 & n16718 ) ;
  assign n16720 = ( n16523 & n16628 ) | ( n16523 & n16718 ) | ( n16628 & n16718 ) ;
  assign n16721 = ( n16523 & n16719 ) | ( n16523 & ~n16720 ) | ( n16719 & ~n16720 ) ;
  assign n16722 = ( ~n16527 & n16529 ) | ( ~n16527 & n16721 ) | ( n16529 & n16721 ) ;
  assign n16723 = ( n16527 & n16529 ) | ( n16527 & n16721 ) | ( n16529 & n16721 ) ;
  assign n16724 = ( n16527 & n16722 ) | ( n16527 & ~n16723 ) | ( n16722 & ~n16723 ) ;
  assign n16725 = n40 & n16724 ;
  assign n16726 = n8721 & ~n16531 ;
  assign n16727 = n8340 & ~n16338 ;
  assign n16728 = n16726 | n16727 ;
  assign n16729 = n16725 | n16728 ;
  assign n16730 = x5 & n16729 ;
  assign n16731 = ~n16540 & n16724 ;
  assign n16732 = n16531 & n16538 ;
  assign n16733 = ( n16540 & n16724 ) | ( n16540 & ~n16732 ) | ( n16724 & ~n16732 ) ;
  assign n16734 = n16724 & ~n16732 ;
  assign n16735 = ( n16731 & n16733 ) | ( n16731 & ~n16734 ) | ( n16733 & ~n16734 ) ;
  assign n16736 = n8341 & n16735 ;
  assign n16737 = ( ~x5 & n16729 ) | ( ~x5 & n16736 ) | ( n16729 & n16736 ) ;
  assign n16738 = x5 & ~n16736 ;
  assign n16739 = ( ~n16730 & n16737 ) | ( ~n16730 & n16738 ) | ( n16737 & n16738 ) ;
  assign n16740 = n7346 & ~n16161 ;
  assign n16741 = x8 & n16740 ;
  assign n16742 = n7341 & ~n15806 ;
  assign n16743 = n7345 | n16742 ;
  assign n16744 = ( ~n16150 & n16742 ) | ( ~n16150 & n16743 ) | ( n16742 & n16743 ) ;
  assign n16745 = n7644 & ~n15954 ;
  assign n16746 = n16744 | n16745 ;
  assign n16747 = x8 & ~n16746 ;
  assign n16748 = ( ~x8 & n16740 ) | ( ~x8 & n16746 ) | ( n16740 & n16746 ) ;
  assign n16749 = ( ~n16741 & n16747 ) | ( ~n16741 & n16748 ) | ( n16747 & n16748 ) ;
  assign n16750 = n6796 & ~n15394 ;
  assign n16751 = x11 & n16750 ;
  assign n16752 = n6567 & ~n15184 ;
  assign n16753 = n6570 | n16752 ;
  assign n16754 = ( n15561 & n16752 ) | ( n15561 & n16753 ) | ( n16752 & n16753 ) ;
  assign n16755 = n6571 | n16754 ;
  assign n16756 = ( n15573 & n16754 ) | ( n15573 & n16755 ) | ( n16754 & n16755 ) ;
  assign n16757 = x11 & ~n16756 ;
  assign n16758 = ( ~x11 & n16750 ) | ( ~x11 & n16756 ) | ( n16750 & n16756 ) ;
  assign n16759 = ( ~n16751 & n16757 ) | ( ~n16751 & n16758 ) | ( n16757 & n16758 ) ;
  assign n16760 = n5584 & n13992 ;
  assign n16761 = x17 & n16760 ;
  assign n16762 = n5413 & n13996 ;
  assign n16763 = n5417 | n16762 ;
  assign n16764 = ( n14352 & n16762 ) | ( n14352 & n16763 ) | ( n16762 & n16763 ) ;
  assign n16765 = n5418 | n16764 ;
  assign n16766 = ( n14363 & n16764 ) | ( n14363 & n16765 ) | ( n16764 & n16765 ) ;
  assign n16767 = x17 & ~n16766 ;
  assign n16768 = ( ~x17 & n16760 ) | ( ~x17 & n16766 ) | ( n16760 & n16766 ) ;
  assign n16769 = ( ~n16761 & n16767 ) | ( ~n16761 & n16768 ) | ( n16767 & n16768 ) ;
  assign n16770 = n5232 & ~n14000 ;
  assign n16771 = x20 & n16770 ;
  assign n16772 = n4874 & ~n14007 ;
  assign n16773 = n4878 | n16772 ;
  assign n16774 = ( n13998 & n16772 ) | ( n13998 & n16773 ) | ( n16772 & n16773 ) ;
  assign n16775 = n4879 | n16774 ;
  assign n16776 = ( n14115 & n16774 ) | ( n14115 & n16775 ) | ( n16774 & n16775 ) ;
  assign n16777 = x20 & ~n16776 ;
  assign n16778 = ( ~x20 & n16770 ) | ( ~x20 & n16776 ) | ( n16770 & n16776 ) ;
  assign n16779 = ( ~n16771 & n16777 ) | ( ~n16771 & n16778 ) | ( n16777 & n16778 ) ;
  assign n16780 = x23 & n16603 ;
  assign n16781 = n4637 & ~n14004 ;
  assign n16782 = n4584 & ~n14014 ;
  assign n16783 = n16781 | n16782 ;
  assign n16784 = n4591 | n16783 ;
  assign n16785 = ( n14072 & n16783 ) | ( n14072 & n16784 ) | ( n16783 & n16784 ) ;
  assign n16786 = n4649 & n14002 ;
  assign n16787 = n16785 | n16786 ;
  assign n16788 = n16780 & ~n16787 ;
  assign n16789 = ~n16780 & n16787 ;
  assign n16790 = n16788 | n16789 ;
  assign n16791 = ( ~n16607 & n16779 ) | ( ~n16607 & n16790 ) | ( n16779 & n16790 ) ;
  assign n16792 = ( n16607 & n16779 ) | ( n16607 & n16790 ) | ( n16779 & n16790 ) ;
  assign n16793 = ( n16607 & n16791 ) | ( n16607 & ~n16792 ) | ( n16791 & ~n16792 ) ;
  assign n16794 = ( ~n16611 & n16769 ) | ( ~n16611 & n16793 ) | ( n16769 & n16793 ) ;
  assign n16795 = ( n16611 & n16769 ) | ( n16611 & n16793 ) | ( n16769 & n16793 ) ;
  assign n16796 = ( n16611 & n16794 ) | ( n16611 & ~n16795 ) | ( n16794 & ~n16795 ) ;
  assign n16797 = n6332 & ~n14723 ;
  assign n16798 = x14 & n16797 ;
  assign n16799 = n5909 & n14520 ;
  assign n16800 = n5914 | n16799 ;
  assign n16801 = ( n14942 & n16799 ) | ( n14942 & n16800 ) | ( n16799 & n16800 ) ;
  assign n16802 = n5915 | n16801 ;
  assign n16803 = ( ~n14953 & n16801 ) | ( ~n14953 & n16802 ) | ( n16801 & n16802 ) ;
  assign n16804 = x14 & ~n16803 ;
  assign n16805 = ( ~x14 & n16797 ) | ( ~x14 & n16803 ) | ( n16797 & n16803 ) ;
  assign n16806 = ( ~n16798 & n16804 ) | ( ~n16798 & n16805 ) | ( n16804 & n16805 ) ;
  assign n16807 = ( ~n16614 & n16796 ) | ( ~n16614 & n16806 ) | ( n16796 & n16806 ) ;
  assign n16808 = ( n16614 & n16796 ) | ( n16614 & n16806 ) | ( n16796 & n16806 ) ;
  assign n16809 = ( n16614 & n16807 ) | ( n16614 & ~n16808 ) | ( n16807 & ~n16808 ) ;
  assign n16810 = ( ~n16616 & n16759 ) | ( ~n16616 & n16809 ) | ( n16759 & n16809 ) ;
  assign n16811 = ( n16616 & n16759 ) | ( n16616 & n16809 ) | ( n16759 & n16809 ) ;
  assign n16812 = ( n16616 & n16810 ) | ( n16616 & ~n16811 ) | ( n16810 & ~n16811 ) ;
  assign n16813 = ( ~n16620 & n16749 ) | ( ~n16620 & n16812 ) | ( n16749 & n16812 ) ;
  assign n16814 = ( n16620 & n16749 ) | ( n16620 & n16812 ) | ( n16749 & n16812 ) ;
  assign n16815 = ( n16620 & n16813 ) | ( n16620 & ~n16814 ) | ( n16813 & ~n16814 ) ;
  assign n16816 = ( n16622 & n16739 ) | ( n16622 & n16815 ) | ( n16739 & n16815 ) ;
  assign n16817 = n5413 & ~n13280 ;
  assign n16818 = n5417 | n16817 ;
  assign n16819 = ( n13475 & n16817 ) | ( n13475 & n16818 ) | ( n16817 & n16818 ) ;
  assign n16820 = n5584 & ~n13473 ;
  assign n16821 = n16819 | n16820 ;
  assign n16822 = x17 & n16821 ;
  assign n16823 = n5418 & n13671 ;
  assign n16824 = ( ~x17 & n16821 ) | ( ~x17 & n16823 ) | ( n16821 & n16823 ) ;
  assign n16825 = x17 & ~n16823 ;
  assign n16826 = ( ~n16822 & n16824 ) | ( ~n16822 & n16825 ) | ( n16824 & n16825 ) ;
  assign n16827 = n4874 & ~n10237 ;
  assign n16828 = n4878 | n16827 ;
  assign n16829 = ( ~n10235 & n16827 ) | ( ~n10235 & n16828 ) | ( n16827 & n16828 ) ;
  assign n16830 = n5232 & n10214 ;
  assign n16831 = n16829 | n16830 ;
  assign n16832 = x20 & n16831 ;
  assign n16833 = n4879 & n10371 ;
  assign n16834 = x20 & ~n16833 ;
  assign n16835 = ( ~x20 & n16831 ) | ( ~x20 & n16833 ) | ( n16831 & n16833 ) ;
  assign n16836 = ( ~n16832 & n16834 ) | ( ~n16832 & n16835 ) | ( n16834 & n16835 ) ;
  assign n16837 = n4637 & n10329 ;
  assign n16838 = x23 & n16837 ;
  assign n16839 = n4584 & n10326 ;
  assign n16840 = n4649 | n16839 ;
  assign n16841 = ( ~n10332 & n16839 ) | ( ~n10332 & n16840 ) | ( n16839 & n16840 ) ;
  assign n16842 = n4591 | n16841 ;
  assign n16843 = ( ~n10383 & n16841 ) | ( ~n10383 & n16842 ) | ( n16841 & n16842 ) ;
  assign n16844 = x23 & ~n16843 ;
  assign n16845 = ( ~x23 & n16837 ) | ( ~x23 & n16843 ) | ( n16837 & n16843 ) ;
  assign n16846 = ( ~n16838 & n16844 ) | ( ~n16838 & n16845 ) | ( n16844 & n16845 ) ;
  assign n16847 = n4203 & n12575 ;
  assign n16848 = n4215 & n10239 ;
  assign n16849 = n4200 & n10241 ;
  assign n16850 = n2083 & n10243 ;
  assign n16851 = n16849 | n16850 ;
  assign n16852 = n16848 | n16851 ;
  assign n16853 = n16847 | n16852 ;
  assign n16854 = n3501 & n10245 ;
  assign n16855 = n3536 & ~n10316 ;
  assign n16856 = n16854 | n16855 ;
  assign n16857 = n3541 | n16856 ;
  assign n16858 = ( ~n10414 & n16856 ) | ( ~n10414 & n16857 ) | ( n16856 & n16857 ) ;
  assign n16859 = n4039 & ~n10320 ;
  assign n16860 = n16858 | n16859 ;
  assign n16861 = n6269 & ~n16860 ;
  assign n16862 = ~n6269 & n16860 ;
  assign n16863 = n16861 | n16862 ;
  assign n16864 = n3273 & ~n10249 ;
  assign n16865 = n3270 | n16864 ;
  assign n16866 = ( n10247 & n16864 ) | ( n10247 & n16865 ) | ( n16864 & n16865 ) ;
  assign n16867 = n390 | n16866 ;
  assign n16868 = ( n10428 & n16866 ) | ( n10428 & n16867 ) | ( n16866 & n16867 ) ;
  assign n16869 = n3274 & n10312 ;
  assign n16870 = n16868 | n16869 ;
  assign n16871 = n2803 | n3747 ;
  assign n16872 = n372 | n3384 ;
  assign n16873 = n1365 | n2917 ;
  assign n16874 = n16872 | n16873 ;
  assign n16875 = n153 | n644 ;
  assign n16876 = n134 | n321 ;
  assign n16877 = n16875 | n16876 ;
  assign n16878 = n16874 | n16877 ;
  assign n16879 = n16871 | n16878 ;
  assign n16880 = n1309 | n4904 ;
  assign n16881 = n13610 | n16880 ;
  assign n16882 = n16879 | n16881 ;
  assign n16883 = n2600 | n13583 ;
  assign n16884 = n16882 | n16883 ;
  assign n16885 = n900 | n947 ;
  assign n16886 = n1074 | n1560 ;
  assign n16887 = n16885 | n16886 ;
  assign n16888 = n524 | n594 ;
  assign n16889 = n2883 | n16888 ;
  assign n16890 = n16887 | n16889 ;
  assign n16891 = n167 | n5076 ;
  assign n16892 = n3280 | n16891 ;
  assign n16893 = n16890 | n16892 ;
  assign n16894 = n616 | n676 ;
  assign n16895 = n103 | n179 ;
  assign n16896 = n16894 | n16895 ;
  assign n16897 = n659 | n16896 ;
  assign n16898 = n474 | n16897 ;
  assign n16899 = n16295 | n16898 ;
  assign n16900 = n16893 | n16899 ;
  assign n16901 = n16884 | n16900 ;
  assign n16902 = ( ~n16700 & n16870 ) | ( ~n16700 & n16901 ) | ( n16870 & n16901 ) ;
  assign n16903 = ( n16700 & n16870 ) | ( n16700 & n16901 ) | ( n16870 & n16901 ) ;
  assign n16904 = ( n16700 & n16902 ) | ( n16700 & ~n16903 ) | ( n16902 & ~n16903 ) ;
  assign n16905 = ( n16701 & n16705 ) | ( n16701 & n16904 ) | ( n16705 & n16904 ) ;
  assign n16906 = ( n16701 & ~n16705 ) | ( n16701 & n16904 ) | ( ~n16705 & n16904 ) ;
  assign n16907 = ( n16705 & ~n16905 ) | ( n16705 & n16906 ) | ( ~n16905 & n16906 ) ;
  assign n16908 = ( n16853 & n16863 ) | ( n16853 & ~n16907 ) | ( n16863 & ~n16907 ) ;
  assign n16909 = ( n16853 & ~n16863 ) | ( n16853 & n16907 ) | ( ~n16863 & n16907 ) ;
  assign n16910 = ( ~n16853 & n16908 ) | ( ~n16853 & n16909 ) | ( n16908 & n16909 ) ;
  assign n16911 = ( ~n16707 & n16846 ) | ( ~n16707 & n16910 ) | ( n16846 & n16910 ) ;
  assign n16912 = ( n16707 & n16846 ) | ( n16707 & n16910 ) | ( n16846 & n16910 ) ;
  assign n16913 = ( n16707 & n16911 ) | ( n16707 & ~n16912 ) | ( n16911 & ~n16912 ) ;
  assign n16914 = ( n16711 & n16836 ) | ( n16711 & n16913 ) | ( n16836 & n16913 ) ;
  assign n16915 = ( n16711 & ~n16836 ) | ( n16711 & n16913 ) | ( ~n16836 & n16913 ) ;
  assign n16916 = ( n16836 & ~n16914 ) | ( n16836 & n16915 ) | ( ~n16914 & n16915 ) ;
  assign n16917 = ( ~n16714 & n16826 ) | ( ~n16714 & n16916 ) | ( n16826 & n16916 ) ;
  assign n16918 = ( n16714 & n16826 ) | ( n16714 & n16916 ) | ( n16826 & n16916 ) ;
  assign n16919 = ( n16714 & n16917 ) | ( n16714 & ~n16918 ) | ( n16917 & ~n16918 ) ;
  assign n16920 = ( ~n16624 & n16717 ) | ( ~n16624 & n16919 ) | ( n16717 & n16919 ) ;
  assign n16921 = ( n16624 & n16717 ) | ( n16624 & n16919 ) | ( n16717 & n16919 ) ;
  assign n16922 = ( n16624 & n16920 ) | ( n16624 & ~n16921 ) | ( n16920 & ~n16921 ) ;
  assign n16923 = ( ~n16720 & n16723 ) | ( ~n16720 & n16922 ) | ( n16723 & n16922 ) ;
  assign n16924 = ( n16720 & n16723 ) | ( n16720 & n16922 ) | ( n16723 & n16922 ) ;
  assign n16925 = ( n16720 & n16923 ) | ( n16720 & ~n16924 ) | ( n16923 & ~n16924 ) ;
  assign n16926 = n40 & n16925 ;
  assign n16927 = n8721 & n16724 ;
  assign n16928 = n8340 & ~n16531 ;
  assign n16929 = n16927 | n16928 ;
  assign n16930 = n16926 | n16929 ;
  assign n16931 = x5 & n16930 ;
  assign n16932 = n16540 & ~n16724 ;
  assign n16933 = n16925 & n16932 ;
  assign n16934 = ( n16734 & ~n16925 ) | ( n16734 & n16932 ) | ( ~n16925 & n16932 ) ;
  assign n16935 = ~n16734 & n16925 ;
  assign n16936 = ( ~n16933 & n16934 ) | ( ~n16933 & n16935 ) | ( n16934 & n16935 ) ;
  assign n16937 = n8341 & ~n16936 ;
  assign n16938 = ( ~x5 & n16930 ) | ( ~x5 & n16937 ) | ( n16930 & n16937 ) ;
  assign n16939 = x5 & ~n16937 ;
  assign n16940 = ( ~n16931 & n16938 ) | ( ~n16931 & n16939 ) | ( n16938 & n16939 ) ;
  assign n16941 = n7644 & ~n16150 ;
  assign n16942 = x8 & n16941 ;
  assign n16943 = n7341 & ~n15954 ;
  assign n16944 = n7345 | n16943 ;
  assign n16945 = ( ~n16338 & n16943 ) | ( ~n16338 & n16944 ) | ( n16943 & n16944 ) ;
  assign n16946 = n7346 | n16945 ;
  assign n16947 = ( ~n16349 & n16945 ) | ( ~n16349 & n16946 ) | ( n16945 & n16946 ) ;
  assign n16948 = x8 & ~n16947 ;
  assign n16949 = ( ~x8 & n16941 ) | ( ~x8 & n16947 ) | ( n16941 & n16947 ) ;
  assign n16950 = ( ~n16942 & n16948 ) | ( ~n16942 & n16949 ) | ( n16948 & n16949 ) ;
  assign n16951 = n6796 & n15561 ;
  assign n16952 = x11 & n16951 ;
  assign n16953 = n6567 & ~n15394 ;
  assign n16954 = n6570 | n16953 ;
  assign n16955 = ( ~n15806 & n16953 ) | ( ~n15806 & n16954 ) | ( n16953 & n16954 ) ;
  assign n16956 = n6571 | n16955 ;
  assign n16957 = ( n15817 & n16955 ) | ( n15817 & n16956 ) | ( n16955 & n16956 ) ;
  assign n16958 = x11 & ~n16957 ;
  assign n16959 = ( ~x11 & n16951 ) | ( ~x11 & n16957 ) | ( n16951 & n16957 ) ;
  assign n16960 = ( ~n16952 & n16958 ) | ( ~n16952 & n16959 ) | ( n16958 & n16959 ) ;
  assign n16961 = n6332 & n14942 ;
  assign n16962 = x14 & n16961 ;
  assign n16963 = n5909 & ~n14723 ;
  assign n16964 = n5914 | n16963 ;
  assign n16965 = ( ~n15184 & n16963 ) | ( ~n15184 & n16964 ) | ( n16963 & n16964 ) ;
  assign n16966 = n5915 | n16965 ;
  assign n16967 = ( ~n15195 & n16965 ) | ( ~n15195 & n16966 ) | ( n16965 & n16966 ) ;
  assign n16968 = x14 & ~n16967 ;
  assign n16969 = ( ~x14 & n16961 ) | ( ~x14 & n16967 ) | ( n16961 & n16967 ) ;
  assign n16970 = ( ~n16962 & n16968 ) | ( ~n16962 & n16969 ) | ( n16968 & n16969 ) ;
  assign n16971 = n5584 & n14352 ;
  assign n16972 = x17 & n16971 ;
  assign n16973 = n5413 & n13992 ;
  assign n16974 = n5417 | n16973 ;
  assign n16975 = ( n14520 & n16973 ) | ( n14520 & n16974 ) | ( n16973 & n16974 ) ;
  assign n16976 = n5418 | n16975 ;
  assign n16977 = ( n14531 & n16975 ) | ( n14531 & n16976 ) | ( n16975 & n16976 ) ;
  assign n16978 = x17 & ~n16977 ;
  assign n16979 = ( ~x17 & n16971 ) | ( ~x17 & n16977 ) | ( n16971 & n16977 ) ;
  assign n16980 = ( ~n16972 & n16978 ) | ( ~n16972 & n16979 ) | ( n16978 & n16979 ) ;
  assign n16981 = n5232 & n13998 ;
  assign n16982 = x20 & n16981 ;
  assign n16983 = n4874 & ~n14000 ;
  assign n16984 = n4878 | n16983 ;
  assign n16985 = ( n13996 & n16983 ) | ( n13996 & n16984 ) | ( n16983 & n16984 ) ;
  assign n16986 = n4879 | n16985 ;
  assign n16987 = ( ~n14130 & n16985 ) | ( ~n14130 & n16986 ) | ( n16985 & n16986 ) ;
  assign n16988 = x20 & ~n16987 ;
  assign n16989 = ( ~x20 & n16981 ) | ( ~x20 & n16987 ) | ( n16981 & n16987 ) ;
  assign n16990 = ( ~n16982 & n16988 ) | ( ~n16982 & n16989 ) | ( n16988 & n16989 ) ;
  assign n16991 = n4584 & ~n14004 ;
  assign n16992 = n4649 | n16991 ;
  assign n16993 = ( ~n14007 & n16991 ) | ( ~n14007 & n16992 ) | ( n16991 & n16992 ) ;
  assign n16994 = n4591 | n16993 ;
  assign n16995 = ( n14066 & n16993 ) | ( n14066 & n16994 ) | ( n16993 & n16994 ) ;
  assign n16996 = n4637 & n14002 ;
  assign n16997 = n16995 | n16996 ;
  assign n16998 = x23 & ~n16603 ;
  assign n16999 = ~n16787 & n16998 ;
  assign n17000 = n16997 & ~n16999 ;
  assign n17001 = n4202 & ~n14014 ;
  assign n17002 = x23 & ~n16999 ;
  assign n17003 = ( n16997 & n17001 ) | ( n16997 & ~n17002 ) | ( n17001 & ~n17002 ) ;
  assign n17004 = ( n16997 & ~n17001 ) | ( n16997 & n17002 ) | ( ~n17001 & n17002 ) ;
  assign n17005 = ( ~n17000 & n17003 ) | ( ~n17000 & n17004 ) | ( n17003 & n17004 ) ;
  assign n17006 = ( ~n16792 & n16990 ) | ( ~n16792 & n17005 ) | ( n16990 & n17005 ) ;
  assign n17007 = ( n16792 & n16990 ) | ( n16792 & n17005 ) | ( n16990 & n17005 ) ;
  assign n17008 = ( n16792 & n17006 ) | ( n16792 & ~n17007 ) | ( n17006 & ~n17007 ) ;
  assign n17009 = ( ~n16795 & n16980 ) | ( ~n16795 & n17008 ) | ( n16980 & n17008 ) ;
  assign n17010 = ( n16795 & n16980 ) | ( n16795 & n17008 ) | ( n16980 & n17008 ) ;
  assign n17011 = ( n16795 & n17009 ) | ( n16795 & ~n17010 ) | ( n17009 & ~n17010 ) ;
  assign n17012 = ( ~n16808 & n16970 ) | ( ~n16808 & n17011 ) | ( n16970 & n17011 ) ;
  assign n17013 = ( n16808 & n16970 ) | ( n16808 & n17011 ) | ( n16970 & n17011 ) ;
  assign n17014 = ( n16808 & n17012 ) | ( n16808 & ~n17013 ) | ( n17012 & ~n17013 ) ;
  assign n17015 = ( ~n16811 & n16960 ) | ( ~n16811 & n17014 ) | ( n16960 & n17014 ) ;
  assign n17016 = ( n16811 & n16960 ) | ( n16811 & n17014 ) | ( n16960 & n17014 ) ;
  assign n17017 = ( n16811 & n17015 ) | ( n16811 & ~n17016 ) | ( n17015 & ~n17016 ) ;
  assign n17018 = ( ~n16814 & n16950 ) | ( ~n16814 & n17017 ) | ( n16950 & n17017 ) ;
  assign n17019 = ( n16814 & n16950 ) | ( n16814 & n17017 ) | ( n16950 & n17017 ) ;
  assign n17020 = ( n16814 & n17018 ) | ( n16814 & ~n17019 ) | ( n17018 & ~n17019 ) ;
  assign n17021 = ( n16816 & n16940 ) | ( n16816 & n17020 ) | ( n16940 & n17020 ) ;
  assign n17022 = n4591 & n12756 ;
  assign n17023 = x23 & n17022 ;
  assign n17024 = n4649 & ~n10237 ;
  assign n17025 = n4637 & ~n10332 ;
  assign n17026 = n4584 & n10329 ;
  assign n17027 = n17025 | n17026 ;
  assign n17028 = n17024 | n17027 ;
  assign n17029 = x23 & ~n17028 ;
  assign n17030 = ( ~x23 & n17022 ) | ( ~x23 & n17028 ) | ( n17022 & n17028 ) ;
  assign n17031 = ( ~n17023 & n17029 ) | ( ~n17023 & n17030 ) | ( n17029 & n17030 ) ;
  assign n17032 = n4215 & n10326 ;
  assign n17033 = n4200 & n10239 ;
  assign n17034 = n2083 & n10241 ;
  assign n17035 = n17033 | n17034 ;
  assign n17036 = n17032 | n17035 ;
  assign n17037 = x26 & n17036 ;
  assign n17038 = n4203 & n12222 ;
  assign n17039 = ( ~x26 & n17036 ) | ( ~x26 & n17038 ) | ( n17036 & n17038 ) ;
  assign n17040 = x26 & ~n17038 ;
  assign n17041 = ( ~n17037 & n17039 ) | ( ~n17037 & n17040 ) | ( n17039 & n17040 ) ;
  assign n17042 = x26 & ~n16853 ;
  assign n17043 = ~x26 & n16853 ;
  assign n17044 = n17042 | n17043 ;
  assign n17045 = x29 & ~n16860 ;
  assign n17046 = ~x29 & n16860 ;
  assign n17047 = n17045 | n17046 ;
  assign n17048 = ( n16907 & n17044 ) | ( n16907 & n17047 ) | ( n17044 & n17047 ) ;
  assign n17049 = n3541 & ~n11989 ;
  assign n17050 = x29 & n17049 ;
  assign n17051 = n4039 & n10243 ;
  assign n17052 = n3501 & ~n10320 ;
  assign n17053 = n3536 & n10245 ;
  assign n17054 = n17052 | n17053 ;
  assign n17055 = n17051 | n17054 ;
  assign n17056 = x29 & ~n17055 ;
  assign n17057 = ( ~x29 & n17049 ) | ( ~x29 & n17055 ) | ( n17049 & n17055 ) ;
  assign n17058 = ( ~n17050 & n17056 ) | ( ~n17050 & n17057 ) | ( n17056 & n17057 ) ;
  assign n17059 = n3273 & n10312 ;
  assign n17060 = n3270 | n17059 ;
  assign n17061 = ( ~n10316 & n17059 ) | ( ~n10316 & n17060 ) | ( n17059 & n17060 ) ;
  assign n17062 = n390 | n17061 ;
  assign n17063 = ( ~n11691 & n17061 ) | ( ~n11691 & n17062 ) | ( n17061 & n17062 ) ;
  assign n17064 = n3274 & n10247 ;
  assign n17065 = n17063 | n17064 ;
  assign n17066 = n2301 & ~n6188 ;
  assign n17067 = n4478 | n15125 ;
  assign n17068 = n3983 | n17067 ;
  assign n17069 = n323 | n442 ;
  assign n17070 = n87 | n17069 ;
  assign n17071 = n984 | n17070 ;
  assign n17072 = n1273 | n17071 ;
  assign n17073 = n17068 | n17072 ;
  assign n17074 = n669 | n915 ;
  assign n17075 = n1253 | n1998 ;
  assign n17076 = n17074 | n17075 ;
  assign n17077 = n13586 | n17076 ;
  assign n17078 = n2092 | n4384 ;
  assign n17079 = n14844 | n17078 ;
  assign n17080 = n17077 | n17079 ;
  assign n17081 = n2341 | n17080 ;
  assign n17082 = n17073 | n17081 ;
  assign n17083 = n17066 & ~n17082 ;
  assign n17084 = ( n16624 & n16700 ) | ( n16624 & ~n17083 ) | ( n16700 & ~n17083 ) ;
  assign n17085 = ( n16624 & ~n16700 ) | ( n16624 & n17083 ) | ( ~n16700 & n17083 ) ;
  assign n17086 = ( ~n16624 & n17084 ) | ( ~n16624 & n17085 ) | ( n17084 & n17085 ) ;
  assign n17087 = ( ~n16902 & n17065 ) | ( ~n16902 & n17086 ) | ( n17065 & n17086 ) ;
  assign n17088 = ( n16902 & n17065 ) | ( n16902 & n17086 ) | ( n17065 & n17086 ) ;
  assign n17089 = ( n16902 & n17087 ) | ( n16902 & ~n17088 ) | ( n17087 & ~n17088 ) ;
  assign n17090 = ( n16906 & n17058 ) | ( n16906 & n17089 ) | ( n17058 & n17089 ) ;
  assign n17091 = ( ~n16906 & n17058 ) | ( ~n16906 & n17089 ) | ( n17058 & n17089 ) ;
  assign n17092 = ( n16906 & ~n17090 ) | ( n16906 & n17091 ) | ( ~n17090 & n17091 ) ;
  assign n17093 = ( n17041 & n17048 ) | ( n17041 & ~n17092 ) | ( n17048 & ~n17092 ) ;
  assign n17094 = ( n17041 & ~n17048 ) | ( n17041 & n17092 ) | ( ~n17048 & n17092 ) ;
  assign n17095 = ( ~n17041 & n17093 ) | ( ~n17041 & n17094 ) | ( n17093 & n17094 ) ;
  assign n17096 = ( n16912 & ~n17031 ) | ( n16912 & n17095 ) | ( ~n17031 & n17095 ) ;
  assign n17097 = ( n16912 & n17031 ) | ( n16912 & ~n17095 ) | ( n17031 & ~n17095 ) ;
  assign n17098 = ( ~n16912 & n17096 ) | ( ~n16912 & n17097 ) | ( n17096 & n17097 ) ;
  assign n17099 = n5232 & ~n10235 ;
  assign n17100 = x20 & n17099 ;
  assign n17101 = n4874 & n10214 ;
  assign n17102 = n4878 | n17101 ;
  assign n17103 = ( ~n13280 & n17101 ) | ( ~n13280 & n17102 ) | ( n17101 & n17102 ) ;
  assign n17104 = n4879 | n17103 ;
  assign n17105 = ( ~n13285 & n17103 ) | ( ~n13285 & n17104 ) | ( n17103 & n17104 ) ;
  assign n17106 = x20 & ~n17105 ;
  assign n17107 = ( ~x20 & n17099 ) | ( ~x20 & n17105 ) | ( n17099 & n17105 ) ;
  assign n17108 = ( ~n17100 & n17106 ) | ( ~n17100 & n17107 ) | ( n17106 & n17107 ) ;
  assign n17109 = ( n16914 & n17098 ) | ( n16914 & ~n17108 ) | ( n17098 & ~n17108 ) ;
  assign n17110 = ( n16914 & ~n17098 ) | ( n16914 & n17108 ) | ( ~n17098 & n17108 ) ;
  assign n17111 = ( ~n16914 & n17109 ) | ( ~n16914 & n17110 ) | ( n17109 & n17110 ) ;
  assign n17112 = n5413 | n5417 ;
  assign n17113 = ( n5417 & ~n13473 ) | ( n5417 & n17112 ) | ( ~n13473 & n17112 ) ;
  assign n17114 = n5584 | n17113 ;
  assign n17115 = ( n13475 & n17113 ) | ( n13475 & n17114 ) | ( n17113 & n17114 ) ;
  assign n17116 = x17 & n17115 ;
  assign n17117 = n5414 & n13477 ;
  assign n17118 = x17 & ~n17117 ;
  assign n17119 = ( ~x17 & n17115 ) | ( ~x17 & n17117 ) | ( n17115 & n17117 ) ;
  assign n17120 = ( ~n17116 & n17118 ) | ( ~n17116 & n17119 ) | ( n17118 & n17119 ) ;
  assign n17121 = ( n16918 & ~n17111 ) | ( n16918 & n17120 ) | ( ~n17111 & n17120 ) ;
  assign n17122 = ( n16918 & n17111 ) | ( n16918 & ~n17120 ) | ( n17111 & ~n17120 ) ;
  assign n17123 = ( ~n16918 & n17121 ) | ( ~n16918 & n17122 ) | ( n17121 & n17122 ) ;
  assign n17124 = ( ~n16921 & n16924 ) | ( ~n16921 & n17123 ) | ( n16924 & n17123 ) ;
  assign n17125 = ( n16921 & n16924 ) | ( n16921 & ~n17123 ) | ( n16924 & ~n17123 ) ;
  assign n17126 = ( ~n16924 & n17124 ) | ( ~n16924 & n17125 ) | ( n17124 & n17125 ) ;
  assign n17127 = n40 & ~n17126 ;
  assign n17128 = n8721 & n16925 ;
  assign n17129 = n8340 & n16724 ;
  assign n17130 = n17128 | n17129 ;
  assign n17131 = n17127 | n17130 ;
  assign n17132 = x5 & n17131 ;
  assign n17133 = n16734 | n16925 ;
  assign n17134 = n16925 & ~n16932 ;
  assign n17135 = n17126 & ~n17134 ;
  assign n17136 = n17133 & n17135 ;
  assign n17137 = ~n17126 & n17133 ;
  assign n17138 = ( ~n16925 & n16933 ) | ( ~n16925 & n17137 ) | ( n16933 & n17137 ) ;
  assign n17139 = ( n17126 & ~n17136 ) | ( n17126 & n17138 ) | ( ~n17136 & n17138 ) ;
  assign n17140 = n8341 & ~n17139 ;
  assign n17141 = ( ~x5 & n17131 ) | ( ~x5 & n17140 ) | ( n17131 & n17140 ) ;
  assign n17142 = x5 & ~n17140 ;
  assign n17143 = ( ~n17132 & n17141 ) | ( ~n17132 & n17142 ) | ( n17141 & n17142 ) ;
  assign n17144 = n7346 & ~n16542 ;
  assign n17145 = x8 & n17144 ;
  assign n17146 = n7341 & ~n16150 ;
  assign n17147 = n7345 | n17146 ;
  assign n17148 = ( ~n16531 & n17146 ) | ( ~n16531 & n17147 ) | ( n17146 & n17147 ) ;
  assign n17149 = n7644 & ~n16338 ;
  assign n17150 = n17148 | n17149 ;
  assign n17151 = x8 & ~n17150 ;
  assign n17152 = ( ~x8 & n17144 ) | ( ~x8 & n17150 ) | ( n17144 & n17150 ) ;
  assign n17153 = ( ~n17145 & n17151 ) | ( ~n17145 & n17152 ) | ( n17151 & n17152 ) ;
  assign n17154 = n6796 & ~n15806 ;
  assign n17155 = x11 & n17154 ;
  assign n17156 = n6567 & n15561 ;
  assign n17157 = n6570 | n17156 ;
  assign n17158 = ( ~n15954 & n17156 ) | ( ~n15954 & n17157 ) | ( n17156 & n17157 ) ;
  assign n17159 = n6571 | n17158 ;
  assign n17160 = ( ~n15965 & n17158 ) | ( ~n15965 & n17159 ) | ( n17158 & n17159 ) ;
  assign n17161 = x11 & ~n17160 ;
  assign n17162 = ( ~x11 & n17154 ) | ( ~x11 & n17160 ) | ( n17154 & n17160 ) ;
  assign n17163 = ( ~n17155 & n17161 ) | ( ~n17155 & n17162 ) | ( n17161 & n17162 ) ;
  assign n17164 = n6332 & ~n15184 ;
  assign n17165 = x14 & n17164 ;
  assign n17166 = n5909 & n14942 ;
  assign n17167 = n5914 | n17166 ;
  assign n17168 = ( ~n15394 & n17166 ) | ( ~n15394 & n17167 ) | ( n17166 & n17167 ) ;
  assign n17169 = n5915 | n17168 ;
  assign n17170 = ( n15405 & n17168 ) | ( n15405 & n17169 ) | ( n17168 & n17169 ) ;
  assign n17171 = x14 & ~n17170 ;
  assign n17172 = ( ~x14 & n17164 ) | ( ~x14 & n17170 ) | ( n17164 & n17170 ) ;
  assign n17173 = ( ~n17165 & n17171 ) | ( ~n17165 & n17172 ) | ( n17171 & n17172 ) ;
  assign n17174 = n5584 & n14520 ;
  assign n17175 = x17 & n17174 ;
  assign n17176 = n5413 & n14352 ;
  assign n17177 = n5417 | n17176 ;
  assign n17178 = ( ~n14723 & n17176 ) | ( ~n14723 & n17177 ) | ( n17176 & n17177 ) ;
  assign n17179 = n5418 | n17178 ;
  assign n17180 = ( ~n14734 & n17178 ) | ( ~n14734 & n17179 ) | ( n17178 & n17179 ) ;
  assign n17181 = x17 & ~n17180 ;
  assign n17182 = ( ~x17 & n17174 ) | ( ~x17 & n17180 ) | ( n17174 & n17180 ) ;
  assign n17183 = ( ~n17175 & n17181 ) | ( ~n17175 & n17182 ) | ( n17181 & n17182 ) ;
  assign n17184 = n4878 & n13992 ;
  assign n17185 = n5232 & n13996 ;
  assign n17186 = n4874 & n13998 ;
  assign n17187 = n17185 | n17186 ;
  assign n17188 = n17184 | n17187 ;
  assign n17189 = x20 & n17188 ;
  assign n17190 = n4879 & n14024 ;
  assign n17191 = x20 & ~n17190 ;
  assign n17192 = ( ~x20 & n17188 ) | ( ~x20 & n17190 ) | ( n17188 & n17190 ) ;
  assign n17193 = ( ~n17189 & n17191 ) | ( ~n17189 & n17192 ) | ( n17191 & n17192 ) ;
  assign n17194 = n4637 & ~n14007 ;
  assign n17195 = x23 & n17194 ;
  assign n17196 = n4584 & n14002 ;
  assign n17197 = n4649 | n17196 ;
  assign n17198 = ( ~n14000 & n17196 ) | ( ~n14000 & n17197 ) | ( n17196 & n17197 ) ;
  assign n17199 = n4591 | n17198 ;
  assign n17200 = ( ~n14042 & n17198 ) | ( ~n14042 & n17199 ) | ( n17198 & n17199 ) ;
  assign n17201 = x23 & ~n17200 ;
  assign n17202 = ( ~x23 & n17194 ) | ( ~x23 & n17200 ) | ( n17194 & n17200 ) ;
  assign n17203 = ( ~n17195 & n17201 ) | ( ~n17195 & n17202 ) | ( n17201 & n17202 ) ;
  assign n17204 = x23 & ~n16997 ;
  assign n17205 = ( n17000 & ~n17004 ) | ( n17000 & n17204 ) | ( ~n17004 & n17204 ) ;
  assign n17206 = n4203 & n14004 ;
  assign n17207 = n4200 & ~n14014 ;
  assign n17208 = ( ~n14014 & n17206 ) | ( ~n14014 & n17207 ) | ( n17206 & n17207 ) ;
  assign n17209 = ( n4202 & n4215 ) | ( n4202 & n14014 ) | ( n4215 & n14014 ) ;
  assign n17210 = ~n14004 & n17209 ;
  assign n17211 = n17208 | n17210 ;
  assign n17212 = n17001 | n17211 ;
  assign n17213 = ( x26 & n17001 ) | ( x26 & ~n17211 ) | ( n17001 & ~n17211 ) ;
  assign n17214 = x26 & ~n17211 ;
  assign n17215 = ( n17212 & ~n17213 ) | ( n17212 & n17214 ) | ( ~n17213 & n17214 ) ;
  assign n17216 = ( n17203 & n17205 ) | ( n17203 & n17215 ) | ( n17205 & n17215 ) ;
  assign n17217 = ( ~n17203 & n17205 ) | ( ~n17203 & n17215 ) | ( n17205 & n17215 ) ;
  assign n17218 = ( n17203 & ~n17216 ) | ( n17203 & n17217 ) | ( ~n17216 & n17217 ) ;
  assign n17219 = ( ~n17007 & n17193 ) | ( ~n17007 & n17218 ) | ( n17193 & n17218 ) ;
  assign n17220 = ( n17007 & n17193 ) | ( n17007 & n17218 ) | ( n17193 & n17218 ) ;
  assign n17221 = ( n17007 & n17219 ) | ( n17007 & ~n17220 ) | ( n17219 & ~n17220 ) ;
  assign n17222 = ( ~n17010 & n17183 ) | ( ~n17010 & n17221 ) | ( n17183 & n17221 ) ;
  assign n17223 = ( n17010 & n17183 ) | ( n17010 & n17221 ) | ( n17183 & n17221 ) ;
  assign n17224 = ( n17010 & n17222 ) | ( n17010 & ~n17223 ) | ( n17222 & ~n17223 ) ;
  assign n17225 = ( ~n17013 & n17173 ) | ( ~n17013 & n17224 ) | ( n17173 & n17224 ) ;
  assign n17226 = ( n17013 & n17173 ) | ( n17013 & n17224 ) | ( n17173 & n17224 ) ;
  assign n17227 = ( n17013 & n17225 ) | ( n17013 & ~n17226 ) | ( n17225 & ~n17226 ) ;
  assign n17228 = ( ~n17016 & n17163 ) | ( ~n17016 & n17227 ) | ( n17163 & n17227 ) ;
  assign n17229 = ( n17016 & n17163 ) | ( n17016 & n17227 ) | ( n17163 & n17227 ) ;
  assign n17230 = ( n17016 & n17228 ) | ( n17016 & ~n17229 ) | ( n17228 & ~n17229 ) ;
  assign n17231 = ( ~n17019 & n17153 ) | ( ~n17019 & n17230 ) | ( n17153 & n17230 ) ;
  assign n17232 = ( n17019 & n17153 ) | ( n17019 & n17230 ) | ( n17153 & n17230 ) ;
  assign n17233 = ( n17019 & n17231 ) | ( n17019 & ~n17232 ) | ( n17231 & ~n17232 ) ;
  assign n17234 = ( n17021 & n17143 ) | ( n17021 & n17233 ) | ( n17143 & n17233 ) ;
  assign n17235 = n5232 & ~n13280 ;
  assign n17236 = x20 & n17235 ;
  assign n17237 = n4878 & ~n13473 ;
  assign n17238 = n4874 & ~n10235 ;
  assign n17239 = n17237 | n17238 ;
  assign n17240 = n4879 | n17239 ;
  assign n17241 = ( ~n13480 & n17239 ) | ( ~n13480 & n17240 ) | ( n17239 & n17240 ) ;
  assign n17242 = x20 & ~n17241 ;
  assign n17243 = ( ~x20 & n17235 ) | ( ~x20 & n17241 ) | ( n17235 & n17241 ) ;
  assign n17244 = ( ~n17236 & n17242 ) | ( ~n17236 & n17243 ) | ( n17242 & n17243 ) ;
  assign n17245 = n4637 & ~n10237 ;
  assign n17246 = x23 & n17245 ;
  assign n17247 = n4584 & ~n10332 ;
  assign n17248 = n4649 | n17247 ;
  assign n17249 = ( n10214 & n17247 ) | ( n10214 & n17248 ) | ( n17247 & n17248 ) ;
  assign n17250 = n4591 | n17249 ;
  assign n17251 = ( n12953 & n17249 ) | ( n12953 & n17250 ) | ( n17249 & n17250 ) ;
  assign n17252 = x23 & ~n17251 ;
  assign n17253 = ( ~x23 & n17245 ) | ( ~x23 & n17251 ) | ( n17245 & n17251 ) ;
  assign n17254 = ( ~n17246 & n17252 ) | ( ~n17246 & n17253 ) | ( n17252 & n17253 ) ;
  assign n17255 = n4215 & n10329 ;
  assign n17256 = n4200 & n10326 ;
  assign n17257 = n2083 & n10239 ;
  assign n17258 = n17256 | n17257 ;
  assign n17259 = n17255 | n17258 ;
  assign n17260 = x26 & n17259 ;
  assign n17261 = n4203 & n10397 ;
  assign n17262 = ( ~x26 & n17259 ) | ( ~x26 & n17261 ) | ( n17259 & n17261 ) ;
  assign n17263 = x26 & ~n17261 ;
  assign n17264 = ( ~n17260 & n17262 ) | ( ~n17260 & n17263 ) | ( n17262 & n17263 ) ;
  assign n17265 = n3501 & n10243 ;
  assign n17266 = x29 & n17265 ;
  assign n17267 = n3536 & ~n10320 ;
  assign n17268 = n4039 | n17267 ;
  assign n17269 = ( n10241 & n17267 ) | ( n10241 & n17268 ) | ( n17267 & n17268 ) ;
  assign n17270 = n3541 | n17269 ;
  assign n17271 = ( n12105 & n17269 ) | ( n12105 & n17270 ) | ( n17269 & n17270 ) ;
  assign n17272 = x29 & ~n17271 ;
  assign n17273 = ( ~x29 & n17265 ) | ( ~x29 & n17271 ) | ( n17265 & n17271 ) ;
  assign n17274 = ( ~n17266 & n17272 ) | ( ~n17266 & n17273 ) | ( n17272 & n17273 ) ;
  assign n17275 = n294 | n916 ;
  assign n17276 = n323 | n689 ;
  assign n17277 = n17275 | n17276 ;
  assign n17278 = n876 | n15763 ;
  assign n17279 = n17277 | n17278 ;
  assign n17280 = n5662 | n17279 ;
  assign n17281 = n431 | n922 ;
  assign n17282 = n477 | n647 ;
  assign n17283 = n17281 | n17282 ;
  assign n17284 = n3427 | n17283 ;
  assign n17285 = n17280 | n17284 ;
  assign n17286 = n2351 | n3116 ;
  assign n17287 = n14882 | n17286 ;
  assign n17288 = n17285 | n17287 ;
  assign n17289 = n4370 | n17288 ;
  assign n17290 = n151 | n3032 ;
  assign n17291 = n17289 | n17290 ;
  assign n17292 = n419 | n533 ;
  assign n17293 = n1914 | n17292 ;
  assign n17294 = n2413 | n17293 ;
  assign n17295 = n137 | n17294 ;
  assign n17296 = n2105 | n2917 ;
  assign n17297 = n5952 | n17296 ;
  assign n17298 = n17295 | n17297 ;
  assign n17299 = n735 | n2448 ;
  assign n17300 = n574 | n1126 ;
  assign n17301 = n17299 | n17300 ;
  assign n17302 = n17298 | n17301 ;
  assign n17303 = n1064 | n3022 ;
  assign n17304 = n268 | n372 ;
  assign n17305 = n1263 | n17304 ;
  assign n17306 = n17303 | n17305 ;
  assign n17307 = n1849 | n3206 ;
  assign n17308 = n393 | n17307 ;
  assign n17309 = n17306 | n17308 ;
  assign n17310 = n17302 | n17309 ;
  assign n17311 = n3200 | n17310 ;
  assign n17312 = n17291 | n17311 ;
  assign n17313 = n3273 & n10247 ;
  assign n17314 = n3270 | n17313 ;
  assign n17315 = ( n10245 & n17313 ) | ( n10245 & n17314 ) | ( n17313 & n17314 ) ;
  assign n17316 = n390 | n17315 ;
  assign n17317 = ( ~n11676 & n17315 ) | ( ~n11676 & n17316 ) | ( n17315 & n17316 ) ;
  assign n17318 = n3274 & ~n10316 ;
  assign n17319 = n17317 | n17318 ;
  assign n17320 = ( n17085 & n17312 ) | ( n17085 & n17319 ) | ( n17312 & n17319 ) ;
  assign n17321 = ( n17085 & ~n17312 ) | ( n17085 & n17319 ) | ( ~n17312 & n17319 ) ;
  assign n17322 = ( n17312 & ~n17320 ) | ( n17312 & n17321 ) | ( ~n17320 & n17321 ) ;
  assign n17323 = ( n17088 & ~n17274 ) | ( n17088 & n17322 ) | ( ~n17274 & n17322 ) ;
  assign n17324 = ( n17088 & n17274 ) | ( n17088 & n17322 ) | ( n17274 & n17322 ) ;
  assign n17325 = ( n17274 & n17323 ) | ( n17274 & ~n17324 ) | ( n17323 & ~n17324 ) ;
  assign n17326 = ( n17091 & n17264 ) | ( n17091 & n17325 ) | ( n17264 & n17325 ) ;
  assign n17327 = ( n17091 & ~n17264 ) | ( n17091 & n17325 ) | ( ~n17264 & n17325 ) ;
  assign n17328 = ( n17264 & ~n17326 ) | ( n17264 & n17327 ) | ( ~n17326 & n17327 ) ;
  assign n17329 = ( n17093 & ~n17254 ) | ( n17093 & n17328 ) | ( ~n17254 & n17328 ) ;
  assign n17330 = ( n17093 & n17254 ) | ( n17093 & n17328 ) | ( n17254 & n17328 ) ;
  assign n17331 = ( n17254 & n17329 ) | ( n17254 & ~n17330 ) | ( n17329 & ~n17330 ) ;
  assign n17332 = ( n17097 & ~n17244 ) | ( n17097 & n17331 ) | ( ~n17244 & n17331 ) ;
  assign n17333 = ( n17097 & n17244 ) | ( n17097 & n17331 ) | ( n17244 & n17331 ) ;
  assign n17334 = ( n17244 & n17332 ) | ( n17244 & ~n17333 ) | ( n17332 & ~n17333 ) ;
  assign n17335 = ( x14 & ~x15 ) | ( x14 & x16 ) | ( ~x15 & x16 ) ;
  assign n17336 = ( x15 & ~x17 ) | ( x15 & n17335 ) | ( ~x17 & n17335 ) ;
  assign n17337 = ~n5412 & n17336 ;
  assign n17338 = ( n13475 & n17336 ) | ( n13475 & n17337 ) | ( n17336 & n17337 ) ;
  assign n17339 = n5409 & ~n13475 ;
  assign n17340 = n17338 | n17339 ;
  assign n17341 = ( ~n17110 & n17334 ) | ( ~n17110 & n17340 ) | ( n17334 & n17340 ) ;
  assign n17342 = ( n17110 & n17334 ) | ( n17110 & n17340 ) | ( n17334 & n17340 ) ;
  assign n17343 = ( n17110 & n17341 ) | ( n17110 & ~n17342 ) | ( n17341 & ~n17342 ) ;
  assign n17344 = ( ~n17121 & n17125 ) | ( ~n17121 & n17343 ) | ( n17125 & n17343 ) ;
  assign n17345 = ( n17121 & n17125 ) | ( n17121 & n17343 ) | ( n17125 & n17343 ) ;
  assign n17346 = ( n17121 & n17344 ) | ( n17121 & ~n17345 ) | ( n17344 & ~n17345 ) ;
  assign n17347 = n40 & n17346 ;
  assign n17348 = n8721 & ~n17126 ;
  assign n17349 = n8340 & n16925 ;
  assign n17350 = n17348 | n17349 ;
  assign n17351 = n17347 | n17350 ;
  assign n17352 = x5 & n17351 ;
  assign n17353 = n17137 & n17346 ;
  assign n17354 = ~n17135 & n17346 ;
  assign n17355 = ( n17135 & n17137 ) | ( n17135 & ~n17346 ) | ( n17137 & ~n17346 ) ;
  assign n17356 = ( ~n17353 & n17354 ) | ( ~n17353 & n17355 ) | ( n17354 & n17355 ) ;
  assign n17357 = n8341 & ~n17356 ;
  assign n17358 = ( ~x5 & n17351 ) | ( ~x5 & n17357 ) | ( n17351 & n17357 ) ;
  assign n17359 = x5 & ~n17357 ;
  assign n17360 = ( ~n17352 & n17358 ) | ( ~n17352 & n17359 ) | ( n17358 & n17359 ) ;
  assign n17361 = n7345 & n16724 ;
  assign n17362 = n7644 & ~n16531 ;
  assign n17363 = n7341 & ~n16338 ;
  assign n17364 = n17362 | n17363 ;
  assign n17365 = n17361 | n17364 ;
  assign n17366 = x8 & n17365 ;
  assign n17367 = n7346 & n16735 ;
  assign n17368 = ( ~x8 & n17365 ) | ( ~x8 & n17367 ) | ( n17365 & n17367 ) ;
  assign n17369 = x8 & ~n17367 ;
  assign n17370 = ( ~n17366 & n17368 ) | ( ~n17366 & n17369 ) | ( n17368 & n17369 ) ;
  assign n17371 = n6571 & ~n16161 ;
  assign n17372 = x11 & n17371 ;
  assign n17373 = n6567 & ~n15806 ;
  assign n17374 = n6570 | n17373 ;
  assign n17375 = ( ~n16150 & n17373 ) | ( ~n16150 & n17374 ) | ( n17373 & n17374 ) ;
  assign n17376 = n6796 & ~n15954 ;
  assign n17377 = n17375 | n17376 ;
  assign n17378 = x11 & ~n17377 ;
  assign n17379 = ( ~x11 & n17371 ) | ( ~x11 & n17377 ) | ( n17371 & n17377 ) ;
  assign n17380 = ( ~n17372 & n17378 ) | ( ~n17372 & n17379 ) | ( n17378 & n17379 ) ;
  assign n17381 = n6332 & ~n15394 ;
  assign n17382 = x14 & n17381 ;
  assign n17383 = n5909 & ~n15184 ;
  assign n17384 = n5914 | n17383 ;
  assign n17385 = ( n15561 & n17383 ) | ( n15561 & n17384 ) | ( n17383 & n17384 ) ;
  assign n17386 = n5915 | n17385 ;
  assign n17387 = ( n15573 & n17385 ) | ( n15573 & n17386 ) | ( n17385 & n17386 ) ;
  assign n17388 = x14 & ~n17387 ;
  assign n17389 = ( ~x14 & n17381 ) | ( ~x14 & n17387 ) | ( n17381 & n17387 ) ;
  assign n17390 = ( ~n17382 & n17388 ) | ( ~n17382 & n17389 ) | ( n17388 & n17389 ) ;
  assign n17391 = n5584 & ~n14723 ;
  assign n17392 = x17 & n17391 ;
  assign n17393 = n5413 & n14520 ;
  assign n17394 = n5417 | n17393 ;
  assign n17395 = ( n14942 & n17393 ) | ( n14942 & n17394 ) | ( n17393 & n17394 ) ;
  assign n17396 = n5418 | n17395 ;
  assign n17397 = ( ~n14953 & n17395 ) | ( ~n14953 & n17396 ) | ( n17395 & n17396 ) ;
  assign n17398 = x17 & ~n17397 ;
  assign n17399 = ( ~x17 & n17391 ) | ( ~x17 & n17397 ) | ( n17391 & n17397 ) ;
  assign n17400 = ( ~n17392 & n17398 ) | ( ~n17392 & n17399 ) | ( n17398 & n17399 ) ;
  assign n17401 = n5232 & n13992 ;
  assign n17402 = x20 & n17401 ;
  assign n17403 = n4874 & n13996 ;
  assign n17404 = n4878 | n17403 ;
  assign n17405 = ( n14352 & n17403 ) | ( n14352 & n17404 ) | ( n17403 & n17404 ) ;
  assign n17406 = n4879 | n17405 ;
  assign n17407 = ( n14363 & n17405 ) | ( n14363 & n17406 ) | ( n17405 & n17406 ) ;
  assign n17408 = x20 & ~n17407 ;
  assign n17409 = ( ~x20 & n17401 ) | ( ~x20 & n17407 ) | ( n17401 & n17407 ) ;
  assign n17410 = ( ~n17402 & n17408 ) | ( ~n17402 & n17409 ) | ( n17408 & n17409 ) ;
  assign n17411 = n4637 & ~n14000 ;
  assign n17412 = x23 & n17411 ;
  assign n17413 = n4584 & ~n14007 ;
  assign n17414 = n4649 | n17413 ;
  assign n17415 = ( n13998 & n17413 ) | ( n13998 & n17414 ) | ( n17413 & n17414 ) ;
  assign n17416 = n4591 | n17415 ;
  assign n17417 = ( n14115 & n17415 ) | ( n14115 & n17416 ) | ( n17415 & n17416 ) ;
  assign n17418 = x23 & ~n17417 ;
  assign n17419 = ( ~x23 & n17411 ) | ( ~x23 & n17417 ) | ( n17411 & n17417 ) ;
  assign n17420 = ( ~n17412 & n17418 ) | ( ~n17412 & n17419 ) | ( n17418 & n17419 ) ;
  assign n17421 = x26 & n17212 ;
  assign n17422 = n4200 & ~n14004 ;
  assign n17423 = n2083 & ~n14014 ;
  assign n17424 = n17422 | n17423 ;
  assign n17425 = n4203 | n17424 ;
  assign n17426 = ( n14072 & n17424 ) | ( n14072 & n17425 ) | ( n17424 & n17425 ) ;
  assign n17427 = n4215 & n14002 ;
  assign n17428 = n17426 | n17427 ;
  assign n17429 = n17421 & ~n17428 ;
  assign n17430 = ~n17421 & n17428 ;
  assign n17431 = n17429 | n17430 ;
  assign n17432 = ( ~n17216 & n17420 ) | ( ~n17216 & n17431 ) | ( n17420 & n17431 ) ;
  assign n17433 = ( n17216 & n17420 ) | ( n17216 & n17431 ) | ( n17420 & n17431 ) ;
  assign n17434 = ( n17216 & n17432 ) | ( n17216 & ~n17433 ) | ( n17432 & ~n17433 ) ;
  assign n17435 = ( n17220 & n17410 ) | ( n17220 & n17434 ) | ( n17410 & n17434 ) ;
  assign n17436 = ( ~n17220 & n17410 ) | ( ~n17220 & n17434 ) | ( n17410 & n17434 ) ;
  assign n17437 = ( n17220 & ~n17435 ) | ( n17220 & n17436 ) | ( ~n17435 & n17436 ) ;
  assign n17438 = ( ~n17223 & n17400 ) | ( ~n17223 & n17437 ) | ( n17400 & n17437 ) ;
  assign n17439 = ( n17223 & n17400 ) | ( n17223 & n17437 ) | ( n17400 & n17437 ) ;
  assign n17440 = ( n17223 & n17438 ) | ( n17223 & ~n17439 ) | ( n17438 & ~n17439 ) ;
  assign n17441 = ( ~n17226 & n17390 ) | ( ~n17226 & n17440 ) | ( n17390 & n17440 ) ;
  assign n17442 = ( n17226 & n17390 ) | ( n17226 & n17440 ) | ( n17390 & n17440 ) ;
  assign n17443 = ( n17226 & n17441 ) | ( n17226 & ~n17442 ) | ( n17441 & ~n17442 ) ;
  assign n17444 = ( ~n17229 & n17380 ) | ( ~n17229 & n17443 ) | ( n17380 & n17443 ) ;
  assign n17445 = ( n17229 & n17380 ) | ( n17229 & n17443 ) | ( n17380 & n17443 ) ;
  assign n17446 = ( n17229 & n17444 ) | ( n17229 & ~n17445 ) | ( n17444 & ~n17445 ) ;
  assign n17447 = ( ~n17232 & n17370 ) | ( ~n17232 & n17446 ) | ( n17370 & n17446 ) ;
  assign n17448 = ( n17232 & n17370 ) | ( n17232 & n17446 ) | ( n17370 & n17446 ) ;
  assign n17449 = ( n17232 & n17447 ) | ( n17232 & ~n17448 ) | ( n17447 & ~n17448 ) ;
  assign n17450 = ( n17234 & n17360 ) | ( n17234 & n17449 ) | ( n17360 & n17449 ) ;
  assign n17451 = n7644 & n16724 ;
  assign n17452 = x8 & n17451 ;
  assign n17453 = n7341 & ~n16531 ;
  assign n17454 = n7345 | n17453 ;
  assign n17455 = ( n16925 & n17453 ) | ( n16925 & n17454 ) | ( n17453 & n17454 ) ;
  assign n17456 = n7346 | n17455 ;
  assign n17457 = ( ~n16936 & n17455 ) | ( ~n16936 & n17456 ) | ( n17455 & n17456 ) ;
  assign n17458 = x8 & ~n17457 ;
  assign n17459 = ( ~x8 & n17451 ) | ( ~x8 & n17457 ) | ( n17451 & n17457 ) ;
  assign n17460 = ( ~n17452 & n17458 ) | ( ~n17452 & n17459 ) | ( n17458 & n17459 ) ;
  assign n17461 = n6796 & ~n16150 ;
  assign n17462 = x11 & n17461 ;
  assign n17463 = n6567 & ~n15954 ;
  assign n17464 = n6570 | n17463 ;
  assign n17465 = ( ~n16338 & n17463 ) | ( ~n16338 & n17464 ) | ( n17463 & n17464 ) ;
  assign n17466 = n6571 | n17465 ;
  assign n17467 = ( ~n16349 & n17465 ) | ( ~n16349 & n17466 ) | ( n17465 & n17466 ) ;
  assign n17468 = x11 & ~n17467 ;
  assign n17469 = ( ~x11 & n17461 ) | ( ~x11 & n17467 ) | ( n17461 & n17467 ) ;
  assign n17470 = ( ~n17462 & n17468 ) | ( ~n17462 & n17469 ) | ( n17468 & n17469 ) ;
  assign n17471 = n6332 & n15561 ;
  assign n17472 = x14 & n17471 ;
  assign n17473 = n5909 & ~n15394 ;
  assign n17474 = n5914 | n17473 ;
  assign n17475 = ( ~n15806 & n17473 ) | ( ~n15806 & n17474 ) | ( n17473 & n17474 ) ;
  assign n17476 = n5915 | n17475 ;
  assign n17477 = ( n15817 & n17475 ) | ( n15817 & n17476 ) | ( n17475 & n17476 ) ;
  assign n17478 = x14 & ~n17477 ;
  assign n17479 = ( ~x14 & n17471 ) | ( ~x14 & n17477 ) | ( n17471 & n17477 ) ;
  assign n17480 = ( ~n17472 & n17478 ) | ( ~n17472 & n17479 ) | ( n17478 & n17479 ) ;
  assign n17481 = n5584 & n14942 ;
  assign n17482 = x17 & n17481 ;
  assign n17483 = n5413 & ~n14723 ;
  assign n17484 = n5417 | n17483 ;
  assign n17485 = ( ~n15184 & n17483 ) | ( ~n15184 & n17484 ) | ( n17483 & n17484 ) ;
  assign n17486 = n5418 | n17485 ;
  assign n17487 = ( ~n15195 & n17485 ) | ( ~n15195 & n17486 ) | ( n17485 & n17486 ) ;
  assign n17488 = x17 & ~n17487 ;
  assign n17489 = ( ~x17 & n17481 ) | ( ~x17 & n17487 ) | ( n17481 & n17487 ) ;
  assign n17490 = ( ~n17482 & n17488 ) | ( ~n17482 & n17489 ) | ( n17488 & n17489 ) ;
  assign n17491 = n5232 & n14352 ;
  assign n17492 = x20 & n17491 ;
  assign n17493 = n4874 & n13992 ;
  assign n17494 = n4878 | n17493 ;
  assign n17495 = ( n14520 & n17493 ) | ( n14520 & n17494 ) | ( n17493 & n17494 ) ;
  assign n17496 = n4879 | n17495 ;
  assign n17497 = ( n14531 & n17495 ) | ( n14531 & n17496 ) | ( n17495 & n17496 ) ;
  assign n17498 = x20 & ~n17497 ;
  assign n17499 = ( ~x20 & n17491 ) | ( ~x20 & n17497 ) | ( n17491 & n17497 ) ;
  assign n17500 = ( ~n17492 & n17498 ) | ( ~n17492 & n17499 ) | ( n17498 & n17499 ) ;
  assign n17501 = n4215 & ~n14007 ;
  assign n17502 = n4200 & n14002 ;
  assign n17503 = n2083 & ~n14004 ;
  assign n17504 = n17502 | n17503 ;
  assign n17505 = n17501 | n17504 ;
  assign n17506 = x26 & n17505 ;
  assign n17507 = n4203 & n14066 ;
  assign n17508 = ( ~x26 & n17505 ) | ( ~x26 & n17507 ) | ( n17505 & n17507 ) ;
  assign n17509 = x26 & ~n17507 ;
  assign n17510 = ( ~n17506 & n17508 ) | ( ~n17506 & n17509 ) | ( n17508 & n17509 ) ;
  assign n17511 = x26 & ~n17212 ;
  assign n17512 = ~n17428 & n17511 ;
  assign n17513 = n3500 & ~n14014 ;
  assign n17514 = ( n17510 & n17512 ) | ( n17510 & n17513 ) | ( n17512 & n17513 ) ;
  assign n17515 = ( ~n17510 & n17512 ) | ( ~n17510 & n17513 ) | ( n17512 & n17513 ) ;
  assign n17516 = ( n17510 & ~n17514 ) | ( n17510 & n17515 ) | ( ~n17514 & n17515 ) ;
  assign n17517 = n4591 & ~n14130 ;
  assign n17518 = x23 & n17517 ;
  assign n17519 = n4584 & ~n14000 ;
  assign n17520 = n4649 | n17519 ;
  assign n17521 = ( n13996 & n17519 ) | ( n13996 & n17520 ) | ( n17519 & n17520 ) ;
  assign n17522 = n4637 & n13998 ;
  assign n17523 = n17521 | n17522 ;
  assign n17524 = x23 & ~n17523 ;
  assign n17525 = ( ~x23 & n17517 ) | ( ~x23 & n17523 ) | ( n17517 & n17523 ) ;
  assign n17526 = ( ~n17518 & n17524 ) | ( ~n17518 & n17525 ) | ( n17524 & n17525 ) ;
  assign n17527 = ( ~n17433 & n17516 ) | ( ~n17433 & n17526 ) | ( n17516 & n17526 ) ;
  assign n17528 = ( n17433 & n17516 ) | ( n17433 & n17526 ) | ( n17516 & n17526 ) ;
  assign n17529 = ( n17433 & n17527 ) | ( n17433 & ~n17528 ) | ( n17527 & ~n17528 ) ;
  assign n17530 = ( ~n17435 & n17500 ) | ( ~n17435 & n17529 ) | ( n17500 & n17529 ) ;
  assign n17531 = ( n17435 & n17500 ) | ( n17435 & n17529 ) | ( n17500 & n17529 ) ;
  assign n17532 = ( n17435 & n17530 ) | ( n17435 & ~n17531 ) | ( n17530 & ~n17531 ) ;
  assign n17533 = ( ~n17439 & n17490 ) | ( ~n17439 & n17532 ) | ( n17490 & n17532 ) ;
  assign n17534 = ( n17439 & n17490 ) | ( n17439 & n17532 ) | ( n17490 & n17532 ) ;
  assign n17535 = ( n17439 & n17533 ) | ( n17439 & ~n17534 ) | ( n17533 & ~n17534 ) ;
  assign n17536 = ( ~n17442 & n17480 ) | ( ~n17442 & n17535 ) | ( n17480 & n17535 ) ;
  assign n17537 = ( n17442 & n17480 ) | ( n17442 & n17535 ) | ( n17480 & n17535 ) ;
  assign n17538 = ( n17442 & n17536 ) | ( n17442 & ~n17537 ) | ( n17536 & ~n17537 ) ;
  assign n17539 = ( ~n17445 & n17470 ) | ( ~n17445 & n17538 ) | ( n17470 & n17538 ) ;
  assign n17540 = ( n17445 & n17470 ) | ( n17445 & n17538 ) | ( n17470 & n17538 ) ;
  assign n17541 = ( n17445 & n17539 ) | ( n17445 & ~n17540 ) | ( n17539 & ~n17540 ) ;
  assign n17542 = ( ~n17448 & n17460 ) | ( ~n17448 & n17541 ) | ( n17460 & n17541 ) ;
  assign n17543 = ( n17448 & n17460 ) | ( n17448 & n17541 ) | ( n17460 & n17541 ) ;
  assign n17544 = ( n17448 & n17542 ) | ( n17448 & ~n17543 ) | ( n17542 & ~n17543 ) ;
  assign n17545 = n4874 & ~n13280 ;
  assign n17546 = n4878 | n17545 ;
  assign n17547 = ( n13475 & n17545 ) | ( n13475 & n17546 ) | ( n17545 & n17546 ) ;
  assign n17548 = n5232 & ~n13473 ;
  assign n17549 = n17547 | n17548 ;
  assign n17550 = x20 & n17549 ;
  assign n17551 = n4879 & n13671 ;
  assign n17552 = ( ~x20 & n17549 ) | ( ~x20 & n17551 ) | ( n17549 & n17551 ) ;
  assign n17553 = x20 & ~n17551 ;
  assign n17554 = ( ~n17550 & n17552 ) | ( ~n17550 & n17553 ) | ( n17552 & n17553 ) ;
  assign n17555 = n4584 & ~n10237 ;
  assign n17556 = n4649 | n17555 ;
  assign n17557 = ( ~n10235 & n17555 ) | ( ~n10235 & n17556 ) | ( n17555 & n17556 ) ;
  assign n17558 = n4637 & n10214 ;
  assign n17559 = n17557 | n17558 ;
  assign n17560 = x23 & n17559 ;
  assign n17561 = n4591 & n10371 ;
  assign n17562 = x23 & ~n17561 ;
  assign n17563 = ( ~x23 & n17559 ) | ( ~x23 & n17561 ) | ( n17559 & n17561 ) ;
  assign n17564 = ( ~n17560 & n17562 ) | ( ~n17560 & n17563 ) | ( n17562 & n17563 ) ;
  assign n17565 = n4215 & ~n10332 ;
  assign n17566 = n4200 & n10329 ;
  assign n17567 = n2083 & n10326 ;
  assign n17568 = n17566 | n17567 ;
  assign n17569 = n17565 | n17568 ;
  assign n17570 = x26 & n17569 ;
  assign n17571 = n4203 & ~n10383 ;
  assign n17572 = ( ~x26 & n17569 ) | ( ~x26 & n17571 ) | ( n17569 & n17571 ) ;
  assign n17573 = x26 & ~n17571 ;
  assign n17574 = ( ~n17570 & n17572 ) | ( ~n17570 & n17573 ) | ( n17572 & n17573 ) ;
  assign n17575 = n3501 & n10241 ;
  assign n17576 = x29 & n17575 ;
  assign n17577 = n3536 & n10243 ;
  assign n17578 = n4039 | n17577 ;
  assign n17579 = ( n10239 & n17577 ) | ( n10239 & n17578 ) | ( n17577 & n17578 ) ;
  assign n17580 = n3541 | n17579 ;
  assign n17581 = ( n12575 & n17579 ) | ( n12575 & n17580 ) | ( n17579 & n17580 ) ;
  assign n17582 = x29 & ~n17581 ;
  assign n17583 = ( ~x29 & n17575 ) | ( ~x29 & n17581 ) | ( n17575 & n17581 ) ;
  assign n17584 = ( ~n17576 & n17582 ) | ( ~n17576 & n17583 ) | ( n17582 & n17583 ) ;
  assign n17585 = n150 | n242 ;
  assign n17586 = n912 | n17585 ;
  assign n17587 = n3037 | n17586 ;
  assign n17588 = n1229 | n2288 ;
  assign n17589 = n17587 | n17588 ;
  assign n17590 = n627 | n896 ;
  assign n17591 = n1698 | n17590 ;
  assign n17592 = n1958 | n17591 ;
  assign n17593 = n17589 | n17592 ;
  assign n17594 = n434 | n712 ;
  assign n17595 = n554 | n17594 ;
  assign n17596 = n13404 | n17595 ;
  assign n17597 = n618 & ~n1069 ;
  assign n17598 = ~n270 & n17597 ;
  assign n17599 = ~n17596 & n17598 ;
  assign n17600 = n2357 | n2933 ;
  assign n17601 = n4384 | n5617 ;
  assign n17602 = n17600 | n17601 ;
  assign n17603 = n17599 & ~n17602 ;
  assign n17604 = ~n17593 & n17603 ;
  assign n17605 = ~n5124 & n17604 ;
  assign n17606 = ~n2797 & n17605 ;
  assign n17607 = ~n3903 & n17606 ;
  assign n17608 = ( n17319 & n17321 ) | ( n17319 & ~n17607 ) | ( n17321 & ~n17607 ) ;
  assign n17609 = ( ~n17085 & n17320 ) | ( ~n17085 & n17607 ) | ( n17320 & n17607 ) ;
  assign n17610 = ( ~n17319 & n17608 ) | ( ~n17319 & n17609 ) | ( n17608 & n17609 ) ;
  assign n17611 = n3274 & n10245 ;
  assign n17612 = n3273 & ~n10316 ;
  assign n17613 = n17611 | n17612 ;
  assign n17614 = n390 | n17613 ;
  assign n17615 = ( ~n10414 & n17613 ) | ( ~n10414 & n17614 ) | ( n17613 & n17614 ) ;
  assign n17616 = n3270 & ~n10320 ;
  assign n17617 = n17615 | n17616 ;
  assign n17618 = ( n17584 & ~n17610 ) | ( n17584 & n17617 ) | ( ~n17610 & n17617 ) ;
  assign n17619 = ( n17584 & n17610 ) | ( n17584 & ~n17617 ) | ( n17610 & ~n17617 ) ;
  assign n17620 = ( ~n17584 & n17618 ) | ( ~n17584 & n17619 ) | ( n17618 & n17619 ) ;
  assign n17621 = ( n17324 & n17574 ) | ( n17324 & ~n17620 ) | ( n17574 & ~n17620 ) ;
  assign n17622 = ( ~n17324 & n17574 ) | ( ~n17324 & n17620 ) | ( n17574 & n17620 ) ;
  assign n17623 = ( ~n17574 & n17621 ) | ( ~n17574 & n17622 ) | ( n17621 & n17622 ) ;
  assign n17624 = ( ~n17326 & n17564 ) | ( ~n17326 & n17623 ) | ( n17564 & n17623 ) ;
  assign n17625 = ( n17326 & n17564 ) | ( n17326 & ~n17623 ) | ( n17564 & ~n17623 ) ;
  assign n17626 = ( ~n17564 & n17624 ) | ( ~n17564 & n17625 ) | ( n17624 & n17625 ) ;
  assign n17627 = ( n17330 & n17554 ) | ( n17330 & ~n17626 ) | ( n17554 & ~n17626 ) ;
  assign n17628 = ( ~n17330 & n17554 ) | ( ~n17330 & n17626 ) | ( n17554 & n17626 ) ;
  assign n17629 = ( ~n17554 & n17627 ) | ( ~n17554 & n17628 ) | ( n17627 & n17628 ) ;
  assign n17630 = ( n17333 & n17336 ) | ( n17333 & ~n17629 ) | ( n17336 & ~n17629 ) ;
  assign n17631 = ( ~n17333 & n17336 ) | ( ~n17333 & n17629 ) | ( n17336 & n17629 ) ;
  assign n17632 = ( ~n17336 & n17630 ) | ( ~n17336 & n17631 ) | ( n17630 & n17631 ) ;
  assign n17633 = ( n17342 & n17345 ) | ( n17342 & ~n17632 ) | ( n17345 & ~n17632 ) ;
  assign n17634 = ( ~n17342 & n17345 ) | ( ~n17342 & n17632 ) | ( n17345 & n17632 ) ;
  assign n17635 = ( ~n17345 & n17633 ) | ( ~n17345 & n17634 ) | ( n17633 & n17634 ) ;
  assign n17636 = n40 & ~n17635 ;
  assign n17637 = n8721 & n17346 ;
  assign n17638 = n8340 & ~n17126 ;
  assign n17639 = n17637 | n17638 ;
  assign n17640 = n17636 | n17639 ;
  assign n17641 = x5 & n17640 ;
  assign n17642 = n17137 | n17346 ;
  assign n17643 = n17635 & ~n17642 ;
  assign n17644 = ~n17354 & n17635 ;
  assign n17645 = ( ~n17354 & n17635 ) | ( ~n17354 & n17642 ) | ( n17635 & n17642 ) ;
  assign n17646 = ( n17643 & ~n17644 ) | ( n17643 & n17645 ) | ( ~n17644 & n17645 ) ;
  assign n17647 = n8341 & ~n17646 ;
  assign n17648 = ( ~x5 & n17640 ) | ( ~x5 & n17647 ) | ( n17640 & n17647 ) ;
  assign n17649 = x5 & ~n17647 ;
  assign n17650 = ( ~n17641 & n17648 ) | ( ~n17641 & n17649 ) | ( n17648 & n17649 ) ;
  assign n17651 = ( n17450 & n17544 ) | ( n17450 & n17650 ) | ( n17544 & n17650 ) ;
  assign n17652 = n4215 & ~n10237 ;
  assign n17653 = n4200 & ~n10332 ;
  assign n17654 = n2083 & n10329 ;
  assign n17655 = n17653 | n17654 ;
  assign n17656 = n17652 | n17655 ;
  assign n17657 = x26 & n17656 ;
  assign n17658 = n4203 & n12756 ;
  assign n17659 = ( ~x26 & n17656 ) | ( ~x26 & n17658 ) | ( n17656 & n17658 ) ;
  assign n17660 = x26 & ~n17658 ;
  assign n17661 = ( ~n17657 & n17659 ) | ( ~n17657 & n17660 ) | ( n17659 & n17660 ) ;
  assign n17662 = n3501 & n10239 ;
  assign n17663 = x29 & n17662 ;
  assign n17664 = n3536 & n10241 ;
  assign n17665 = n4039 | n17664 ;
  assign n17666 = ( n10326 & n17664 ) | ( n10326 & n17665 ) | ( n17664 & n17665 ) ;
  assign n17667 = n3541 | n17666 ;
  assign n17668 = ( n12222 & n17666 ) | ( n12222 & n17667 ) | ( n17666 & n17667 ) ;
  assign n17669 = x29 & ~n17668 ;
  assign n17670 = ( ~x29 & n17662 ) | ( ~x29 & n17668 ) | ( n17662 & n17668 ) ;
  assign n17671 = ( ~n17663 & n17669 ) | ( ~n17663 & n17670 ) | ( n17669 & n17670 ) ;
  assign n17672 = n390 & ~n11989 ;
  assign n17673 = n3270 & n10243 ;
  assign n17674 = n3274 & ~n10320 ;
  assign n17675 = n3273 & n10245 ;
  assign n17676 = n17674 | n17675 ;
  assign n17677 = n17673 | n17676 ;
  assign n17678 = n17672 | n17677 ;
  assign n17679 = n2285 | n4341 ;
  assign n17680 = n339 | n524 ;
  assign n17681 = n17679 | n17680 ;
  assign n17682 = n1127 | n3729 ;
  assign n17683 = n276 | n471 ;
  assign n17684 = n629 | n17683 ;
  assign n17685 = n17682 | n17684 ;
  assign n17686 = n17681 | n17685 ;
  assign n17687 = n10164 | n17686 ;
  assign n17688 = n4802 | n17687 ;
  assign n17689 = n2867 | n15499 ;
  assign n17690 = n308 | n1302 ;
  assign n17691 = n756 | n17690 ;
  assign n17692 = n5479 | n17691 ;
  assign n17693 = n17689 | n17692 ;
  assign n17694 = n178 | n242 ;
  assign n17695 = n1573 | n17694 ;
  assign n17696 = n134 | n335 ;
  assign n17697 = n322 | n17696 ;
  assign n17698 = n17695 | n17697 ;
  assign n17699 = n5944 | n17698 ;
  assign n17700 = n17693 | n17699 ;
  assign n17701 = n3121 | n17700 ;
  assign n17702 = n17688 | n17701 ;
  assign n17703 = ( n17336 & n17607 ) | ( n17336 & ~n17702 ) | ( n17607 & ~n17702 ) ;
  assign n17704 = ( n17336 & ~n17607 ) | ( n17336 & n17702 ) | ( ~n17607 & n17702 ) ;
  assign n17705 = ( ~n17336 & n17703 ) | ( ~n17336 & n17704 ) | ( n17703 & n17704 ) ;
  assign n17706 = ( ~n17609 & n17678 ) | ( ~n17609 & n17705 ) | ( n17678 & n17705 ) ;
  assign n17707 = ( n17609 & n17678 ) | ( n17609 & n17705 ) | ( n17678 & n17705 ) ;
  assign n17708 = ( n17609 & n17706 ) | ( n17609 & ~n17707 ) | ( n17706 & ~n17707 ) ;
  assign n17709 = ( n17618 & ~n17671 ) | ( n17618 & n17708 ) | ( ~n17671 & n17708 ) ;
  assign n17710 = ( n17618 & n17671 ) | ( n17618 & n17708 ) | ( n17671 & n17708 ) ;
  assign n17711 = ( n17671 & n17709 ) | ( n17671 & ~n17710 ) | ( n17709 & ~n17710 ) ;
  assign n17712 = ( ~n17621 & n17661 ) | ( ~n17621 & n17711 ) | ( n17661 & n17711 ) ;
  assign n17713 = ( n17621 & n17661 ) | ( n17621 & n17711 ) | ( n17661 & n17711 ) ;
  assign n17714 = ( n17621 & n17712 ) | ( n17621 & ~n17713 ) | ( n17712 & ~n17713 ) ;
  assign n17715 = n4637 & ~n10235 ;
  assign n17716 = x23 & n17715 ;
  assign n17717 = n4584 & n10214 ;
  assign n17718 = n4649 | n17717 ;
  assign n17719 = ( ~n13280 & n17717 ) | ( ~n13280 & n17718 ) | ( n17717 & n17718 ) ;
  assign n17720 = n4591 | n17719 ;
  assign n17721 = ( ~n13285 & n17719 ) | ( ~n13285 & n17720 ) | ( n17719 & n17720 ) ;
  assign n17722 = x23 & ~n17721 ;
  assign n17723 = ( ~x23 & n17715 ) | ( ~x23 & n17721 ) | ( n17715 & n17721 ) ;
  assign n17724 = ( ~n17716 & n17722 ) | ( ~n17716 & n17723 ) | ( n17722 & n17723 ) ;
  assign n17725 = ( ~n17625 & n17714 ) | ( ~n17625 & n17724 ) | ( n17714 & n17724 ) ;
  assign n17726 = ( n17625 & n17714 ) | ( n17625 & n17724 ) | ( n17714 & n17724 ) ;
  assign n17727 = ( n17625 & n17725 ) | ( n17625 & ~n17726 ) | ( n17725 & ~n17726 ) ;
  assign n17728 = n4874 | n4878 ;
  assign n17729 = ( n4878 & ~n13473 ) | ( n4878 & n17728 ) | ( ~n13473 & n17728 ) ;
  assign n17730 = n5232 | n17729 ;
  assign n17731 = ( n13475 & n17729 ) | ( n13475 & n17730 ) | ( n17729 & n17730 ) ;
  assign n17732 = x20 & n17731 ;
  assign n17733 = n4875 & n13477 ;
  assign n17734 = x20 & ~n17733 ;
  assign n17735 = ( ~x20 & n17731 ) | ( ~x20 & n17733 ) | ( n17731 & n17733 ) ;
  assign n17736 = ( ~n17732 & n17734 ) | ( ~n17732 & n17735 ) | ( n17734 & n17735 ) ;
  assign n17737 = ( n17627 & n17727 ) | ( n17627 & n17736 ) | ( n17727 & n17736 ) ;
  assign n17738 = ( ~n17627 & n17727 ) | ( ~n17627 & n17736 ) | ( n17727 & n17736 ) ;
  assign n17739 = ( n17627 & ~n17737 ) | ( n17627 & n17738 ) | ( ~n17737 & n17738 ) ;
  assign n17740 = ( n17630 & ~n17633 ) | ( n17630 & n17739 ) | ( ~n17633 & n17739 ) ;
  assign n17741 = ( n17630 & n17633 ) | ( n17630 & n17739 ) | ( n17633 & n17739 ) ;
  assign n17742 = ( n17633 & n17740 ) | ( n17633 & ~n17741 ) | ( n17740 & ~n17741 ) ;
  assign n17743 = n40 & n17742 ;
  assign n17744 = x5 & n17743 ;
  assign n17745 = n17644 & n17742 ;
  assign n17746 = ~n17635 & n17642 ;
  assign n17747 = ( n17644 & ~n17742 ) | ( n17644 & n17746 ) | ( ~n17742 & n17746 ) ;
  assign n17748 = n17742 & ~n17746 ;
  assign n17749 = ( ~n17745 & n17747 ) | ( ~n17745 & n17748 ) | ( n17747 & n17748 ) ;
  assign n17750 = n8721 & ~n17635 ;
  assign n17751 = n8340 & n17346 ;
  assign n17752 = n17750 | n17751 ;
  assign n17753 = n8341 | n17752 ;
  assign n17754 = ( ~n17749 & n17752 ) | ( ~n17749 & n17753 ) | ( n17752 & n17753 ) ;
  assign n17755 = x5 & ~n17754 ;
  assign n17756 = ( ~x5 & n17743 ) | ( ~x5 & n17754 ) | ( n17743 & n17754 ) ;
  assign n17757 = ( ~n17744 & n17755 ) | ( ~n17744 & n17756 ) | ( n17755 & n17756 ) ;
  assign n17758 = n7346 & ~n17139 ;
  assign n17759 = x8 & n17758 ;
  assign n17760 = n7341 & n16724 ;
  assign n17761 = n7345 | n17760 ;
  assign n17762 = ( ~n17126 & n17760 ) | ( ~n17126 & n17761 ) | ( n17760 & n17761 ) ;
  assign n17763 = n7644 & n16925 ;
  assign n17764 = n17762 | n17763 ;
  assign n17765 = x8 & ~n17764 ;
  assign n17766 = ( ~x8 & n17758 ) | ( ~x8 & n17764 ) | ( n17758 & n17764 ) ;
  assign n17767 = ( ~n17759 & n17765 ) | ( ~n17759 & n17766 ) | ( n17765 & n17766 ) ;
  assign n17768 = n6796 & ~n16338 ;
  assign n17769 = x11 & n17768 ;
  assign n17770 = n6567 & ~n16150 ;
  assign n17771 = n6570 | n17770 ;
  assign n17772 = ( ~n16531 & n17770 ) | ( ~n16531 & n17771 ) | ( n17770 & n17771 ) ;
  assign n17773 = n6571 | n17772 ;
  assign n17774 = ( ~n16542 & n17772 ) | ( ~n16542 & n17773 ) | ( n17772 & n17773 ) ;
  assign n17775 = x11 & ~n17774 ;
  assign n17776 = ( ~x11 & n17768 ) | ( ~x11 & n17774 ) | ( n17768 & n17774 ) ;
  assign n17777 = ( ~n17769 & n17775 ) | ( ~n17769 & n17776 ) | ( n17775 & n17776 ) ;
  assign n17778 = n5915 & ~n15965 ;
  assign n17779 = x14 & n17778 ;
  assign n17780 = n5909 & n15561 ;
  assign n17781 = n5914 | n17780 ;
  assign n17782 = ( ~n15954 & n17780 ) | ( ~n15954 & n17781 ) | ( n17780 & n17781 ) ;
  assign n17783 = n6332 & ~n15806 ;
  assign n17784 = n17782 | n17783 ;
  assign n17785 = x14 & ~n17784 ;
  assign n17786 = ( ~x14 & n17778 ) | ( ~x14 & n17784 ) | ( n17778 & n17784 ) ;
  assign n17787 = ( ~n17779 & n17785 ) | ( ~n17779 & n17786 ) | ( n17785 & n17786 ) ;
  assign n17788 = n5584 & ~n15184 ;
  assign n17789 = x17 & n17788 ;
  assign n17790 = n5413 & n14942 ;
  assign n17791 = n5417 | n17790 ;
  assign n17792 = ( ~n15394 & n17790 ) | ( ~n15394 & n17791 ) | ( n17790 & n17791 ) ;
  assign n17793 = n5418 | n17792 ;
  assign n17794 = ( n15405 & n17792 ) | ( n15405 & n17793 ) | ( n17792 & n17793 ) ;
  assign n17795 = x17 & ~n17794 ;
  assign n17796 = ( ~x17 & n17788 ) | ( ~x17 & n17794 ) | ( n17788 & n17794 ) ;
  assign n17797 = ( ~n17789 & n17795 ) | ( ~n17789 & n17796 ) | ( n17795 & n17796 ) ;
  assign n17798 = n4879 & ~n14734 ;
  assign n17799 = x20 & n17798 ;
  assign n17800 = n4874 & n14352 ;
  assign n17801 = n4878 | n17800 ;
  assign n17802 = ( ~n14723 & n17800 ) | ( ~n14723 & n17801 ) | ( n17800 & n17801 ) ;
  assign n17803 = n5232 & n14520 ;
  assign n17804 = n17802 | n17803 ;
  assign n17805 = x20 & ~n17804 ;
  assign n17806 = ( ~x20 & n17798 ) | ( ~x20 & n17804 ) | ( n17798 & n17804 ) ;
  assign n17807 = ( ~n17799 & n17805 ) | ( ~n17799 & n17806 ) | ( n17805 & n17806 ) ;
  assign n17808 = n4649 & n13992 ;
  assign n17809 = x23 & n17808 ;
  assign n17810 = n4637 & n13996 ;
  assign n17811 = n4584 & n13998 ;
  assign n17812 = n17810 | n17811 ;
  assign n17813 = n4591 | n17812 ;
  assign n17814 = ( n14024 & n17812 ) | ( n14024 & n17813 ) | ( n17812 & n17813 ) ;
  assign n17815 = x23 & ~n17814 ;
  assign n17816 = ( ~x23 & n17808 ) | ( ~x23 & n17814 ) | ( n17808 & n17814 ) ;
  assign n17817 = ( ~n17809 & n17815 ) | ( ~n17809 & n17816 ) | ( n17815 & n17816 ) ;
  assign n17818 = n4215 & ~n14000 ;
  assign n17819 = n4200 & ~n14007 ;
  assign n17820 = n2083 & n14002 ;
  assign n17821 = n17819 | n17820 ;
  assign n17822 = n17818 | n17821 ;
  assign n17823 = x26 & n17822 ;
  assign n17824 = n4203 & ~n14042 ;
  assign n17825 = ( ~x26 & n17822 ) | ( ~x26 & n17824 ) | ( n17822 & n17824 ) ;
  assign n17826 = x26 & ~n17824 ;
  assign n17827 = ( ~n17823 & n17825 ) | ( ~n17823 & n17826 ) | ( n17825 & n17826 ) ;
  assign n17828 = n4039 & ~n14004 ;
  assign n17829 = ( n3501 & n6605 ) | ( n3501 & n14004 ) | ( n6605 & n14004 ) ;
  assign n17830 = ~n14014 & n17829 ;
  assign n17831 = n17828 | n17830 ;
  assign n17832 = n3500 & n14015 ;
  assign n17833 = n17831 | n17832 ;
  assign n17834 = n17513 | n17833 ;
  assign n17835 = ( x29 & n17513 ) | ( x29 & ~n17833 ) | ( n17513 & ~n17833 ) ;
  assign n17836 = x29 & ~n17831 ;
  assign n17837 = ( n17834 & ~n17835 ) | ( n17834 & n17836 ) | ( ~n17835 & n17836 ) ;
  assign n17838 = n17510 & n17514 ;
  assign n17839 = ( n17827 & n17837 ) | ( n17827 & n17838 ) | ( n17837 & n17838 ) ;
  assign n17840 = ( ~n17827 & n17837 ) | ( ~n17827 & n17838 ) | ( n17837 & n17838 ) ;
  assign n17841 = ( n17827 & ~n17839 ) | ( n17827 & n17840 ) | ( ~n17839 & n17840 ) ;
  assign n17842 = ( ~n17528 & n17817 ) | ( ~n17528 & n17841 ) | ( n17817 & n17841 ) ;
  assign n17843 = ( n17528 & n17817 ) | ( n17528 & n17841 ) | ( n17817 & n17841 ) ;
  assign n17844 = ( n17528 & n17842 ) | ( n17528 & ~n17843 ) | ( n17842 & ~n17843 ) ;
  assign n17845 = ( ~n17531 & n17807 ) | ( ~n17531 & n17844 ) | ( n17807 & n17844 ) ;
  assign n17846 = ( n17531 & n17807 ) | ( n17531 & n17844 ) | ( n17807 & n17844 ) ;
  assign n17847 = ( n17531 & n17845 ) | ( n17531 & ~n17846 ) | ( n17845 & ~n17846 ) ;
  assign n17848 = ( n17534 & n17797 ) | ( n17534 & n17847 ) | ( n17797 & n17847 ) ;
  assign n17849 = ( ~n17534 & n17797 ) | ( ~n17534 & n17847 ) | ( n17797 & n17847 ) ;
  assign n17850 = ( n17534 & ~n17848 ) | ( n17534 & n17849 ) | ( ~n17848 & n17849 ) ;
  assign n17851 = ( ~n17537 & n17787 ) | ( ~n17537 & n17850 ) | ( n17787 & n17850 ) ;
  assign n17852 = ( n17537 & n17787 ) | ( n17537 & n17850 ) | ( n17787 & n17850 ) ;
  assign n17853 = ( n17537 & n17851 ) | ( n17537 & ~n17852 ) | ( n17851 & ~n17852 ) ;
  assign n17854 = ( ~n17540 & n17777 ) | ( ~n17540 & n17853 ) | ( n17777 & n17853 ) ;
  assign n17855 = ( n17540 & n17777 ) | ( n17540 & n17853 ) | ( n17777 & n17853 ) ;
  assign n17856 = ( n17540 & n17854 ) | ( n17540 & ~n17855 ) | ( n17854 & ~n17855 ) ;
  assign n17857 = ( ~n17543 & n17767 ) | ( ~n17543 & n17856 ) | ( n17767 & n17856 ) ;
  assign n17858 = ( n17543 & n17767 ) | ( n17543 & n17856 ) | ( n17767 & n17856 ) ;
  assign n17859 = ( n17543 & n17857 ) | ( n17543 & ~n17858 ) | ( n17857 & ~n17858 ) ;
  assign n17860 = ( n17651 & n17757 ) | ( n17651 & n17859 ) | ( n17757 & n17859 ) ;
  assign n17861 = ( x17 & ~x18 ) | ( x17 & x19 ) | ( ~x18 & x19 ) ;
  assign n17862 = ( x18 & ~x20 ) | ( x18 & n17861 ) | ( ~x20 & n17861 ) ;
  assign n17863 = ~n4870 & n17862 ;
  assign n17864 = ( n13475 & n17862 ) | ( n13475 & n17863 ) | ( n17862 & n17863 ) ;
  assign n17865 = n4873 & ~n13475 ;
  assign n17866 = n17864 | n17865 ;
  assign n17867 = n4637 & ~n13280 ;
  assign n17868 = x23 & n17867 ;
  assign n17869 = n4649 & ~n13473 ;
  assign n17870 = n4584 & ~n10235 ;
  assign n17871 = n17869 | n17870 ;
  assign n17872 = n4591 | n17871 ;
  assign n17873 = ( ~n13480 & n17871 ) | ( ~n13480 & n17872 ) | ( n17871 & n17872 ) ;
  assign n17874 = x23 & ~n17873 ;
  assign n17875 = ( ~x23 & n17867 ) | ( ~x23 & n17873 ) | ( n17867 & n17873 ) ;
  assign n17876 = ( ~n17868 & n17874 ) | ( ~n17868 & n17875 ) | ( n17874 & n17875 ) ;
  assign n17877 = n4215 & n10214 ;
  assign n17878 = n4200 & ~n10237 ;
  assign n17879 = n2083 & ~n10332 ;
  assign n17880 = n17878 | n17879 ;
  assign n17881 = n17877 | n17880 ;
  assign n17882 = x26 & n17881 ;
  assign n17883 = n4203 & n12953 ;
  assign n17884 = ( ~x26 & n17881 ) | ( ~x26 & n17883 ) | ( n17881 & n17883 ) ;
  assign n17885 = x26 & ~n17883 ;
  assign n17886 = ( ~n17882 & n17884 ) | ( ~n17882 & n17885 ) | ( n17884 & n17885 ) ;
  assign n17887 = n3501 & n10326 ;
  assign n17888 = x29 & n17887 ;
  assign n17889 = n3536 & n10239 ;
  assign n17890 = n4039 | n17889 ;
  assign n17891 = ( n10329 & n17889 ) | ( n10329 & n17890 ) | ( n17889 & n17890 ) ;
  assign n17892 = n3541 | n17891 ;
  assign n17893 = ( n10397 & n17891 ) | ( n10397 & n17892 ) | ( n17891 & n17892 ) ;
  assign n17894 = x29 & ~n17893 ;
  assign n17895 = ( ~x29 & n17887 ) | ( ~x29 & n17893 ) | ( n17887 & n17893 ) ;
  assign n17896 = ( ~n17888 & n17894 ) | ( ~n17888 & n17895 ) | ( n17894 & n17895 ) ;
  assign n17897 = n3273 & ~n10320 ;
  assign n17898 = n3270 | n17897 ;
  assign n17899 = ( n10241 & n17897 ) | ( n10241 & n17898 ) | ( n17897 & n17898 ) ;
  assign n17900 = n390 | n17899 ;
  assign n17901 = ( n12105 & n17899 ) | ( n12105 & n17900 ) | ( n17899 & n17900 ) ;
  assign n17902 = n3274 & n10243 ;
  assign n17903 = n17901 | n17902 ;
  assign n17904 = n2690 | n6160 ;
  assign n17905 = n2321 | n3546 ;
  assign n17906 = n17904 | n17905 ;
  assign n17907 = n188 | n968 ;
  assign n17908 = n4279 | n17907 ;
  assign n17909 = n17906 | n17908 ;
  assign n17910 = n220 | n419 ;
  assign n17911 = n2544 | n17910 ;
  assign n17912 = n2399 | n17911 ;
  assign n17913 = n1048 | n17912 ;
  assign n17914 = n1285 | n2293 ;
  assign n17915 = n2851 | n17914 ;
  assign n17916 = n17913 | n17915 ;
  assign n17917 = n17909 | n17916 ;
  assign n17918 = n1388 | n4894 ;
  assign n17919 = n17917 | n17918 ;
  assign n17920 = n494 | n916 ;
  assign n17921 = n2890 | n17920 ;
  assign n17922 = n4382 | n17921 ;
  assign n17923 = n189 | n987 ;
  assign n17924 = n17922 | n17923 ;
  assign n17925 = n1391 | n1872 ;
  assign n17926 = n262 | n17925 ;
  assign n17927 = n17924 | n17926 ;
  assign n17928 = n526 | n794 ;
  assign n17929 = n360 | n17928 ;
  assign n17930 = n200 | n17929 ;
  assign n17931 = ~n556 & n618 ;
  assign n17932 = ~n83 & n17931 ;
  assign n17933 = ~n17930 & n17932 ;
  assign n17934 = ~n17927 & n17933 ;
  assign n17935 = n432 | n2744 ;
  assign n17936 = n378 | n487 ;
  assign n17937 = n17935 | n17936 ;
  assign n17938 = n184 | n207 ;
  assign n17939 = n518 | n17938 ;
  assign n17940 = n17937 | n17939 ;
  assign n17941 = n1135 | n17940 ;
  assign n17942 = n17686 | n17941 ;
  assign n17943 = n17934 & ~n17942 ;
  assign n17944 = ~n17919 & n17943 ;
  assign n17945 = ~n3122 & n17944 ;
  assign n17946 = ( ~n17703 & n17903 ) | ( ~n17703 & n17945 ) | ( n17903 & n17945 ) ;
  assign n17947 = ( n17703 & n17903 ) | ( n17703 & ~n17945 ) | ( n17903 & ~n17945 ) ;
  assign n17948 = ( ~n17903 & n17946 ) | ( ~n17903 & n17947 ) | ( n17946 & n17947 ) ;
  assign n17949 = ( n17707 & n17896 ) | ( n17707 & ~n17948 ) | ( n17896 & ~n17948 ) ;
  assign n17950 = ( ~n17707 & n17896 ) | ( ~n17707 & n17948 ) | ( n17896 & n17948 ) ;
  assign n17951 = ( ~n17896 & n17949 ) | ( ~n17896 & n17950 ) | ( n17949 & n17950 ) ;
  assign n17952 = ( ~n17710 & n17886 ) | ( ~n17710 & n17951 ) | ( n17886 & n17951 ) ;
  assign n17953 = ( n17710 & n17886 ) | ( n17710 & ~n17951 ) | ( n17886 & ~n17951 ) ;
  assign n17954 = ( ~n17886 & n17952 ) | ( ~n17886 & n17953 ) | ( n17952 & n17953 ) ;
  assign n17955 = ( n17713 & ~n17876 ) | ( n17713 & n17954 ) | ( ~n17876 & n17954 ) ;
  assign n17956 = ( n17713 & n17876 ) | ( n17713 & ~n17954 ) | ( n17876 & ~n17954 ) ;
  assign n17957 = ( ~n17713 & n17955 ) | ( ~n17713 & n17956 ) | ( n17955 & n17956 ) ;
  assign n17958 = ( ~n17726 & n17866 ) | ( ~n17726 & n17957 ) | ( n17866 & n17957 ) ;
  assign n17959 = ( n17726 & n17866 ) | ( n17726 & ~n17957 ) | ( n17866 & ~n17957 ) ;
  assign n17960 = ( ~n17866 & n17958 ) | ( ~n17866 & n17959 ) | ( n17958 & n17959 ) ;
  assign n17961 = ( ~n17737 & n17741 ) | ( ~n17737 & n17960 ) | ( n17741 & n17960 ) ;
  assign n17962 = ( n17737 & n17741 ) | ( n17737 & ~n17960 ) | ( n17741 & ~n17960 ) ;
  assign n17963 = ( ~n17741 & n17961 ) | ( ~n17741 & n17962 ) | ( n17961 & n17962 ) ;
  assign n17964 = n40 & ~n17963 ;
  assign n17965 = n8721 & n17742 ;
  assign n17966 = n8340 & ~n17635 ;
  assign n17967 = n17965 | n17966 ;
  assign n17968 = n17964 | n17967 ;
  assign n17969 = x5 & n17968 ;
  assign n17970 = n17742 | n17746 ;
  assign n17971 = ~n17644 & n17742 ;
  assign n17972 = n17963 & ~n17971 ;
  assign n17973 = n17970 & n17972 ;
  assign n17974 = ~n17963 & n17970 ;
  assign n17975 = ( ~n17742 & n17745 ) | ( ~n17742 & n17974 ) | ( n17745 & n17974 ) ;
  assign n17976 = ( n17963 & ~n17973 ) | ( n17963 & n17975 ) | ( ~n17973 & n17975 ) ;
  assign n17977 = n8341 & ~n17976 ;
  assign n17978 = ( ~x5 & n17968 ) | ( ~x5 & n17977 ) | ( n17968 & n17977 ) ;
  assign n17979 = x5 & ~n17977 ;
  assign n17980 = ( ~n17969 & n17978 ) | ( ~n17969 & n17979 ) | ( n17978 & n17979 ) ;
  assign n17981 = n7644 & ~n17126 ;
  assign n17982 = x8 & n17981 ;
  assign n17983 = n7341 & n16925 ;
  assign n17984 = n7345 | n17983 ;
  assign n17985 = ( n17346 & n17983 ) | ( n17346 & n17984 ) | ( n17983 & n17984 ) ;
  assign n17986 = n7346 | n17985 ;
  assign n17987 = ( ~n17356 & n17985 ) | ( ~n17356 & n17986 ) | ( n17985 & n17986 ) ;
  assign n17988 = x8 & ~n17987 ;
  assign n17989 = ( ~x8 & n17981 ) | ( ~x8 & n17987 ) | ( n17981 & n17987 ) ;
  assign n17990 = ( ~n17982 & n17988 ) | ( ~n17982 & n17989 ) | ( n17988 & n17989 ) ;
  assign n17991 = n6796 & ~n16531 ;
  assign n17992 = x11 & n17991 ;
  assign n17993 = n6567 & ~n16338 ;
  assign n17994 = n6570 | n17993 ;
  assign n17995 = ( n16724 & n17993 ) | ( n16724 & n17994 ) | ( n17993 & n17994 ) ;
  assign n17996 = n6571 | n17995 ;
  assign n17997 = ( n16735 & n17995 ) | ( n16735 & n17996 ) | ( n17995 & n17996 ) ;
  assign n17998 = x11 & ~n17997 ;
  assign n17999 = ( ~x11 & n17991 ) | ( ~x11 & n17997 ) | ( n17991 & n17997 ) ;
  assign n18000 = ( ~n17992 & n17998 ) | ( ~n17992 & n17999 ) | ( n17998 & n17999 ) ;
  assign n18001 = n5584 & ~n15394 ;
  assign n18002 = x17 & n18001 ;
  assign n18003 = n5413 & ~n15184 ;
  assign n18004 = n5417 | n18003 ;
  assign n18005 = ( n15561 & n18003 ) | ( n15561 & n18004 ) | ( n18003 & n18004 ) ;
  assign n18006 = n5418 | n18005 ;
  assign n18007 = ( n15573 & n18005 ) | ( n15573 & n18006 ) | ( n18005 & n18006 ) ;
  assign n18008 = x17 & ~n18007 ;
  assign n18009 = ( ~x17 & n18001 ) | ( ~x17 & n18007 ) | ( n18001 & n18007 ) ;
  assign n18010 = ( ~n18002 & n18008 ) | ( ~n18002 & n18009 ) | ( n18008 & n18009 ) ;
  assign n18011 = n5232 & ~n14723 ;
  assign n18012 = x20 & n18011 ;
  assign n18013 = n4874 & n14520 ;
  assign n18014 = n4878 | n18013 ;
  assign n18015 = ( n14942 & n18013 ) | ( n14942 & n18014 ) | ( n18013 & n18014 ) ;
  assign n18016 = n4879 | n18015 ;
  assign n18017 = ( ~n14953 & n18015 ) | ( ~n14953 & n18016 ) | ( n18015 & n18016 ) ;
  assign n18018 = x20 & ~n18017 ;
  assign n18019 = ( ~x20 & n18011 ) | ( ~x20 & n18017 ) | ( n18011 & n18017 ) ;
  assign n18020 = ( ~n18012 & n18018 ) | ( ~n18012 & n18019 ) | ( n18018 & n18019 ) ;
  assign n18021 = n4637 & n13992 ;
  assign n18022 = x23 & n18021 ;
  assign n18023 = n4584 & n13996 ;
  assign n18024 = n4649 | n18023 ;
  assign n18025 = ( n14352 & n18023 ) | ( n14352 & n18024 ) | ( n18023 & n18024 ) ;
  assign n18026 = n4591 | n18025 ;
  assign n18027 = ( n14363 & n18025 ) | ( n14363 & n18026 ) | ( n18025 & n18026 ) ;
  assign n18028 = x23 & ~n18027 ;
  assign n18029 = ( ~x23 & n18021 ) | ( ~x23 & n18027 ) | ( n18021 & n18027 ) ;
  assign n18030 = ( ~n18022 & n18028 ) | ( ~n18022 & n18029 ) | ( n18028 & n18029 ) ;
  assign n18031 = n3501 & ~n14004 ;
  assign n18032 = n3536 & ~n14014 ;
  assign n18033 = n18031 | n18032 ;
  assign n18034 = n3541 | n18033 ;
  assign n18035 = ( n14072 & n18033 ) | ( n14072 & n18034 ) | ( n18033 & n18034 ) ;
  assign n18036 = n4039 & n14002 ;
  assign n18037 = n18035 | n18036 ;
  assign n18038 = ~x29 & n18037 ;
  assign n18039 = ( x29 & n17834 ) | ( x29 & n18037 ) | ( n17834 & n18037 ) ;
  assign n18040 = n17834 & n18037 ;
  assign n18041 = ( n18038 & n18039 ) | ( n18038 & ~n18040 ) | ( n18039 & ~n18040 ) ;
  assign n18042 = n4215 & n13998 ;
  assign n18043 = n4200 & ~n14000 ;
  assign n18044 = n2083 & ~n14007 ;
  assign n18045 = n18043 | n18044 ;
  assign n18046 = n18042 | n18045 ;
  assign n18047 = x26 & n18046 ;
  assign n18048 = n4203 & n14115 ;
  assign n18049 = ( ~x26 & n18046 ) | ( ~x26 & n18048 ) | ( n18046 & n18048 ) ;
  assign n18050 = x26 & ~n18048 ;
  assign n18051 = ( ~n18047 & n18049 ) | ( ~n18047 & n18050 ) | ( n18049 & n18050 ) ;
  assign n18052 = ( ~n17839 & n18041 ) | ( ~n17839 & n18051 ) | ( n18041 & n18051 ) ;
  assign n18053 = ( n17839 & n18041 ) | ( n17839 & n18051 ) | ( n18041 & n18051 ) ;
  assign n18054 = ( n17839 & n18052 ) | ( n17839 & ~n18053 ) | ( n18052 & ~n18053 ) ;
  assign n18055 = ( ~n17843 & n18030 ) | ( ~n17843 & n18054 ) | ( n18030 & n18054 ) ;
  assign n18056 = ( n17843 & n18030 ) | ( n17843 & n18054 ) | ( n18030 & n18054 ) ;
  assign n18057 = ( n17843 & n18055 ) | ( n17843 & ~n18056 ) | ( n18055 & ~n18056 ) ;
  assign n18058 = ( ~n17846 & n18020 ) | ( ~n17846 & n18057 ) | ( n18020 & n18057 ) ;
  assign n18059 = ( n17846 & n18020 ) | ( n17846 & n18057 ) | ( n18020 & n18057 ) ;
  assign n18060 = ( n17846 & n18058 ) | ( n17846 & ~n18059 ) | ( n18058 & ~n18059 ) ;
  assign n18061 = ( ~n17848 & n18010 ) | ( ~n17848 & n18060 ) | ( n18010 & n18060 ) ;
  assign n18062 = ( n17848 & n18010 ) | ( n17848 & n18060 ) | ( n18010 & n18060 ) ;
  assign n18063 = ( n17848 & n18061 ) | ( n17848 & ~n18062 ) | ( n18061 & ~n18062 ) ;
  assign n18064 = n5915 & ~n16161 ;
  assign n18065 = x14 & n18064 ;
  assign n18066 = n5914 & ~n16150 ;
  assign n18067 = n6332 & ~n15954 ;
  assign n18068 = n5909 & ~n15806 ;
  assign n18069 = n18067 | n18068 ;
  assign n18070 = n18066 | n18069 ;
  assign n18071 = x14 & ~n18070 ;
  assign n18072 = ( ~x14 & n18064 ) | ( ~x14 & n18070 ) | ( n18064 & n18070 ) ;
  assign n18073 = ( ~n18065 & n18071 ) | ( ~n18065 & n18072 ) | ( n18071 & n18072 ) ;
  assign n18074 = ( ~n17852 & n18063 ) | ( ~n17852 & n18073 ) | ( n18063 & n18073 ) ;
  assign n18075 = ( n17852 & n18063 ) | ( n17852 & n18073 ) | ( n18063 & n18073 ) ;
  assign n18076 = ( n17852 & n18074 ) | ( n17852 & ~n18075 ) | ( n18074 & ~n18075 ) ;
  assign n18077 = ( ~n17855 & n18000 ) | ( ~n17855 & n18076 ) | ( n18000 & n18076 ) ;
  assign n18078 = ( n17855 & n18000 ) | ( n17855 & n18076 ) | ( n18000 & n18076 ) ;
  assign n18079 = ( n17855 & n18077 ) | ( n17855 & ~n18078 ) | ( n18077 & ~n18078 ) ;
  assign n18080 = ( n17858 & n17990 ) | ( n17858 & n18079 ) | ( n17990 & n18079 ) ;
  assign n18081 = ( ~n17858 & n17990 ) | ( ~n17858 & n18079 ) | ( n17990 & n18079 ) ;
  assign n18082 = ( n17858 & ~n18080 ) | ( n17858 & n18081 ) | ( ~n18080 & n18081 ) ;
  assign n18083 = ( n17860 & n17980 ) | ( n17860 & n18082 ) | ( n17980 & n18082 ) ;
  assign n18084 = n5915 & ~n16349 ;
  assign n18085 = x14 & n18084 ;
  assign n18086 = n5909 & ~n15954 ;
  assign n18087 = n5914 | n18086 ;
  assign n18088 = ( ~n16338 & n18086 ) | ( ~n16338 & n18087 ) | ( n18086 & n18087 ) ;
  assign n18089 = n6332 & ~n16150 ;
  assign n18090 = n18088 | n18089 ;
  assign n18091 = x14 & ~n18090 ;
  assign n18092 = ( ~x14 & n18084 ) | ( ~x14 & n18090 ) | ( n18084 & n18090 ) ;
  assign n18093 = ( ~n18085 & n18091 ) | ( ~n18085 & n18092 ) | ( n18091 & n18092 ) ;
  assign n18094 = n5584 & n15561 ;
  assign n18095 = x17 & n18094 ;
  assign n18096 = n5413 & ~n15394 ;
  assign n18097 = n5417 | n18096 ;
  assign n18098 = ( ~n15806 & n18096 ) | ( ~n15806 & n18097 ) | ( n18096 & n18097 ) ;
  assign n18099 = n5418 | n18098 ;
  assign n18100 = ( n15817 & n18098 ) | ( n15817 & n18099 ) | ( n18098 & n18099 ) ;
  assign n18101 = x17 & ~n18100 ;
  assign n18102 = ( ~x17 & n18094 ) | ( ~x17 & n18100 ) | ( n18094 & n18100 ) ;
  assign n18103 = ( ~n18095 & n18101 ) | ( ~n18095 & n18102 ) | ( n18101 & n18102 ) ;
  assign n18104 = n5232 & n14942 ;
  assign n18105 = x20 & n18104 ;
  assign n18106 = n4874 & ~n14723 ;
  assign n18107 = n4878 | n18106 ;
  assign n18108 = ( ~n15184 & n18106 ) | ( ~n15184 & n18107 ) | ( n18106 & n18107 ) ;
  assign n18109 = n4879 | n18108 ;
  assign n18110 = ( ~n15195 & n18108 ) | ( ~n15195 & n18109 ) | ( n18108 & n18109 ) ;
  assign n18111 = x20 & ~n18110 ;
  assign n18112 = ( ~x20 & n18104 ) | ( ~x20 & n18110 ) | ( n18104 & n18110 ) ;
  assign n18113 = ( ~n18105 & n18111 ) | ( ~n18105 & n18112 ) | ( n18111 & n18112 ) ;
  assign n18114 = n4649 & n14520 ;
  assign n18115 = n4591 | n18114 ;
  assign n18116 = ( n14531 & n18114 ) | ( n14531 & n18115 ) | ( n18114 & n18115 ) ;
  assign n18117 = n4584 & n13992 ;
  assign n18118 = ( ~x23 & n18116 ) | ( ~x23 & n18117 ) | ( n18116 & n18117 ) ;
  assign n18119 = n4637 & n14352 ;
  assign n18120 = x23 & ~n18117 ;
  assign n18121 = n18119 | n18120 ;
  assign n18122 = ( n18116 & n18119 ) | ( n18116 & n18120 ) | ( n18119 & n18120 ) ;
  assign n18123 = ( n18118 & n18121 ) | ( n18118 & ~n18122 ) | ( n18121 & ~n18122 ) ;
  assign n18124 = x29 & n18039 ;
  assign n18125 = ~n18038 & n18124 ;
  assign n18126 = n389 & ~n14014 ;
  assign n18127 = n3541 & n14066 ;
  assign n18128 = n4039 & ~n14007 ;
  assign n18129 = n3501 & n14002 ;
  assign n18130 = n3536 & ~n14004 ;
  assign n18131 = n18129 | n18130 ;
  assign n18132 = n18128 | n18131 ;
  assign n18133 = n18127 | n18132 ;
  assign n18134 = ( n18125 & ~n18126 ) | ( n18125 & n18133 ) | ( ~n18126 & n18133 ) ;
  assign n18135 = ( n18125 & n18126 ) | ( n18125 & ~n18133 ) | ( n18126 & ~n18133 ) ;
  assign n18136 = ( ~n18125 & n18134 ) | ( ~n18125 & n18135 ) | ( n18134 & n18135 ) ;
  assign n18137 = n4215 & n13996 ;
  assign n18138 = n4200 & n13998 ;
  assign n18139 = n2083 & ~n14000 ;
  assign n18140 = n18138 | n18139 ;
  assign n18141 = n18137 | n18140 ;
  assign n18142 = x26 & n18141 ;
  assign n18143 = n4203 & ~n14130 ;
  assign n18144 = ( ~x26 & n18141 ) | ( ~x26 & n18143 ) | ( n18141 & n18143 ) ;
  assign n18145 = x26 & ~n18143 ;
  assign n18146 = ( ~n18142 & n18144 ) | ( ~n18142 & n18145 ) | ( n18144 & n18145 ) ;
  assign n18147 = ( ~n18053 & n18136 ) | ( ~n18053 & n18146 ) | ( n18136 & n18146 ) ;
  assign n18148 = ( n18053 & n18136 ) | ( n18053 & n18146 ) | ( n18136 & n18146 ) ;
  assign n18149 = ( n18053 & n18147 ) | ( n18053 & ~n18148 ) | ( n18147 & ~n18148 ) ;
  assign n18150 = ( ~n18056 & n18123 ) | ( ~n18056 & n18149 ) | ( n18123 & n18149 ) ;
  assign n18151 = ( n18056 & n18123 ) | ( n18056 & n18149 ) | ( n18123 & n18149 ) ;
  assign n18152 = ( n18056 & n18150 ) | ( n18056 & ~n18151 ) | ( n18150 & ~n18151 ) ;
  assign n18153 = ( ~n18059 & n18113 ) | ( ~n18059 & n18152 ) | ( n18113 & n18152 ) ;
  assign n18154 = ( n18059 & n18113 ) | ( n18059 & n18152 ) | ( n18113 & n18152 ) ;
  assign n18155 = ( n18059 & n18153 ) | ( n18059 & ~n18154 ) | ( n18153 & ~n18154 ) ;
  assign n18156 = ( ~n18062 & n18103 ) | ( ~n18062 & n18155 ) | ( n18103 & n18155 ) ;
  assign n18157 = ( n18062 & n18103 ) | ( n18062 & n18155 ) | ( n18103 & n18155 ) ;
  assign n18158 = ( n18062 & n18156 ) | ( n18062 & ~n18157 ) | ( n18156 & ~n18157 ) ;
  assign n18159 = ( ~n18075 & n18093 ) | ( ~n18075 & n18158 ) | ( n18093 & n18158 ) ;
  assign n18160 = ( n18075 & n18093 ) | ( n18075 & n18158 ) | ( n18093 & n18158 ) ;
  assign n18161 = ( n18075 & n18159 ) | ( n18075 & ~n18160 ) | ( n18159 & ~n18160 ) ;
  assign n18162 = n6796 & n16724 ;
  assign n18163 = x11 & n18162 ;
  assign n18164 = n6567 & ~n16531 ;
  assign n18165 = n6570 | n18164 ;
  assign n18166 = ( n16925 & n18164 ) | ( n16925 & n18165 ) | ( n18164 & n18165 ) ;
  assign n18167 = n6571 | n18166 ;
  assign n18168 = ( ~n16936 & n18166 ) | ( ~n16936 & n18167 ) | ( n18166 & n18167 ) ;
  assign n18169 = x11 & ~n18168 ;
  assign n18170 = ( ~x11 & n18162 ) | ( ~x11 & n18168 ) | ( n18162 & n18168 ) ;
  assign n18171 = ( ~n18163 & n18169 ) | ( ~n18163 & n18170 ) | ( n18169 & n18170 ) ;
  assign n18172 = ( ~n18078 & n18161 ) | ( ~n18078 & n18171 ) | ( n18161 & n18171 ) ;
  assign n18173 = ( n18078 & n18161 ) | ( n18078 & n18171 ) | ( n18161 & n18171 ) ;
  assign n18174 = ( n18078 & n18172 ) | ( n18078 & ~n18173 ) | ( n18172 & ~n18173 ) ;
  assign n18175 = n7644 & n17346 ;
  assign n18176 = x8 & n18175 ;
  assign n18177 = n7341 & ~n17126 ;
  assign n18178 = n7345 | n18177 ;
  assign n18179 = ( ~n17635 & n18177 ) | ( ~n17635 & n18178 ) | ( n18177 & n18178 ) ;
  assign n18180 = n7346 | n18179 ;
  assign n18181 = ( ~n17646 & n18179 ) | ( ~n17646 & n18180 ) | ( n18179 & n18180 ) ;
  assign n18182 = x8 & ~n18181 ;
  assign n18183 = ( ~x8 & n18175 ) | ( ~x8 & n18181 ) | ( n18175 & n18181 ) ;
  assign n18184 = ( ~n18176 & n18182 ) | ( ~n18176 & n18183 ) | ( n18182 & n18183 ) ;
  assign n18185 = ( ~n18080 & n18174 ) | ( ~n18080 & n18184 ) | ( n18174 & n18184 ) ;
  assign n18186 = ( n18080 & n18174 ) | ( n18080 & n18184 ) | ( n18174 & n18184 ) ;
  assign n18187 = ( n18080 & n18185 ) | ( n18080 & ~n18186 ) | ( n18185 & ~n18186 ) ;
  assign n18188 = n4584 & ~n13280 ;
  assign n18189 = n4649 | n18188 ;
  assign n18190 = ( n13475 & n18188 ) | ( n13475 & n18189 ) | ( n18188 & n18189 ) ;
  assign n18191 = n4637 & ~n13473 ;
  assign n18192 = n18190 | n18191 ;
  assign n18193 = x23 & n18192 ;
  assign n18194 = n4591 & n13671 ;
  assign n18195 = ( ~x23 & n18192 ) | ( ~x23 & n18194 ) | ( n18192 & n18194 ) ;
  assign n18196 = x23 & ~n18194 ;
  assign n18197 = ( ~n18193 & n18195 ) | ( ~n18193 & n18196 ) | ( n18195 & n18196 ) ;
  assign n18198 = n4203 & n10371 ;
  assign n18199 = n4215 & ~n10235 ;
  assign n18200 = n4200 & n10214 ;
  assign n18201 = n2083 & ~n10237 ;
  assign n18202 = n18200 | n18201 ;
  assign n18203 = n18199 | n18202 ;
  assign n18204 = n18198 | n18203 ;
  assign n18205 = n3541 & ~n10383 ;
  assign n18206 = n4039 & ~n10332 ;
  assign n18207 = n3501 & n10329 ;
  assign n18208 = n3536 & n10326 ;
  assign n18209 = n18207 | n18208 ;
  assign n18210 = n18206 | n18209 ;
  assign n18211 = n18205 | n18210 ;
  assign n18212 = n6269 & ~n18211 ;
  assign n18213 = ~n6269 & n18211 ;
  assign n18214 = n18212 | n18213 ;
  assign n18215 = n3273 & n10243 ;
  assign n18216 = n3270 | n18215 ;
  assign n18217 = ( n10239 & n18215 ) | ( n10239 & n18216 ) | ( n18215 & n18216 ) ;
  assign n18218 = n390 | n18217 ;
  assign n18219 = ( n12575 & n18217 ) | ( n12575 & n18218 ) | ( n18217 & n18218 ) ;
  assign n18220 = n3274 & n10241 ;
  assign n18221 = n18219 | n18220 ;
  assign n18222 = n2982 | n3384 ;
  assign n18223 = n173 | n558 ;
  assign n18224 = n18222 | n18223 ;
  assign n18225 = n148 | n279 ;
  assign n18226 = n695 | n18225 ;
  assign n18227 = n237 | n407 ;
  assign n18228 = n18226 | n18227 ;
  assign n18229 = n18224 | n18228 ;
  assign n18230 = n456 | n16108 ;
  assign n18231 = n1877 | n18230 ;
  assign n18232 = n18229 | n18231 ;
  assign n18233 = n1228 | n1665 ;
  assign n18234 = n3937 | n4967 ;
  assign n18235 = n18233 | n18234 ;
  assign n18236 = n1815 | n18235 ;
  assign n18237 = n18232 | n18236 ;
  assign n18238 = n2436 | n18237 ;
  assign n18239 = n5030 & ~n18238 ;
  assign n18240 = ~n14669 & n18239 ;
  assign n18241 = ( n17945 & n18221 ) | ( n17945 & ~n18240 ) | ( n18221 & ~n18240 ) ;
  assign n18242 = ( n17945 & ~n18221 ) | ( n17945 & n18240 ) | ( ~n18221 & n18240 ) ;
  assign n18243 = ( ~n17945 & n18241 ) | ( ~n17945 & n18242 ) | ( n18241 & n18242 ) ;
  assign n18244 = ( ~n17946 & n17949 ) | ( ~n17946 & n18243 ) | ( n17949 & n18243 ) ;
  assign n18245 = ( n17946 & n17949 ) | ( n17946 & ~n18243 ) | ( n17949 & ~n18243 ) ;
  assign n18246 = ( ~n17949 & n18244 ) | ( ~n17949 & n18245 ) | ( n18244 & n18245 ) ;
  assign n18247 = ( n18204 & ~n18214 ) | ( n18204 & n18246 ) | ( ~n18214 & n18246 ) ;
  assign n18248 = ( n18204 & n18214 ) | ( n18204 & ~n18246 ) | ( n18214 & ~n18246 ) ;
  assign n18249 = ( ~n18204 & n18247 ) | ( ~n18204 & n18248 ) | ( n18247 & n18248 ) ;
  assign n18250 = ( ~n17953 & n18197 ) | ( ~n17953 & n18249 ) | ( n18197 & n18249 ) ;
  assign n18251 = ( n17953 & n18197 ) | ( n17953 & ~n18249 ) | ( n18197 & ~n18249 ) ;
  assign n18252 = ( ~n18197 & n18250 ) | ( ~n18197 & n18251 ) | ( n18250 & n18251 ) ;
  assign n18253 = ( n17862 & n17956 ) | ( n17862 & ~n18252 ) | ( n17956 & ~n18252 ) ;
  assign n18254 = ( ~n17862 & n17956 ) | ( ~n17862 & n18252 ) | ( n17956 & n18252 ) ;
  assign n18255 = ( ~n17956 & n18253 ) | ( ~n17956 & n18254 ) | ( n18253 & n18254 ) ;
  assign n18256 = ( n17959 & n17962 ) | ( n17959 & ~n18255 ) | ( n17962 & ~n18255 ) ;
  assign n18257 = ( ~n17959 & n17962 ) | ( ~n17959 & n18255 ) | ( n17962 & n18255 ) ;
  assign n18258 = ( ~n17962 & n18256 ) | ( ~n17962 & n18257 ) | ( n18256 & n18257 ) ;
  assign n18259 = n40 & ~n18258 ;
  assign n18260 = n8721 & ~n17963 ;
  assign n18261 = n8340 & n17742 ;
  assign n18262 = n18260 | n18261 ;
  assign n18263 = n18259 | n18262 ;
  assign n18264 = x5 & n18263 ;
  assign n18265 = n17974 & ~n18258 ;
  assign n18266 = n17972 | n18258 ;
  assign n18267 = ( n17972 & n17974 ) | ( n17972 & n18258 ) | ( n17974 & n18258 ) ;
  assign n18268 = ( n18265 & n18266 ) | ( n18265 & ~n18267 ) | ( n18266 & ~n18267 ) ;
  assign n18269 = n8341 & n18268 ;
  assign n18270 = ( ~x5 & n18263 ) | ( ~x5 & n18269 ) | ( n18263 & n18269 ) ;
  assign n18271 = x5 & ~n18269 ;
  assign n18272 = ( ~n18264 & n18270 ) | ( ~n18264 & n18271 ) | ( n18270 & n18271 ) ;
  assign n18273 = ( n18083 & n18187 ) | ( n18083 & n18272 ) | ( n18187 & n18272 ) ;
  assign n18274 = n4584 | n4649 ;
  assign n18275 = ( n4649 & ~n13473 ) | ( n4649 & n18274 ) | ( ~n13473 & n18274 ) ;
  assign n18276 = n4637 | n18275 ;
  assign n18277 = ( n13475 & n18275 ) | ( n13475 & n18276 ) | ( n18275 & n18276 ) ;
  assign n18278 = x23 & n18277 ;
  assign n18279 = n4590 & n13477 ;
  assign n18280 = x23 & ~n18279 ;
  assign n18281 = ( ~x23 & n18277 ) | ( ~x23 & n18279 ) | ( n18277 & n18279 ) ;
  assign n18282 = ( ~n18278 & n18280 ) | ( ~n18278 & n18281 ) | ( n18280 & n18281 ) ;
  assign n18283 = x26 & ~n18204 ;
  assign n18284 = ~x26 & n18204 ;
  assign n18285 = n18283 | n18284 ;
  assign n18286 = x29 & ~n18211 ;
  assign n18287 = ~x29 & n18211 ;
  assign n18288 = n18286 | n18287 ;
  assign n18289 = ( ~n18246 & n18285 ) | ( ~n18246 & n18288 ) | ( n18285 & n18288 ) ;
  assign n18290 = n4203 & ~n13285 ;
  assign n18291 = x26 & n18290 ;
  assign n18292 = n4215 & ~n13280 ;
  assign n18293 = n4200 & ~n10235 ;
  assign n18294 = n2083 & n10214 ;
  assign n18295 = n18293 | n18294 ;
  assign n18296 = n18292 | n18295 ;
  assign n18297 = x26 & ~n18296 ;
  assign n18298 = ( ~x26 & n18290 ) | ( ~x26 & n18296 ) | ( n18290 & n18296 ) ;
  assign n18299 = ( ~n18291 & n18297 ) | ( ~n18291 & n18298 ) | ( n18297 & n18298 ) ;
  assign n18300 = n4039 & ~n10237 ;
  assign n18301 = n3501 & ~n10332 ;
  assign n18302 = n3536 & n10329 ;
  assign n18303 = n18301 | n18302 ;
  assign n18304 = n18300 | n18303 ;
  assign n18305 = x29 & n18304 ;
  assign n18306 = n3541 & n12756 ;
  assign n18307 = ( ~x29 & n18304 ) | ( ~x29 & n18306 ) | ( n18304 & n18306 ) ;
  assign n18308 = x29 & ~n18306 ;
  assign n18309 = ( ~n18305 & n18307 ) | ( ~n18305 & n18308 ) | ( n18307 & n18308 ) ;
  assign n18310 = n3273 & n10241 ;
  assign n18311 = n3270 | n18310 ;
  assign n18312 = ( n10326 & n18310 ) | ( n10326 & n18311 ) | ( n18310 & n18311 ) ;
  assign n18313 = n390 | n18312 ;
  assign n18314 = ( n12222 & n18312 ) | ( n12222 & n18313 ) | ( n18312 & n18313 ) ;
  assign n18315 = n3274 & n10239 ;
  assign n18316 = n18314 | n18315 ;
  assign n18317 = n1339 | n1401 ;
  assign n18318 = n2935 | n3928 ;
  assign n18319 = n18317 | n18318 ;
  assign n18320 = n1065 | n1365 ;
  assign n18321 = n305 | n912 ;
  assign n18322 = n18320 | n18321 ;
  assign n18323 = n488 | n1006 ;
  assign n18324 = n624 | n18323 ;
  assign n18325 = n1130 | n18324 ;
  assign n18326 = n18322 | n18325 ;
  assign n18327 = n18319 | n18326 ;
  assign n18328 = n1684 | n18327 ;
  assign n18329 = n3178 | n18328 ;
  assign n18330 = n2221 & ~n18329 ;
  assign n18331 = n497 | n1196 ;
  assign n18332 = n347 | n379 ;
  assign n18333 = n2381 | n18332 ;
  assign n18334 = n18331 | n18333 ;
  assign n18335 = n44 & n231 ;
  assign n18336 = n18334 | n18335 ;
  assign n18337 = n1137 | n2516 ;
  assign n18338 = n17300 | n18337 ;
  assign n18339 = n672 | n18338 ;
  assign n18340 = n18336 | n18339 ;
  assign n18341 = n1157 | n3112 ;
  assign n18342 = n1938 | n18341 ;
  assign n18343 = n18340 | n18342 ;
  assign n18344 = n18330 & ~n18343 ;
  assign n18345 = ( n17862 & ~n17945 ) | ( n17862 & n18344 ) | ( ~n17945 & n18344 ) ;
  assign n18346 = ( n17862 & n17945 ) | ( n17862 & n18344 ) | ( n17945 & n18344 ) ;
  assign n18347 = ( n17945 & n18345 ) | ( n17945 & ~n18346 ) | ( n18345 & ~n18346 ) ;
  assign n18348 = ( n18241 & n18316 ) | ( n18241 & ~n18347 ) | ( n18316 & ~n18347 ) ;
  assign n18349 = ( ~n18241 & n18316 ) | ( ~n18241 & n18347 ) | ( n18316 & n18347 ) ;
  assign n18350 = ( ~n18316 & n18348 ) | ( ~n18316 & n18349 ) | ( n18348 & n18349 ) ;
  assign n18351 = ( n18245 & n18309 ) | ( n18245 & ~n18350 ) | ( n18309 & ~n18350 ) ;
  assign n18352 = ( ~n18245 & n18309 ) | ( ~n18245 & n18350 ) | ( n18309 & n18350 ) ;
  assign n18353 = ( ~n18309 & n18351 ) | ( ~n18309 & n18352 ) | ( n18351 & n18352 ) ;
  assign n18354 = ( n18289 & n18299 ) | ( n18289 & ~n18353 ) | ( n18299 & ~n18353 ) ;
  assign n18355 = ( n18289 & ~n18299 ) | ( n18289 & n18353 ) | ( ~n18299 & n18353 ) ;
  assign n18356 = ( ~n18289 & n18354 ) | ( ~n18289 & n18355 ) | ( n18354 & n18355 ) ;
  assign n18357 = ( n18251 & n18282 ) | ( n18251 & ~n18356 ) | ( n18282 & ~n18356 ) ;
  assign n18358 = ( n18251 & ~n18282 ) | ( n18251 & n18356 ) | ( ~n18282 & n18356 ) ;
  assign n18359 = ( ~n18251 & n18357 ) | ( ~n18251 & n18358 ) | ( n18357 & n18358 ) ;
  assign n18360 = ( n18253 & n18256 ) | ( n18253 & ~n18359 ) | ( n18256 & ~n18359 ) ;
  assign n18361 = ( ~n18253 & n18256 ) | ( ~n18253 & n18359 ) | ( n18256 & n18359 ) ;
  assign n18362 = ( ~n18256 & n18360 ) | ( ~n18256 & n18361 ) | ( n18360 & n18361 ) ;
  assign n18363 = n40 & ~n18362 ;
  assign n18364 = n8721 & ~n18258 ;
  assign n18365 = n8340 & ~n17963 ;
  assign n18366 = n18364 | n18365 ;
  assign n18367 = n18363 | n18366 ;
  assign n18368 = x5 & n18367 ;
  assign n18369 = ~n18266 & n18362 ;
  assign n18370 = ~n17974 & n18258 ;
  assign n18371 = ( n18266 & n18362 ) | ( n18266 & ~n18370 ) | ( n18362 & ~n18370 ) ;
  assign n18372 = n18362 & ~n18370 ;
  assign n18373 = ( n18369 & n18371 ) | ( n18369 & ~n18372 ) | ( n18371 & ~n18372 ) ;
  assign n18374 = n8341 & ~n18373 ;
  assign n18375 = ( ~x5 & n18367 ) | ( ~x5 & n18374 ) | ( n18367 & n18374 ) ;
  assign n18376 = x5 & ~n18374 ;
  assign n18377 = ( ~n18368 & n18375 ) | ( ~n18368 & n18376 ) | ( n18375 & n18376 ) ;
  assign n18378 = n7345 & n17742 ;
  assign n18379 = x8 & n18378 ;
  assign n18380 = n7644 & ~n17635 ;
  assign n18381 = n7341 & n17346 ;
  assign n18382 = n18380 | n18381 ;
  assign n18383 = n7346 | n18382 ;
  assign n18384 = ( ~n17749 & n18382 ) | ( ~n17749 & n18383 ) | ( n18382 & n18383 ) ;
  assign n18385 = x8 & ~n18384 ;
  assign n18386 = ( ~x8 & n18378 ) | ( ~x8 & n18384 ) | ( n18378 & n18384 ) ;
  assign n18387 = ( ~n18379 & n18385 ) | ( ~n18379 & n18386 ) | ( n18385 & n18386 ) ;
  assign n18388 = n6796 & n16925 ;
  assign n18389 = x11 & n18388 ;
  assign n18390 = n6567 & n16724 ;
  assign n18391 = n6570 | n18390 ;
  assign n18392 = ( ~n17126 & n18390 ) | ( ~n17126 & n18391 ) | ( n18390 & n18391 ) ;
  assign n18393 = n6571 | n18392 ;
  assign n18394 = ( ~n17139 & n18392 ) | ( ~n17139 & n18393 ) | ( n18392 & n18393 ) ;
  assign n18395 = x11 & ~n18394 ;
  assign n18396 = ( ~x11 & n18388 ) | ( ~x11 & n18394 ) | ( n18388 & n18394 ) ;
  assign n18397 = ( ~n18389 & n18395 ) | ( ~n18389 & n18396 ) | ( n18395 & n18396 ) ;
  assign n18398 = n6332 & ~n16338 ;
  assign n18399 = x14 & n18398 ;
  assign n18400 = n5909 & ~n16150 ;
  assign n18401 = n5914 | n18400 ;
  assign n18402 = ( ~n16531 & n18400 ) | ( ~n16531 & n18401 ) | ( n18400 & n18401 ) ;
  assign n18403 = n5915 | n18402 ;
  assign n18404 = ( ~n16542 & n18402 ) | ( ~n16542 & n18403 ) | ( n18402 & n18403 ) ;
  assign n18405 = x14 & ~n18404 ;
  assign n18406 = ( ~x14 & n18398 ) | ( ~x14 & n18404 ) | ( n18398 & n18404 ) ;
  assign n18407 = ( ~n18399 & n18405 ) | ( ~n18399 & n18406 ) | ( n18405 & n18406 ) ;
  assign n18408 = n5584 & ~n15806 ;
  assign n18409 = x17 & n18408 ;
  assign n18410 = n5413 & n15561 ;
  assign n18411 = n5417 | n18410 ;
  assign n18412 = ( ~n15954 & n18410 ) | ( ~n15954 & n18411 ) | ( n18410 & n18411 ) ;
  assign n18413 = n5418 | n18412 ;
  assign n18414 = ( ~n15965 & n18412 ) | ( ~n15965 & n18413 ) | ( n18412 & n18413 ) ;
  assign n18415 = x17 & ~n18414 ;
  assign n18416 = ( ~x17 & n18408 ) | ( ~x17 & n18414 ) | ( n18408 & n18414 ) ;
  assign n18417 = ( ~n18409 & n18415 ) | ( ~n18409 & n18416 ) | ( n18415 & n18416 ) ;
  assign n18418 = n5232 & ~n15184 ;
  assign n18419 = x20 & n18418 ;
  assign n18420 = n4874 & n14942 ;
  assign n18421 = n4878 | n18420 ;
  assign n18422 = ( ~n15394 & n18420 ) | ( ~n15394 & n18421 ) | ( n18420 & n18421 ) ;
  assign n18423 = n4879 | n18422 ;
  assign n18424 = ( n15405 & n18422 ) | ( n15405 & n18423 ) | ( n18422 & n18423 ) ;
  assign n18425 = x20 & ~n18424 ;
  assign n18426 = ( ~x20 & n18418 ) | ( ~x20 & n18424 ) | ( n18418 & n18424 ) ;
  assign n18427 = ( ~n18419 & n18425 ) | ( ~n18419 & n18426 ) | ( n18425 & n18426 ) ;
  assign n18428 = n4591 & ~n14734 ;
  assign n18429 = x23 & n18428 ;
  assign n18430 = n4584 & n14352 ;
  assign n18431 = n4649 | n18430 ;
  assign n18432 = ( ~n14723 & n18430 ) | ( ~n14723 & n18431 ) | ( n18430 & n18431 ) ;
  assign n18433 = n4637 & n14520 ;
  assign n18434 = n18432 | n18433 ;
  assign n18435 = x23 & ~n18434 ;
  assign n18436 = ( ~x23 & n18428 ) | ( ~x23 & n18434 ) | ( n18428 & n18434 ) ;
  assign n18437 = ( ~n18429 & n18435 ) | ( ~n18429 & n18436 ) | ( n18435 & n18436 ) ;
  assign n18438 = n4215 & n13992 ;
  assign n18439 = x26 & n18438 ;
  assign n18440 = n4200 & n13996 ;
  assign n18441 = n2083 & n13998 ;
  assign n18442 = n18440 | n18441 ;
  assign n18443 = n4203 | n18442 ;
  assign n18444 = ( n14024 & n18442 ) | ( n14024 & n18443 ) | ( n18442 & n18443 ) ;
  assign n18445 = x26 & ~n18444 ;
  assign n18446 = ( ~x26 & n18438 ) | ( ~x26 & n18444 ) | ( n18438 & n18444 ) ;
  assign n18447 = ( ~n18439 & n18445 ) | ( ~n18439 & n18446 ) | ( n18445 & n18446 ) ;
  assign n18448 = n3501 & ~n14007 ;
  assign n18449 = x29 & n18448 ;
  assign n18450 = n3536 & n14002 ;
  assign n18451 = n4039 | n18450 ;
  assign n18452 = ( ~n14000 & n18450 ) | ( ~n14000 & n18451 ) | ( n18450 & n18451 ) ;
  assign n18453 = n3541 | n18452 ;
  assign n18454 = ( ~n14042 & n18452 ) | ( ~n14042 & n18453 ) | ( n18452 & n18453 ) ;
  assign n18455 = x29 & ~n18454 ;
  assign n18456 = ( ~x29 & n18448 ) | ( ~x29 & n18454 ) | ( n18448 & n18454 ) ;
  assign n18457 = ( ~n18449 & n18455 ) | ( ~n18449 & n18456 ) | ( n18455 & n18456 ) ;
  assign n18458 = n389 & n14015 ;
  assign n18459 = ( x29 & x30 ) | ( x29 & ~n14004 ) | ( x30 & ~n14004 ) ;
  assign n18460 = ( x31 & ~n14014 ) | ( x31 & n18459 ) | ( ~n14014 & n18459 ) ;
  assign n18461 = x31 & n18459 ;
  assign n18462 = ( n18458 & n18460 ) | ( n18458 & ~n18461 ) | ( n18460 & ~n18461 ) ;
  assign n18463 = n835 | n1151 ;
  assign n18464 = n278 | n953 ;
  assign n18465 = n2103 | n18464 ;
  assign n18466 = n18463 | n18465 ;
  assign n18467 = n328 | n528 ;
  assign n18468 = n131 | n18467 ;
  assign n18469 = n1868 | n18468 ;
  assign n18470 = n18466 | n18469 ;
  assign n18471 = n975 | n1542 ;
  assign n18472 = n18470 | n18471 ;
  assign n18473 = n865 | n1720 ;
  assign n18474 = n243 | n3508 ;
  assign n18475 = n1816 | n18474 ;
  assign n18476 = n18473 | n18475 ;
  assign n18477 = n2590 | n13221 ;
  assign n18478 = n18476 | n18477 ;
  assign n18479 = n1737 | n3285 ;
  assign n18480 = n3909 | n18479 ;
  assign n18481 = n1629 | n18480 ;
  assign n18482 = n18478 | n18481 ;
  assign n18483 = n18472 | n18482 ;
  assign n18484 = n983 | n1005 ;
  assign n18485 = n4262 | n18484 ;
  assign n18486 = n257 | n794 ;
  assign n18487 = n82 | n18486 ;
  assign n18488 = n1399 | n18487 ;
  assign n18489 = n18485 | n18488 ;
  assign n18490 = n416 | n3791 ;
  assign n18491 = n16897 | n18490 ;
  assign n18492 = ~n1333 & n3161 ;
  assign n18493 = ~n18491 & n18492 ;
  assign n18494 = ~n18489 & n18493 ;
  assign n18495 = n1767 | n1963 ;
  assign n18496 = n3946 | n18495 ;
  assign n18497 = n18494 & ~n18496 ;
  assign n18498 = ~n18483 & n18497 ;
  assign n18499 = ~n13613 & n18498 ;
  assign n18500 = ~n18462 & n18499 ;
  assign n18501 = n18462 & ~n18499 ;
  assign n18502 = n18500 | n18501 ;
  assign n18503 = x29 & ~n18133 ;
  assign n18504 = ( x29 & n18133 ) | ( x29 & n18134 ) | ( n18133 & n18134 ) ;
  assign n18505 = ( n18133 & n18503 ) | ( n18133 & ~n18504 ) | ( n18503 & ~n18504 ) ;
  assign n18506 = ( n18457 & ~n18502 ) | ( n18457 & n18505 ) | ( ~n18502 & n18505 ) ;
  assign n18507 = ( n18457 & n18502 ) | ( n18457 & ~n18505 ) | ( n18502 & ~n18505 ) ;
  assign n18508 = ( ~n18457 & n18506 ) | ( ~n18457 & n18507 ) | ( n18506 & n18507 ) ;
  assign n18509 = ( n18148 & ~n18447 ) | ( n18148 & n18508 ) | ( ~n18447 & n18508 ) ;
  assign n18510 = ( n18148 & n18447 ) | ( n18148 & ~n18508 ) | ( n18447 & ~n18508 ) ;
  assign n18511 = ( ~n18148 & n18509 ) | ( ~n18148 & n18510 ) | ( n18509 & n18510 ) ;
  assign n18512 = ( n18151 & n18437 ) | ( n18151 & ~n18511 ) | ( n18437 & ~n18511 ) ;
  assign n18513 = ( n18151 & ~n18437 ) | ( n18151 & n18511 ) | ( ~n18437 & n18511 ) ;
  assign n18514 = ( ~n18151 & n18512 ) | ( ~n18151 & n18513 ) | ( n18512 & n18513 ) ;
  assign n18515 = ( n18154 & n18427 ) | ( n18154 & ~n18514 ) | ( n18427 & ~n18514 ) ;
  assign n18516 = ( n18154 & ~n18427 ) | ( n18154 & n18514 ) | ( ~n18427 & n18514 ) ;
  assign n18517 = ( ~n18154 & n18515 ) | ( ~n18154 & n18516 ) | ( n18515 & n18516 ) ;
  assign n18518 = ( n18157 & n18417 ) | ( n18157 & ~n18517 ) | ( n18417 & ~n18517 ) ;
  assign n18519 = ( n18157 & ~n18417 ) | ( n18157 & n18517 ) | ( ~n18417 & n18517 ) ;
  assign n18520 = ( ~n18157 & n18518 ) | ( ~n18157 & n18519 ) | ( n18518 & n18519 ) ;
  assign n18521 = ( n18160 & ~n18407 ) | ( n18160 & n18520 ) | ( ~n18407 & n18520 ) ;
  assign n18522 = ( n18160 & n18407 ) | ( n18160 & ~n18520 ) | ( n18407 & ~n18520 ) ;
  assign n18523 = ( ~n18160 & n18521 ) | ( ~n18160 & n18522 ) | ( n18521 & n18522 ) ;
  assign n18524 = ( n18173 & n18397 ) | ( n18173 & ~n18523 ) | ( n18397 & ~n18523 ) ;
  assign n18525 = ( n18173 & ~n18397 ) | ( n18173 & n18523 ) | ( ~n18397 & n18523 ) ;
  assign n18526 = ( ~n18173 & n18524 ) | ( ~n18173 & n18525 ) | ( n18524 & n18525 ) ;
  assign n18527 = ( n18186 & n18387 ) | ( n18186 & ~n18526 ) | ( n18387 & ~n18526 ) ;
  assign n18528 = ( n18186 & ~n18387 ) | ( n18186 & n18526 ) | ( ~n18387 & n18526 ) ;
  assign n18529 = ( ~n18186 & n18527 ) | ( ~n18186 & n18528 ) | ( n18527 & n18528 ) ;
  assign n18530 = ( n18273 & n18377 ) | ( n18273 & ~n18529 ) | ( n18377 & ~n18529 ) ;
  assign n18531 = n6796 & ~n17126 ;
  assign n18532 = x11 & n18531 ;
  assign n18533 = n6567 & n16925 ;
  assign n18534 = n6570 | n18533 ;
  assign n18535 = ( n17346 & n18533 ) | ( n17346 & n18534 ) | ( n18533 & n18534 ) ;
  assign n18536 = n6571 | n18535 ;
  assign n18537 = ( ~n17356 & n18535 ) | ( ~n17356 & n18536 ) | ( n18535 & n18536 ) ;
  assign n18538 = x11 & ~n18537 ;
  assign n18539 = ( ~x11 & n18531 ) | ( ~x11 & n18537 ) | ( n18531 & n18537 ) ;
  assign n18540 = ( ~n18532 & n18538 ) | ( ~n18532 & n18539 ) | ( n18538 & n18539 ) ;
  assign n18541 = n5418 & ~n16161 ;
  assign n18542 = x17 & n18541 ;
  assign n18543 = n5413 & ~n15806 ;
  assign n18544 = n5417 | n18543 ;
  assign n18545 = ( ~n16150 & n18543 ) | ( ~n16150 & n18544 ) | ( n18543 & n18544 ) ;
  assign n18546 = n5584 & ~n15954 ;
  assign n18547 = n18545 | n18546 ;
  assign n18548 = x17 & ~n18547 ;
  assign n18549 = ( ~x17 & n18541 ) | ( ~x17 & n18547 ) | ( n18541 & n18547 ) ;
  assign n18550 = ( ~n18542 & n18548 ) | ( ~n18542 & n18549 ) | ( n18548 & n18549 ) ;
  assign n18551 = n5232 & ~n15394 ;
  assign n18552 = x20 & n18551 ;
  assign n18553 = n4874 & ~n15184 ;
  assign n18554 = n4878 | n18553 ;
  assign n18555 = ( n15561 & n18553 ) | ( n15561 & n18554 ) | ( n18553 & n18554 ) ;
  assign n18556 = n4879 | n18555 ;
  assign n18557 = ( n15573 & n18555 ) | ( n15573 & n18556 ) | ( n18555 & n18556 ) ;
  assign n18558 = x20 & ~n18557 ;
  assign n18559 = ( ~x20 & n18551 ) | ( ~x20 & n18557 ) | ( n18551 & n18557 ) ;
  assign n18560 = ( ~n18552 & n18558 ) | ( ~n18552 & n18559 ) | ( n18558 & n18559 ) ;
  assign n18561 = n4637 & ~n14723 ;
  assign n18562 = x23 & n18561 ;
  assign n18563 = n4584 & n14520 ;
  assign n18564 = n4649 | n18563 ;
  assign n18565 = ( n14942 & n18563 ) | ( n14942 & n18564 ) | ( n18563 & n18564 ) ;
  assign n18566 = n4591 | n18565 ;
  assign n18567 = ( ~n14953 & n18565 ) | ( ~n14953 & n18566 ) | ( n18565 & n18566 ) ;
  assign n18568 = x23 & ~n18567 ;
  assign n18569 = ( ~x23 & n18561 ) | ( ~x23 & n18567 ) | ( n18561 & n18567 ) ;
  assign n18570 = ( ~n18562 & n18568 ) | ( ~n18562 & n18569 ) | ( n18568 & n18569 ) ;
  assign n18571 = n4215 & n14352 ;
  assign n18572 = n4200 & n13992 ;
  assign n18573 = n2083 & n13996 ;
  assign n18574 = n18572 | n18573 ;
  assign n18575 = n18571 | n18574 ;
  assign n18576 = x26 & n18575 ;
  assign n18577 = n4203 & n14363 ;
  assign n18578 = ( ~x26 & n18575 ) | ( ~x26 & n18577 ) | ( n18575 & n18577 ) ;
  assign n18579 = x26 & ~n18577 ;
  assign n18580 = ( ~n18576 & n18578 ) | ( ~n18576 & n18579 ) | ( n18578 & n18579 ) ;
  assign n18581 = n3501 & ~n14000 ;
  assign n18582 = x29 & n18581 ;
  assign n18583 = n3536 & ~n14007 ;
  assign n18584 = n4039 | n18583 ;
  assign n18585 = ( n13998 & n18583 ) | ( n13998 & n18584 ) | ( n18583 & n18584 ) ;
  assign n18586 = n3541 | n18585 ;
  assign n18587 = ( n14115 & n18585 ) | ( n14115 & n18586 ) | ( n18585 & n18586 ) ;
  assign n18588 = x29 & ~n18587 ;
  assign n18589 = ( ~x29 & n18581 ) | ( ~x29 & n18587 ) | ( n18581 & n18587 ) ;
  assign n18590 = ( ~n18582 & n18588 ) | ( ~n18582 & n18589 ) | ( n18588 & n18589 ) ;
  assign n18591 = n3273 & ~n14014 ;
  assign n18592 = n3270 | n18591 ;
  assign n18593 = ( n14002 & n18591 ) | ( n14002 & n18592 ) | ( n18591 & n18592 ) ;
  assign n18594 = n390 | n18593 ;
  assign n18595 = ( n14072 & n18593 ) | ( n14072 & n18594 ) | ( n18593 & n18594 ) ;
  assign n18596 = n3274 & ~n14004 ;
  assign n18597 = n18595 | n18596 ;
  assign n18598 = n150 | n616 ;
  assign n18599 = n331 | n18598 ;
  assign n18600 = n550 | n704 ;
  assign n18601 = n131 | n413 ;
  assign n18602 = n18600 | n18601 ;
  assign n18603 = n18599 | n18602 ;
  assign n18604 = n1196 | n18603 ;
  assign n18605 = n3807 | n18604 ;
  assign n18606 = n1640 | n14882 ;
  assign n18607 = n18605 | n18606 ;
  assign n18608 = n13613 | n18607 ;
  assign n18609 = n262 | n1100 ;
  assign n18610 = n696 | n18609 ;
  assign n18611 = n4113 | n18610 ;
  assign n18612 = n16102 | n16688 ;
  assign n18613 = n18611 | n18612 ;
  assign n18614 = n5026 & ~n18613 ;
  assign n18615 = ~n6100 & n18614 ;
  assign n18616 = ~n18608 & n18615 ;
  assign n18617 = ( n18501 & n18597 ) | ( n18501 & ~n18616 ) | ( n18597 & ~n18616 ) ;
  assign n18618 = ( n18501 & ~n18597 ) | ( n18501 & n18616 ) | ( ~n18597 & n18616 ) ;
  assign n18619 = ( ~n18501 & n18617 ) | ( ~n18501 & n18618 ) | ( n18617 & n18618 ) ;
  assign n18620 = ( n18506 & ~n18590 ) | ( n18506 & n18619 ) | ( ~n18590 & n18619 ) ;
  assign n18621 = ( n18506 & n18590 ) | ( n18506 & ~n18619 ) | ( n18590 & ~n18619 ) ;
  assign n18622 = ( ~n18506 & n18620 ) | ( ~n18506 & n18621 ) | ( n18620 & n18621 ) ;
  assign n18623 = ( n18510 & ~n18580 ) | ( n18510 & n18622 ) | ( ~n18580 & n18622 ) ;
  assign n18624 = ( n18510 & n18580 ) | ( n18510 & ~n18622 ) | ( n18580 & ~n18622 ) ;
  assign n18625 = ( ~n18510 & n18623 ) | ( ~n18510 & n18624 ) | ( n18623 & n18624 ) ;
  assign n18626 = ( n18512 & n18570 ) | ( n18512 & ~n18625 ) | ( n18570 & ~n18625 ) ;
  assign n18627 = ( n18512 & ~n18570 ) | ( n18512 & n18625 ) | ( ~n18570 & n18625 ) ;
  assign n18628 = ( ~n18512 & n18626 ) | ( ~n18512 & n18627 ) | ( n18626 & n18627 ) ;
  assign n18629 = ( n18515 & n18560 ) | ( n18515 & ~n18628 ) | ( n18560 & ~n18628 ) ;
  assign n18630 = ( n18515 & ~n18560 ) | ( n18515 & n18628 ) | ( ~n18560 & n18628 ) ;
  assign n18631 = ( ~n18515 & n18629 ) | ( ~n18515 & n18630 ) | ( n18629 & n18630 ) ;
  assign n18632 = ( n18518 & ~n18550 ) | ( n18518 & n18631 ) | ( ~n18550 & n18631 ) ;
  assign n18633 = ( n18518 & n18550 ) | ( n18518 & ~n18631 ) | ( n18550 & ~n18631 ) ;
  assign n18634 = ( ~n18518 & n18632 ) | ( ~n18518 & n18633 ) | ( n18632 & n18633 ) ;
  assign n18635 = n6332 & ~n16531 ;
  assign n18636 = x14 & n18635 ;
  assign n18637 = n5909 & ~n16338 ;
  assign n18638 = n5914 | n18637 ;
  assign n18639 = ( n16724 & n18637 ) | ( n16724 & n18638 ) | ( n18637 & n18638 ) ;
  assign n18640 = n5915 | n18639 ;
  assign n18641 = ( n16735 & n18639 ) | ( n16735 & n18640 ) | ( n18639 & n18640 ) ;
  assign n18642 = x14 & ~n18641 ;
  assign n18643 = ( ~x14 & n18635 ) | ( ~x14 & n18641 ) | ( n18635 & n18641 ) ;
  assign n18644 = ( ~n18636 & n18642 ) | ( ~n18636 & n18643 ) | ( n18642 & n18643 ) ;
  assign n18645 = ( n18522 & n18634 ) | ( n18522 & ~n18644 ) | ( n18634 & ~n18644 ) ;
  assign n18646 = ( n18522 & ~n18634 ) | ( n18522 & n18644 ) | ( ~n18634 & n18644 ) ;
  assign n18647 = ( ~n18522 & n18645 ) | ( ~n18522 & n18646 ) | ( n18645 & n18646 ) ;
  assign n18648 = ( n18524 & ~n18540 ) | ( n18524 & n18647 ) | ( ~n18540 & n18647 ) ;
  assign n18649 = ( n18524 & n18540 ) | ( n18524 & ~n18647 ) | ( n18540 & ~n18647 ) ;
  assign n18650 = ( ~n18524 & n18648 ) | ( ~n18524 & n18649 ) | ( n18648 & n18649 ) ;
  assign n18651 = n7346 & ~n17976 ;
  assign n18652 = x8 & n18651 ;
  assign n18653 = n7341 & ~n17635 ;
  assign n18654 = n7345 | n18653 ;
  assign n18655 = ( ~n17963 & n18653 ) | ( ~n17963 & n18654 ) | ( n18653 & n18654 ) ;
  assign n18656 = n7644 & n17742 ;
  assign n18657 = n18655 | n18656 ;
  assign n18658 = x8 & ~n18657 ;
  assign n18659 = ( ~x8 & n18651 ) | ( ~x8 & n18657 ) | ( n18651 & n18657 ) ;
  assign n18660 = ( ~n18652 & n18658 ) | ( ~n18652 & n18659 ) | ( n18658 & n18659 ) ;
  assign n18661 = ( n18527 & ~n18650 ) | ( n18527 & n18660 ) | ( ~n18650 & n18660 ) ;
  assign n18662 = ( n18527 & n18650 ) | ( n18527 & ~n18660 ) | ( n18650 & ~n18660 ) ;
  assign n18663 = ( ~n18527 & n18661 ) | ( ~n18527 & n18662 ) | ( n18661 & n18662 ) ;
  assign n18664 = n18362 | n18370 ;
  assign n18665 = n2083 & ~n10235 ;
  assign n18666 = x26 & n18665 ;
  assign n18667 = n4215 & ~n13473 ;
  assign n18668 = n4200 & ~n13280 ;
  assign n18669 = n18667 | n18668 ;
  assign n18670 = n4203 | n18669 ;
  assign n18671 = ( ~n13480 & n18669 ) | ( ~n13480 & n18670 ) | ( n18669 & n18670 ) ;
  assign n18672 = x26 & ~n18671 ;
  assign n18673 = ( ~x26 & n18665 ) | ( ~x26 & n18671 ) | ( n18665 & n18671 ) ;
  assign n18674 = ( ~n18666 & n18672 ) | ( ~n18666 & n18673 ) | ( n18672 & n18673 ) ;
  assign n18675 = n3501 & ~n10237 ;
  assign n18676 = x29 & n18675 ;
  assign n18677 = n3536 & ~n10332 ;
  assign n18678 = n4039 | n18677 ;
  assign n18679 = ( n10214 & n18677 ) | ( n10214 & n18678 ) | ( n18677 & n18678 ) ;
  assign n18680 = n3541 | n18679 ;
  assign n18681 = ( n12953 & n18679 ) | ( n12953 & n18680 ) | ( n18679 & n18680 ) ;
  assign n18682 = x29 & ~n18681 ;
  assign n18683 = ( ~x29 & n18675 ) | ( ~x29 & n18681 ) | ( n18675 & n18681 ) ;
  assign n18684 = ( ~n18676 & n18682 ) | ( ~n18676 & n18683 ) | ( n18682 & n18683 ) ;
  assign n18685 = n2178 | n2214 ;
  assign n18686 = n12837 | n18685 ;
  assign n18687 = n14872 | n18686 ;
  assign n18688 = n3182 | n3450 ;
  assign n18689 = n18687 | n18688 ;
  assign n18690 = n233 | n497 ;
  assign n18691 = n329 | n356 ;
  assign n18692 = n18690 | n18691 ;
  assign n18693 = n1862 | n18692 ;
  assign n18694 = n373 | n533 ;
  assign n18695 = n97 | n18694 ;
  assign n18696 = n18693 | n18695 ;
  assign n18697 = n208 | n270 ;
  assign n18698 = n206 | n18697 ;
  assign n18699 = n18696 | n18698 ;
  assign n18700 = n18689 | n18699 ;
  assign n18701 = n2100 | n18700 ;
  assign n18702 = n3341 | n18701 ;
  assign n18703 = n3273 & n10239 ;
  assign n18704 = n3270 | n18703 ;
  assign n18705 = ( n10329 & n18703 ) | ( n10329 & n18704 ) | ( n18703 & n18704 ) ;
  assign n18706 = n390 | n18705 ;
  assign n18707 = ( n10397 & n18705 ) | ( n10397 & n18706 ) | ( n18705 & n18706 ) ;
  assign n18708 = n3274 & n10326 ;
  assign n18709 = n18707 | n18708 ;
  assign n18710 = ( n18346 & n18702 ) | ( n18346 & n18709 ) | ( n18702 & n18709 ) ;
  assign n18711 = ( n18346 & ~n18702 ) | ( n18346 & n18709 ) | ( ~n18702 & n18709 ) ;
  assign n18712 = ( n18702 & ~n18710 ) | ( n18702 & n18711 ) | ( ~n18710 & n18711 ) ;
  assign n18713 = ( ~n18348 & n18684 ) | ( ~n18348 & n18712 ) | ( n18684 & n18712 ) ;
  assign n18714 = ( n18348 & n18684 ) | ( n18348 & n18712 ) | ( n18684 & n18712 ) ;
  assign n18715 = ( n18348 & n18713 ) | ( n18348 & ~n18714 ) | ( n18713 & ~n18714 ) ;
  assign n18716 = ( n18351 & n18674 ) | ( n18351 & n18715 ) | ( n18674 & n18715 ) ;
  assign n18717 = ( n18351 & ~n18674 ) | ( n18351 & n18715 ) | ( ~n18674 & n18715 ) ;
  assign n18718 = ( n18674 & ~n18716 ) | ( n18674 & n18717 ) | ( ~n18716 & n18717 ) ;
  assign n18719 = ( x20 & ~x21 ) | ( x20 & x22 ) | ( ~x21 & x22 ) ;
  assign n18720 = ( x21 & ~x23 ) | ( x21 & n18719 ) | ( ~x23 & n18719 ) ;
  assign n18721 = ~n4583 & n18720 ;
  assign n18722 = ( n13475 & n18720 ) | ( n13475 & n18721 ) | ( n18720 & n18721 ) ;
  assign n18723 = n4580 & ~n13475 ;
  assign n18724 = n18722 | n18723 ;
  assign n18725 = ( n18354 & ~n18718 ) | ( n18354 & n18724 ) | ( ~n18718 & n18724 ) ;
  assign n18726 = ( n18354 & n18718 ) | ( n18354 & n18724 ) | ( n18718 & n18724 ) ;
  assign n18727 = ( n18718 & n18725 ) | ( n18718 & ~n18726 ) | ( n18725 & ~n18726 ) ;
  assign n18728 = ( n18357 & ~n18360 ) | ( n18357 & n18727 ) | ( ~n18360 & n18727 ) ;
  assign n18729 = ( n18357 & n18360 ) | ( n18357 & n18727 ) | ( n18360 & n18727 ) ;
  assign n18730 = ( n18360 & n18728 ) | ( n18360 & ~n18729 ) | ( n18728 & ~n18729 ) ;
  assign n18731 = ~n18664 & n18730 ;
  assign n18732 = n18266 & n18362 ;
  assign n18733 = ( n18664 & n18730 ) | ( n18664 & ~n18732 ) | ( n18730 & ~n18732 ) ;
  assign n18734 = n18730 & ~n18732 ;
  assign n18735 = ( n18731 & n18733 ) | ( n18731 & ~n18734 ) | ( n18733 & ~n18734 ) ;
  assign n18736 = n40 & n18730 ;
  assign n18737 = n8341 | n18736 ;
  assign n18738 = ( n18735 & n18736 ) | ( n18735 & n18737 ) | ( n18736 & n18737 ) ;
  assign n18739 = n8340 & ~n18258 ;
  assign n18740 = ( ~x5 & n18738 ) | ( ~x5 & n18739 ) | ( n18738 & n18739 ) ;
  assign n18741 = n8721 & ~n18362 ;
  assign n18742 = x5 & ~n18739 ;
  assign n18743 = n18741 | n18742 ;
  assign n18744 = ( n18738 & n18741 ) | ( n18738 & n18742 ) | ( n18741 & n18742 ) ;
  assign n18745 = ( n18740 & n18743 ) | ( n18740 & ~n18744 ) | ( n18743 & ~n18744 ) ;
  assign n18746 = ( n18530 & ~n18663 ) | ( n18530 & n18745 ) | ( ~n18663 & n18745 ) ;
  assign n18747 = ( n18530 & n18663 ) | ( n18530 & ~n18745 ) | ( n18663 & ~n18745 ) ;
  assign n18748 = ( ~n18530 & n18746 ) | ( ~n18530 & n18747 ) | ( n18746 & n18747 ) ;
  assign n18749 = ( ~n9590 & n9591 ) | ( ~n9590 & n15195 ) | ( n9591 & n15195 ) ;
  assign n18750 = n9600 & ~n14723 ;
  assign n18751 = n9592 | n18750 ;
  assign n18752 = ~n18749 & n18751 ;
  assign n18753 = n9591 & ~n15195 ;
  assign n18754 = n9593 & ~n15184 ;
  assign n18755 = n41 & n14942 ;
  assign n18756 = n18754 | n18755 ;
  assign n18757 = ~x2 & n18756 ;
  assign n18758 = ( ~x2 & n18753 ) | ( ~x2 & n18757 ) | ( n18753 & n18757 ) ;
  assign n18759 = x2 | n18756 ;
  assign n18760 = ( n18752 & ~n18756 ) | ( n18752 & n18759 ) | ( ~n18756 & n18759 ) ;
  assign n18761 = ( ~n18752 & n18758 ) | ( ~n18752 & n18760 ) | ( n18758 & n18760 ) ;
  assign n18762 = ( ~n14368 & n14535 ) | ( ~n14368 & n14564 ) | ( n14535 & n14564 ) ;
  assign n18763 = ( n14368 & ~n14565 ) | ( n14368 & n18762 ) | ( ~n14565 & n18762 ) ;
  assign n18764 = n41 & ~n14723 ;
  assign n18765 = x2 & n18764 ;
  assign n18766 = n9600 & n14520 ;
  assign n18767 = n9593 | n18766 ;
  assign n18768 = ( n14942 & n18766 ) | ( n14942 & n18767 ) | ( n18766 & n18767 ) ;
  assign n18769 = n9592 | n18768 ;
  assign n18770 = ( ~n14953 & n18768 ) | ( ~n14953 & n18769 ) | ( n18768 & n18769 ) ;
  assign n18771 = x2 & ~n18770 ;
  assign n18772 = ( ~x2 & n18764 ) | ( ~x2 & n18770 ) | ( n18764 & n18770 ) ;
  assign n18773 = ( ~n18765 & n18771 ) | ( ~n18765 & n18772 ) | ( n18771 & n18772 ) ;
  assign n18774 = ( ~n14177 & n14203 ) | ( ~n14177 & n14367 ) | ( n14203 & n14367 ) ;
  assign n18775 = ( n14177 & ~n14368 ) | ( n14177 & n18774 ) | ( ~n14368 & n18774 ) ;
  assign n18776 = n41 & n14520 ;
  assign n18777 = x2 & n18776 ;
  assign n18778 = n9600 & n14352 ;
  assign n18779 = n9593 | n18778 ;
  assign n18780 = ( ~n14723 & n18778 ) | ( ~n14723 & n18779 ) | ( n18778 & n18779 ) ;
  assign n18781 = n9592 | n18780 ;
  assign n18782 = ( ~n14734 & n18780 ) | ( ~n14734 & n18781 ) | ( n18780 & n18781 ) ;
  assign n18783 = x2 & ~n18782 ;
  assign n18784 = ( ~x2 & n18776 ) | ( ~x2 & n18782 ) | ( n18776 & n18782 ) ;
  assign n18785 = ( ~n18777 & n18783 ) | ( ~n18777 & n18784 ) | ( n18783 & n18784 ) ;
  assign n18786 = ( ~n14032 & n14152 ) | ( ~n14032 & n14176 ) | ( n14152 & n14176 ) ;
  assign n18787 = ( n14032 & ~n14177 ) | ( n14032 & n18786 ) | ( ~n14177 & n18786 ) ;
  assign n18788 = n9592 & ~n14130 ;
  assign n18789 = x2 & n18788 ;
  assign n18790 = n9600 & ~n14000 ;
  assign n18791 = n9593 | n18790 ;
  assign n18792 = ( n13996 & n18790 ) | ( n13996 & n18791 ) | ( n18790 & n18791 ) ;
  assign n18793 = n41 & n13998 ;
  assign n18794 = n18792 | n18793 ;
  assign n18795 = x2 & ~n18794 ;
  assign n18796 = ( ~x2 & n18788 ) | ( ~x2 & n18794 ) | ( n18788 & n18794 ) ;
  assign n18797 = ( ~n18789 & n18795 ) | ( ~n18789 & n18796 ) | ( n18795 & n18796 ) ;
  assign n18798 = n41 & ~n14000 ;
  assign n18799 = n9592 | n18798 ;
  assign n18800 = ( n14115 & n18798 ) | ( n14115 & n18799 ) | ( n18798 & n18799 ) ;
  assign n18801 = n9593 & n13998 ;
  assign n18802 = ( x2 & ~n18800 ) | ( x2 & n18801 ) | ( ~n18800 & n18801 ) ;
  assign n18803 = ~x2 & n18800 ;
  assign n18804 = n9600 & ~n14007 ;
  assign n18805 = ( x2 & n18801 ) | ( x2 & n18804 ) | ( n18801 & n18804 ) ;
  assign n18806 = ( n18802 & n18803 ) | ( n18802 & ~n18805 ) | ( n18803 & ~n18805 ) ;
  assign n18807 = n9158 & ~n14042 ;
  assign n18808 = n9593 & ~n14000 ;
  assign n18809 = n41 & ~n14007 ;
  assign n18810 = n18808 | n18809 ;
  assign n18811 = x2 | n18810 ;
  assign n18812 = n18807 | n18811 ;
  assign n18813 = n9589 & ~n14042 ;
  assign n18814 = n9600 & n14002 ;
  assign n18815 = ( x2 & n18810 ) | ( x2 & n18814 ) | ( n18810 & n18814 ) ;
  assign n18816 = n18813 | n18815 ;
  assign n18817 = n18812 & ~n18816 ;
  assign n18818 = ~x0 & n14004 ;
  assign n18819 = ( ~n14002 & n14004 ) | ( ~n14002 & n18818 ) | ( n14004 & n18818 ) ;
  assign n18820 = n34 & ~n14014 ;
  assign n18821 = n9155 & n14014 ;
  assign n18822 = n18820 | n18821 ;
  assign n18823 = ( ~n18819 & n18820 ) | ( ~n18819 & n18822 ) | ( n18820 & n18822 ) ;
  assign n18824 = n9600 & ~n14004 ;
  assign n18825 = n9593 | n18824 ;
  assign n18826 = ( ~n14007 & n18824 ) | ( ~n14007 & n18825 ) | ( n18824 & n18825 ) ;
  assign n18827 = n9592 | n18826 ;
  assign n18828 = ( n14066 & n18826 ) | ( n14066 & n18827 ) | ( n18826 & n18827 ) ;
  assign n18829 = n41 & n14002 ;
  assign n18830 = n18828 | n18829 ;
  assign n18831 = x3 & ~n14014 ;
  assign n18832 = n18830 & n18831 ;
  assign n18833 = x2 & ~n18830 ;
  assign n18834 = ( ~n18823 & n18832 ) | ( ~n18823 & n18833 ) | ( n18832 & n18833 ) ;
  assign n18835 = ~n14084 & n14085 ;
  assign n18836 = n14084 & ~n14085 ;
  assign n18837 = n18835 | n18836 ;
  assign n18838 = ( n18817 & n18834 ) | ( n18817 & n18837 ) | ( n18834 & n18837 ) ;
  assign n18839 = n14079 & n14086 ;
  assign n18840 = n14087 & ~n18839 ;
  assign n18841 = ( n18806 & n18838 ) | ( n18806 & n18840 ) | ( n18838 & n18840 ) ;
  assign n18842 = ( n14092 & n18797 ) | ( n14092 & n18841 ) | ( n18797 & n18841 ) ;
  assign n18843 = n9593 & n13992 ;
  assign n18844 = x2 & n18843 ;
  assign n18845 = n41 & n13996 ;
  assign n18846 = n9600 & n13998 ;
  assign n18847 = n18845 | n18846 ;
  assign n18848 = n9592 | n18847 ;
  assign n18849 = ( n14024 & n18847 ) | ( n14024 & n18848 ) | ( n18847 & n18848 ) ;
  assign n18850 = x2 & ~n18849 ;
  assign n18851 = ( ~x2 & n18843 ) | ( ~x2 & n18849 ) | ( n18843 & n18849 ) ;
  assign n18852 = ( ~n18844 & n18850 ) | ( ~n18844 & n18851 ) | ( n18850 & n18851 ) ;
  assign n18853 = ( ~n14046 & n14057 ) | ( ~n14046 & n14093 ) | ( n14057 & n14093 ) ;
  assign n18854 = ( n14046 & ~n14094 ) | ( n14046 & n18853 ) | ( ~n14094 & n18853 ) ;
  assign n18855 = ( n18842 & n18852 ) | ( n18842 & n18854 ) | ( n18852 & n18854 ) ;
  assign n18856 = ( ~n14094 & n14106 ) | ( ~n14094 & n14119 ) | ( n14106 & n14119 ) ;
  assign n18857 = ( n14094 & ~n14120 ) | ( n14094 & n18856 ) | ( ~n14120 & n18856 ) ;
  assign n18858 = n9592 & n14363 ;
  assign n18859 = n9593 & n14352 ;
  assign n18860 = n41 & n13992 ;
  assign n18861 = n18859 | n18860 ;
  assign n18862 = x2 | n18861 ;
  assign n18863 = ( ~n18858 & n18861 ) | ( ~n18858 & n18862 ) | ( n18861 & n18862 ) ;
  assign n18864 = n9591 & n14363 ;
  assign n18865 = n18863 | n18864 ;
  assign n18866 = n9600 & n13996 ;
  assign n18867 = ( x2 & n18861 ) | ( x2 & n18866 ) | ( n18861 & n18866 ) ;
  assign n18868 = n18865 & ~n18867 ;
  assign n18869 = ( n18855 & n18857 ) | ( n18855 & n18868 ) | ( n18857 & n18868 ) ;
  assign n18870 = n9592 & n14531 ;
  assign n18871 = n9593 & n14520 ;
  assign n18872 = n41 & n14352 ;
  assign n18873 = n18871 | n18872 ;
  assign n18874 = x2 | n18873 ;
  assign n18875 = ( ~n18870 & n18873 ) | ( ~n18870 & n18874 ) | ( n18873 & n18874 ) ;
  assign n18876 = n9591 & n14531 ;
  assign n18877 = n18875 | n18876 ;
  assign n18878 = n9600 & n13992 ;
  assign n18879 = ( x2 & n18873 ) | ( x2 & n18878 ) | ( n18873 & n18878 ) ;
  assign n18880 = n18877 & ~n18879 ;
  assign n18881 = ( ~n14120 & n14134 ) | ( ~n14120 & n14151 ) | ( n14134 & n14151 ) ;
  assign n18882 = ( n14120 & ~n14152 ) | ( n14120 & n18881 ) | ( ~n14152 & n18881 ) ;
  assign n18883 = ( n18869 & n18880 ) | ( n18869 & n18882 ) | ( n18880 & n18882 ) ;
  assign n18884 = ( n18785 & n18787 ) | ( n18785 & n18883 ) | ( n18787 & n18883 ) ;
  assign n18885 = ( n18773 & n18775 ) | ( n18773 & n18884 ) | ( n18775 & n18884 ) ;
  assign n18886 = ( n18761 & n18763 ) | ( n18761 & n18885 ) | ( n18763 & n18885 ) ;
  assign n18887 = n41 & ~n15184 ;
  assign n18888 = x2 & n18887 ;
  assign n18889 = n9600 & n14942 ;
  assign n18890 = n9593 | n18889 ;
  assign n18891 = ( ~n15394 & n18889 ) | ( ~n15394 & n18890 ) | ( n18889 & n18890 ) ;
  assign n18892 = n9592 | n18891 ;
  assign n18893 = ( n15405 & n18891 ) | ( n15405 & n18892 ) | ( n18891 & n18892 ) ;
  assign n18894 = x2 & ~n18893 ;
  assign n18895 = ( ~x2 & n18887 ) | ( ~x2 & n18893 ) | ( n18887 & n18893 ) ;
  assign n18896 = ( ~n18888 & n18894 ) | ( ~n18888 & n18895 ) | ( n18894 & n18895 ) ;
  assign n18897 = ( ~n14565 & n14738 ) | ( ~n14565 & n14774 ) | ( n14738 & n14774 ) ;
  assign n18898 = ( n14565 & ~n14775 ) | ( n14565 & n18897 ) | ( ~n14775 & n18897 ) ;
  assign n18899 = ( n18886 & n18896 ) | ( n18886 & n18898 ) | ( n18896 & n18898 ) ;
  assign n18900 = n9593 & n15561 ;
  assign n18901 = n41 & ~n15394 ;
  assign n18902 = n18900 | n18901 ;
  assign n18903 = x2 & n18902 ;
  assign n18904 = ~x2 & n18902 ;
  assign n18905 = n9600 & ~n15184 ;
  assign n18906 = ( x2 & n9590 ) | ( x2 & ~n15573 ) | ( n9590 & ~n15573 ) ;
  assign n18907 = n9591 & n15573 ;
  assign n18908 = ( ~n18905 & n18906 ) | ( ~n18905 & n18907 ) | ( n18906 & n18907 ) ;
  assign n18909 = ( ~n18903 & n18904 ) | ( ~n18903 & n18908 ) | ( n18904 & n18908 ) ;
  assign n18910 = ( ~n14775 & n14957 ) | ( ~n14775 & n14996 ) | ( n14957 & n14996 ) ;
  assign n18911 = ( n14775 & ~n14997 ) | ( n14775 & n18910 ) | ( ~n14997 & n18910 ) ;
  assign n18912 = ( n18899 & n18909 ) | ( n18899 & n18911 ) | ( n18909 & n18911 ) ;
  assign n18913 = n9593 & ~n15806 ;
  assign n18914 = n41 & n15561 ;
  assign n18915 = n18913 | n18914 ;
  assign n18916 = n9639 | n18915 ;
  assign n18917 = x2 | n15817 ;
  assign n18918 = ~n9158 & n15817 ;
  assign n18919 = ( n18916 & n18917 ) | ( n18916 & ~n18918 ) | ( n18917 & ~n18918 ) ;
  assign n18920 = n9600 & ~n15394 ;
  assign n18921 = ( x2 & n18915 ) | ( x2 & n18920 ) | ( n18915 & n18920 ) ;
  assign n18922 = n18919 & ~n18921 ;
  assign n18923 = ( ~n14997 & n15039 ) | ( ~n14997 & n15199 ) | ( n15039 & n15199 ) ;
  assign n18924 = ( n14997 & ~n15200 ) | ( n14997 & n18923 ) | ( ~n15200 & n18923 ) ;
  assign n18925 = ( n18912 & n18922 ) | ( n18912 & n18924 ) | ( n18922 & n18924 ) ;
  assign n18926 = n41 & ~n15806 ;
  assign n18927 = x2 & n18926 ;
  assign n18928 = n9600 & n15561 ;
  assign n18929 = n9593 | n18928 ;
  assign n18930 = ( ~n15954 & n18928 ) | ( ~n15954 & n18929 ) | ( n18928 & n18929 ) ;
  assign n18931 = n9592 | n18930 ;
  assign n18932 = ( ~n15965 & n18930 ) | ( ~n15965 & n18931 ) | ( n18930 & n18931 ) ;
  assign n18933 = x2 & ~n18932 ;
  assign n18934 = ( ~x2 & n18926 ) | ( ~x2 & n18932 ) | ( n18926 & n18932 ) ;
  assign n18935 = ( ~n18927 & n18933 ) | ( ~n18927 & n18934 ) | ( n18933 & n18934 ) ;
  assign n18936 = ( ~n15200 & n15249 ) | ( ~n15200 & n15409 ) | ( n15249 & n15409 ) ;
  assign n18937 = ( n15200 & ~n15410 ) | ( n15200 & n18936 ) | ( ~n15410 & n18936 ) ;
  assign n18938 = ( n18925 & n18935 ) | ( n18925 & n18937 ) | ( n18935 & n18937 ) ;
  assign n18939 = n9592 & ~n16161 ;
  assign n18940 = n9593 & ~n16150 ;
  assign n18941 = n41 & ~n15954 ;
  assign n18942 = n18940 | n18941 ;
  assign n18943 = x2 | n18942 ;
  assign n18944 = ( ~n18939 & n18942 ) | ( ~n18939 & n18943 ) | ( n18942 & n18943 ) ;
  assign n18945 = n9591 & ~n16161 ;
  assign n18946 = n18944 | n18945 ;
  assign n18947 = n9600 & ~n15806 ;
  assign n18948 = ( x2 & n18942 ) | ( x2 & n18947 ) | ( n18942 & n18947 ) ;
  assign n18949 = n18946 & ~n18948 ;
  assign n18950 = ( ~n15410 & n15577 ) | ( ~n15410 & n15629 ) | ( n15577 & n15629 ) ;
  assign n18951 = ( n15410 & ~n15630 ) | ( n15410 & n18950 ) | ( ~n15630 & n18950 ) ;
  assign n18952 = ( n18938 & n18949 ) | ( n18938 & n18951 ) | ( n18949 & n18951 ) ;
  assign n18953 = n9593 & ~n16338 ;
  assign n18954 = n41 & ~n16150 ;
  assign n18955 = n18953 | n18954 ;
  assign n18956 = ~x2 & n18955 ;
  assign n18957 = n9591 & ~n16349 ;
  assign n18958 = ( x2 & ~n18955 ) | ( x2 & n18957 ) | ( ~n18955 & n18957 ) ;
  assign n18959 = ( ~n9590 & n9591 ) | ( ~n9590 & n16349 ) | ( n9591 & n16349 ) ;
  assign n18960 = n9600 & ~n15954 ;
  assign n18961 = n9592 | n18960 ;
  assign n18962 = ~n18959 & n18961 ;
  assign n18963 = n18958 & ~n18962 ;
  assign n18964 = n18956 | n18963 ;
  assign n18965 = ( ~n15630 & n15685 ) | ( ~n15630 & n15821 ) | ( n15685 & n15821 ) ;
  assign n18966 = ( n15630 & ~n15822 ) | ( n15630 & n18965 ) | ( ~n15822 & n18965 ) ;
  assign n18967 = ( n18952 & n18964 ) | ( n18952 & n18966 ) | ( n18964 & n18966 ) ;
  assign n18968 = n41 & ~n16338 ;
  assign n18969 = x2 & n18968 ;
  assign n18970 = n9600 & ~n16150 ;
  assign n18971 = n9593 | n18970 ;
  assign n18972 = ( ~n16531 & n18970 ) | ( ~n16531 & n18971 ) | ( n18970 & n18971 ) ;
  assign n18973 = n9592 | n18972 ;
  assign n18974 = ( ~n16542 & n18972 ) | ( ~n16542 & n18973 ) | ( n18972 & n18973 ) ;
  assign n18975 = x2 & ~n18974 ;
  assign n18976 = ( ~x2 & n18968 ) | ( ~x2 & n18974 ) | ( n18968 & n18974 ) ;
  assign n18977 = ( ~n18969 & n18975 ) | ( ~n18969 & n18976 ) | ( n18975 & n18976 ) ;
  assign n18978 = ( ~n15822 & n15969 ) | ( ~n15822 & n16031 ) | ( n15969 & n16031 ) ;
  assign n18979 = ( n15822 & ~n16032 ) | ( n15822 & n18978 ) | ( ~n16032 & n18978 ) ;
  assign n18980 = ( n18967 & n18977 ) | ( n18967 & n18979 ) | ( n18977 & n18979 ) ;
  assign n18981 = n41 & ~n16531 ;
  assign n18982 = x2 & n18981 ;
  assign n18983 = n9600 & ~n16338 ;
  assign n18984 = n9593 | n18983 ;
  assign n18985 = ( n16724 & n18983 ) | ( n16724 & n18984 ) | ( n18983 & n18984 ) ;
  assign n18986 = n9592 | n18985 ;
  assign n18987 = ( n16735 & n18985 ) | ( n16735 & n18986 ) | ( n18985 & n18986 ) ;
  assign n18988 = x2 & ~n18987 ;
  assign n18989 = ( ~x2 & n18981 ) | ( ~x2 & n18987 ) | ( n18981 & n18987 ) ;
  assign n18990 = ( ~n18982 & n18988 ) | ( ~n18982 & n18989 ) | ( n18988 & n18989 ) ;
  assign n18991 = ( ~n16032 & n16165 ) | ( ~n16032 & n16230 ) | ( n16165 & n16230 ) ;
  assign n18992 = ( n16032 & ~n16231 ) | ( n16032 & n18991 ) | ( ~n16231 & n18991 ) ;
  assign n18993 = ( n18980 & n18990 ) | ( n18980 & n18992 ) | ( n18990 & n18992 ) ;
  assign n18994 = n41 & n16724 ;
  assign n18995 = x2 & n18994 ;
  assign n18996 = n9600 & ~n16531 ;
  assign n18997 = n9593 | n18996 ;
  assign n18998 = ( n16925 & n18996 ) | ( n16925 & n18997 ) | ( n18996 & n18997 ) ;
  assign n18999 = n9592 | n18998 ;
  assign n19000 = ( ~n16936 & n18998 ) | ( ~n16936 & n18999 ) | ( n18998 & n18999 ) ;
  assign n19001 = x2 & ~n19000 ;
  assign n19002 = ( ~x2 & n18994 ) | ( ~x2 & n19000 ) | ( n18994 & n19000 ) ;
  assign n19003 = ( ~n18995 & n19001 ) | ( ~n18995 & n19002 ) | ( n19001 & n19002 ) ;
  assign n19004 = ( ~n16231 & n16353 ) | ( ~n16231 & n16421 ) | ( n16353 & n16421 ) ;
  assign n19005 = ( n16231 & ~n16422 ) | ( n16231 & n19004 ) | ( ~n16422 & n19004 ) ;
  assign n19006 = ( n18993 & n19003 ) | ( n18993 & n19005 ) | ( n19003 & n19005 ) ;
  assign n19007 = n41 & n16925 ;
  assign n19008 = x2 & n19007 ;
  assign n19009 = n9600 & n16724 ;
  assign n19010 = n9593 | n19009 ;
  assign n19011 = ( ~n17126 & n19009 ) | ( ~n17126 & n19010 ) | ( n19009 & n19010 ) ;
  assign n19012 = n9592 | n19011 ;
  assign n19013 = ( ~n17139 & n19011 ) | ( ~n17139 & n19012 ) | ( n19011 & n19012 ) ;
  assign n19014 = x2 & ~n19013 ;
  assign n19015 = ( ~x2 & n19007 ) | ( ~x2 & n19013 ) | ( n19007 & n19013 ) ;
  assign n19016 = ( ~n19008 & n19014 ) | ( ~n19008 & n19015 ) | ( n19014 & n19015 ) ;
  assign n19017 = ( ~n16422 & n16546 ) | ( ~n16422 & n16621 ) | ( n16546 & n16621 ) ;
  assign n19018 = ( n16422 & ~n16622 ) | ( n16422 & n19017 ) | ( ~n16622 & n19017 ) ;
  assign n19019 = ( n19006 & n19016 ) | ( n19006 & n19018 ) | ( n19016 & n19018 ) ;
  assign n19020 = ( ~n16622 & n16739 ) | ( ~n16622 & n16815 ) | ( n16739 & n16815 ) ;
  assign n19021 = ( n16622 & ~n16816 ) | ( n16622 & n19020 ) | ( ~n16816 & n19020 ) ;
  assign n19022 = n41 & ~n17126 ;
  assign n19023 = x2 & n19022 ;
  assign n19024 = n9600 & n16925 ;
  assign n19025 = n9593 | n19024 ;
  assign n19026 = ( n17346 & n19024 ) | ( n17346 & n19025 ) | ( n19024 & n19025 ) ;
  assign n19027 = n9592 | n19026 ;
  assign n19028 = ( ~n17356 & n19026 ) | ( ~n17356 & n19027 ) | ( n19026 & n19027 ) ;
  assign n19029 = x2 & ~n19028 ;
  assign n19030 = ( ~x2 & n19022 ) | ( ~x2 & n19028 ) | ( n19022 & n19028 ) ;
  assign n19031 = ( ~n19023 & n19029 ) | ( ~n19023 & n19030 ) | ( n19029 & n19030 ) ;
  assign n19032 = ( n19019 & n19021 ) | ( n19019 & n19031 ) | ( n19021 & n19031 ) ;
  assign n19033 = ( ~n16816 & n16940 ) | ( ~n16816 & n17020 ) | ( n16940 & n17020 ) ;
  assign n19034 = ( n16816 & ~n17021 ) | ( n16816 & n19033 ) | ( ~n17021 & n19033 ) ;
  assign n19035 = n41 & n17346 ;
  assign n19036 = n9592 | n19035 ;
  assign n19037 = ( ~n17646 & n19035 ) | ( ~n17646 & n19036 ) | ( n19035 & n19036 ) ;
  assign n19038 = n9593 & ~n17635 ;
  assign n19039 = ( x2 & ~n19037 ) | ( x2 & n19038 ) | ( ~n19037 & n19038 ) ;
  assign n19040 = ~x2 & n19037 ;
  assign n19041 = n9600 & ~n17126 ;
  assign n19042 = ( x2 & n19038 ) | ( x2 & n19041 ) | ( n19038 & n19041 ) ;
  assign n19043 = ( n19039 & n19040 ) | ( n19039 & ~n19042 ) | ( n19040 & ~n19042 ) ;
  assign n19044 = ( n19032 & n19034 ) | ( n19032 & n19043 ) | ( n19034 & n19043 ) ;
  assign n19045 = n9592 & ~n17749 ;
  assign n19046 = n9593 & n17742 ;
  assign n19047 = n41 & ~n17635 ;
  assign n19048 = n19046 | n19047 ;
  assign n19049 = x2 | n19048 ;
  assign n19050 = ( ~n19045 & n19048 ) | ( ~n19045 & n19049 ) | ( n19048 & n19049 ) ;
  assign n19051 = n9591 & ~n17749 ;
  assign n19052 = n19050 | n19051 ;
  assign n19053 = n9600 & n17346 ;
  assign n19054 = ( x2 & n19048 ) | ( x2 & n19053 ) | ( n19048 & n19053 ) ;
  assign n19055 = n19052 & ~n19054 ;
  assign n19056 = ( ~n17021 & n17143 ) | ( ~n17021 & n17233 ) | ( n17143 & n17233 ) ;
  assign n19057 = ( n17021 & ~n17234 ) | ( n17021 & n19056 ) | ( ~n17234 & n19056 ) ;
  assign n19058 = ( n19044 & n19055 ) | ( n19044 & n19057 ) | ( n19055 & n19057 ) ;
  assign n19059 = n41 & n17742 ;
  assign n19060 = x2 & n19059 ;
  assign n19061 = n9600 & ~n17635 ;
  assign n19062 = n9593 | n19061 ;
  assign n19063 = ( ~n17963 & n19061 ) | ( ~n17963 & n19062 ) | ( n19061 & n19062 ) ;
  assign n19064 = n9592 | n19063 ;
  assign n19065 = ( ~n17976 & n19063 ) | ( ~n17976 & n19064 ) | ( n19063 & n19064 ) ;
  assign n19066 = x2 & ~n19065 ;
  assign n19067 = ( ~x2 & n19059 ) | ( ~x2 & n19065 ) | ( n19059 & n19065 ) ;
  assign n19068 = ( ~n19060 & n19066 ) | ( ~n19060 & n19067 ) | ( n19066 & n19067 ) ;
  assign n19069 = ( ~n17234 & n17360 ) | ( ~n17234 & n17449 ) | ( n17360 & n17449 ) ;
  assign n19070 = ( n17234 & ~n17450 ) | ( n17234 & n19069 ) | ( ~n17450 & n19069 ) ;
  assign n19071 = ( n19058 & n19068 ) | ( n19058 & n19070 ) | ( n19068 & n19070 ) ;
  assign n19072 = n9593 & ~n18258 ;
  assign n19073 = n41 & ~n17963 ;
  assign n19074 = n19072 | n19073 ;
  assign n19075 = ~x2 & n19074 ;
  assign n19076 = x2 & n19074 ;
  assign n19077 = x2 & ~n18268 ;
  assign n19078 = n9591 & n18268 ;
  assign n19079 = ( ~n9590 & n19077 ) | ( ~n9590 & n19078 ) | ( n19077 & n19078 ) ;
  assign n19080 = ( n9159 & n9590 ) | ( n9159 & ~n17742 ) | ( n9590 & ~n17742 ) ;
  assign n19081 = n19079 | n19080 ;
  assign n19082 = ( n19075 & ~n19076 ) | ( n19075 & n19081 ) | ( ~n19076 & n19081 ) ;
  assign n19083 = ( ~n17450 & n17544 ) | ( ~n17450 & n17650 ) | ( n17544 & n17650 ) ;
  assign n19084 = ( n17450 & ~n17651 ) | ( n17450 & n19083 ) | ( ~n17651 & n19083 ) ;
  assign n19085 = ( n19071 & n19082 ) | ( n19071 & n19084 ) | ( n19082 & n19084 ) ;
  assign n19086 = ( ~n9590 & n9591 ) | ( ~n9590 & n18373 ) | ( n9591 & n18373 ) ;
  assign n19087 = n9600 & ~n17963 ;
  assign n19088 = n9592 | n19087 ;
  assign n19089 = ~n19086 & n19088 ;
  assign n19090 = n9591 & ~n18373 ;
  assign n19091 = n9593 & ~n18362 ;
  assign n19092 = n41 & ~n18258 ;
  assign n19093 = n19091 | n19092 ;
  assign n19094 = ~x2 & n19093 ;
  assign n19095 = ( ~x2 & n19090 ) | ( ~x2 & n19094 ) | ( n19090 & n19094 ) ;
  assign n19096 = x2 | n19093 ;
  assign n19097 = ( n19089 & ~n19093 ) | ( n19089 & n19096 ) | ( ~n19093 & n19096 ) ;
  assign n19098 = ( ~n19089 & n19095 ) | ( ~n19089 & n19097 ) | ( n19095 & n19097 ) ;
  assign n19099 = ( ~n17651 & n17757 ) | ( ~n17651 & n17859 ) | ( n17757 & n17859 ) ;
  assign n19100 = ( n17651 & ~n17860 ) | ( n17651 & n19099 ) | ( ~n17860 & n19099 ) ;
  assign n19101 = ( n19085 & n19098 ) | ( n19085 & n19100 ) | ( n19098 & n19100 ) ;
  assign n19102 = ( ~n17860 & n17980 ) | ( ~n17860 & n18082 ) | ( n17980 & n18082 ) ;
  assign n19103 = ( n17860 & ~n18083 ) | ( n17860 & n19102 ) | ( ~n18083 & n19102 ) ;
  assign n19104 = n41 & ~n18362 ;
  assign n19105 = n9592 | n19104 ;
  assign n19106 = ( n18735 & n19104 ) | ( n18735 & n19105 ) | ( n19104 & n19105 ) ;
  assign n19107 = n9593 & n18730 ;
  assign n19108 = ( x2 & ~n19106 ) | ( x2 & n19107 ) | ( ~n19106 & n19107 ) ;
  assign n19109 = ~x2 & n19106 ;
  assign n19110 = n9600 & ~n18258 ;
  assign n19111 = ( x2 & n19107 ) | ( x2 & n19110 ) | ( n19107 & n19110 ) ;
  assign n19112 = ( n19108 & n19109 ) | ( n19108 & ~n19111 ) | ( n19109 & ~n19111 ) ;
  assign n19113 = ( n19101 & n19103 ) | ( n19101 & n19112 ) | ( n19103 & n19112 ) ;
  assign n19114 = ( ~n18083 & n18187 ) | ( ~n18083 & n18272 ) | ( n18187 & n18272 ) ;
  assign n19115 = ( n18083 & ~n18273 ) | ( n18083 & n19114 ) | ( ~n18273 & n19114 ) ;
  assign n19116 = n3501 & n10214 ;
  assign n19117 = x29 & n19116 ;
  assign n19118 = n3536 & ~n10237 ;
  assign n19119 = n4039 | n19118 ;
  assign n19120 = ( ~n10235 & n19118 ) | ( ~n10235 & n19119 ) | ( n19118 & n19119 ) ;
  assign n19121 = n3541 | n19120 ;
  assign n19122 = ( n10371 & n19120 ) | ( n10371 & n19121 ) | ( n19120 & n19121 ) ;
  assign n19123 = x29 & ~n19122 ;
  assign n19124 = ( ~x29 & n19116 ) | ( ~x29 & n19122 ) | ( n19116 & n19122 ) ;
  assign n19125 = ( ~n19117 & n19123 ) | ( ~n19117 & n19124 ) | ( n19123 & n19124 ) ;
  assign n19126 = n1672 | n3080 ;
  assign n19127 = n1984 | n19126 ;
  assign n19128 = n3383 | n19127 ;
  assign n19129 = n3282 | n19128 ;
  assign n19130 = n532 | n1378 ;
  assign n19131 = n3293 | n19130 ;
  assign n19132 = n19129 | n19131 ;
  assign n19133 = n63 | n3448 ;
  assign n19134 = n1533 | n19133 ;
  assign n19135 = n650 | n19134 ;
  assign n19136 = n3804 | n5477 ;
  assign n19137 = n19135 | n19136 ;
  assign n19138 = n750 | n922 ;
  assign n19139 = n270 | n19138 ;
  assign n19140 = n3946 | n13047 ;
  assign n19141 = n19139 | n19140 ;
  assign n19142 = n19137 | n19141 ;
  assign n19143 = n19132 | n19142 ;
  assign n19144 = n4415 | n19143 ;
  assign n19145 = n17919 | n19144 ;
  assign n19146 = ( ~n18709 & n18711 ) | ( ~n18709 & n19145 ) | ( n18711 & n19145 ) ;
  assign n19147 = ( n18709 & n18711 ) | ( n18709 & n19145 ) | ( n18711 & n19145 ) ;
  assign n19148 = ( n18709 & n19146 ) | ( n18709 & ~n19147 ) | ( n19146 & ~n19147 ) ;
  assign n19149 = n3273 & n10326 ;
  assign n19150 = n3270 | n19149 ;
  assign n19151 = ( ~n10332 & n19149 ) | ( ~n10332 & n19150 ) | ( n19149 & n19150 ) ;
  assign n19152 = n390 | n19151 ;
  assign n19153 = ( ~n10383 & n19151 ) | ( ~n10383 & n19152 ) | ( n19151 & n19152 ) ;
  assign n19154 = n3274 & n10329 ;
  assign n19155 = n19153 | n19154 ;
  assign n19156 = ( ~n19125 & n19148 ) | ( ~n19125 & n19155 ) | ( n19148 & n19155 ) ;
  assign n19157 = ( n19125 & n19148 ) | ( n19125 & n19155 ) | ( n19148 & n19155 ) ;
  assign n19158 = ( n19125 & n19156 ) | ( n19125 & ~n19157 ) | ( n19156 & ~n19157 ) ;
  assign n19159 = n4200 & ~n13473 ;
  assign n19160 = n4215 | n19159 ;
  assign n19161 = ( n13475 & n19159 ) | ( n13475 & n19160 ) | ( n19159 & n19160 ) ;
  assign n19162 = n2083 & ~n13280 ;
  assign n19163 = n19161 | n19162 ;
  assign n19164 = x26 & n19163 ;
  assign n19165 = n4203 & n13671 ;
  assign n19166 = ( ~x26 & n19163 ) | ( ~x26 & n19165 ) | ( n19163 & n19165 ) ;
  assign n19167 = x26 & ~n19165 ;
  assign n19168 = ( ~n19164 & n19166 ) | ( ~n19164 & n19167 ) | ( n19166 & n19167 ) ;
  assign n19169 = ( n18714 & n19158 ) | ( n18714 & n19168 ) | ( n19158 & n19168 ) ;
  assign n19170 = ( n18714 & ~n19158 ) | ( n18714 & n19168 ) | ( ~n19158 & n19168 ) ;
  assign n19171 = ( n19158 & ~n19169 ) | ( n19158 & n19170 ) | ( ~n19169 & n19170 ) ;
  assign n19172 = ( ~n18716 & n18720 ) | ( ~n18716 & n19171 ) | ( n18720 & n19171 ) ;
  assign n19173 = ( n18716 & n18720 ) | ( n18716 & n19171 ) | ( n18720 & n19171 ) ;
  assign n19174 = ( n18716 & n19172 ) | ( n18716 & ~n19173 ) | ( n19172 & ~n19173 ) ;
  assign n19175 = ( n18726 & ~n18729 ) | ( n18726 & n19174 ) | ( ~n18729 & n19174 ) ;
  assign n19176 = ( n18726 & n18729 ) | ( n18726 & n19174 ) | ( n18729 & n19174 ) ;
  assign n19177 = ( n18729 & n19175 ) | ( n18729 & ~n19176 ) | ( n19175 & ~n19176 ) ;
  assign n19178 = n18664 & ~n18730 ;
  assign n19179 = ~n19177 & n19178 ;
  assign n19180 = n18734 | n19177 ;
  assign n19181 = ( n18734 & n19177 ) | ( n18734 & n19178 ) | ( n19177 & n19178 ) ;
  assign n19182 = ( n19179 & n19180 ) | ( n19179 & ~n19181 ) | ( n19180 & ~n19181 ) ;
  assign n19183 = n9592 & ~n19182 ;
  assign n19184 = n9593 & n19177 ;
  assign n19185 = n41 & n18730 ;
  assign n19186 = n19184 | n19185 ;
  assign n19187 = x2 | n19186 ;
  assign n19188 = ( ~n19183 & n19186 ) | ( ~n19183 & n19187 ) | ( n19186 & n19187 ) ;
  assign n19189 = n9591 & ~n19182 ;
  assign n19190 = n19188 | n19189 ;
  assign n19191 = n9600 & ~n18362 ;
  assign n19192 = ( x2 & n19186 ) | ( x2 & n19191 ) | ( n19186 & n19191 ) ;
  assign n19193 = n19190 & ~n19192 ;
  assign n19194 = ( n19113 & n19115 ) | ( n19113 & n19193 ) | ( n19115 & n19193 ) ;
  assign n19195 = n2083 | n4215 ;
  assign n19196 = ( n4215 & ~n13473 ) | ( n4215 & n19195 ) | ( ~n13473 & n19195 ) ;
  assign n19197 = n4200 | n19196 ;
  assign n19198 = ( n13475 & n19196 ) | ( n13475 & n19197 ) | ( n19196 & n19197 ) ;
  assign n19199 = x26 & n19198 ;
  assign n19200 = n4202 & n13477 ;
  assign n19201 = x26 & ~n19200 ;
  assign n19202 = ( ~x26 & n19198 ) | ( ~x26 & n19200 ) | ( n19198 & n19200 ) ;
  assign n19203 = ( ~n19199 & n19201 ) | ( ~n19199 & n19202 ) | ( n19201 & n19202 ) ;
  assign n19204 = n3541 & ~n13285 ;
  assign n19205 = x29 & n19204 ;
  assign n19206 = n3536 & n10214 ;
  assign n19207 = n4039 | n19206 ;
  assign n19208 = ( ~n13280 & n19206 ) | ( ~n13280 & n19207 ) | ( n19206 & n19207 ) ;
  assign n19209 = n3501 & ~n10235 ;
  assign n19210 = n19208 | n19209 ;
  assign n19211 = x29 & ~n19210 ;
  assign n19212 = ( ~x29 & n19204 ) | ( ~x29 & n19210 ) | ( n19204 & n19210 ) ;
  assign n19213 = ( ~n19205 & n19211 ) | ( ~n19205 & n19212 ) | ( n19211 & n19212 ) ;
  assign n19214 = n3270 & ~n10237 ;
  assign n19215 = n3274 & ~n10332 ;
  assign n19216 = n3273 & n10329 ;
  assign n19217 = n19215 | n19216 ;
  assign n19218 = n19214 | n19217 ;
  assign n19219 = n390 & n12756 ;
  assign n19220 = n19218 | n19219 ;
  assign n19221 = n12888 | n15507 ;
  assign n19222 = n17289 | n19221 ;
  assign n19223 = n2801 | n3992 ;
  assign n19224 = n3786 | n14457 ;
  assign n19225 = n19223 | n19224 ;
  assign n19226 = n6131 | n19225 ;
  assign n19227 = n55 | n3454 ;
  assign n19228 = n766 | n19227 ;
  assign n19229 = n865 | n19228 ;
  assign n19230 = n421 | n19229 ;
  assign n19231 = n19226 | n19230 ;
  assign n19232 = n4767 | n19231 ;
  assign n19233 = n19222 | n19232 ;
  assign n19234 = ( ~n18720 & n19145 ) | ( ~n18720 & n19233 ) | ( n19145 & n19233 ) ;
  assign n19235 = ( n18720 & n19145 ) | ( n18720 & n19233 ) | ( n19145 & n19233 ) ;
  assign n19236 = ( n18720 & n19234 ) | ( n18720 & ~n19235 ) | ( n19234 & ~n19235 ) ;
  assign n19237 = ( n19146 & ~n19220 ) | ( n19146 & n19236 ) | ( ~n19220 & n19236 ) ;
  assign n19238 = ( n19146 & n19220 ) | ( n19146 & ~n19236 ) | ( n19220 & ~n19236 ) ;
  assign n19239 = ( ~n19146 & n19237 ) | ( ~n19146 & n19238 ) | ( n19237 & n19238 ) ;
  assign n19240 = ( n19157 & n19213 ) | ( n19157 & n19239 ) | ( n19213 & n19239 ) ;
  assign n19241 = ( ~n19157 & n19213 ) | ( ~n19157 & n19239 ) | ( n19213 & n19239 ) ;
  assign n19242 = ( n19157 & ~n19240 ) | ( n19157 & n19241 ) | ( ~n19240 & n19241 ) ;
  assign n19243 = ( ~n19169 & n19203 ) | ( ~n19169 & n19242 ) | ( n19203 & n19242 ) ;
  assign n19244 = ( n19169 & n19203 ) | ( n19169 & n19242 ) | ( n19203 & n19242 ) ;
  assign n19245 = ( n19169 & n19243 ) | ( n19169 & ~n19244 ) | ( n19243 & ~n19244 ) ;
  assign n19246 = ( n19173 & ~n19176 ) | ( n19173 & n19245 ) | ( ~n19176 & n19245 ) ;
  assign n19247 = ( n19173 & n19176 ) | ( n19173 & n19245 ) | ( n19176 & n19245 ) ;
  assign n19248 = ( n19176 & n19246 ) | ( n19176 & ~n19247 ) | ( n19246 & ~n19247 ) ;
  assign n19249 = n19177 & ~n19178 ;
  assign n19250 = n19248 & n19249 ;
  assign n19251 = n19180 & n19248 ;
  assign n19252 = ( n19180 & n19248 ) | ( n19180 & ~n19249 ) | ( n19248 & ~n19249 ) ;
  assign n19253 = ( n19250 & ~n19251 ) | ( n19250 & n19252 ) | ( ~n19251 & n19252 ) ;
  assign n19254 = n9593 & n19248 ;
  assign n19255 = n9592 | n19254 ;
  assign n19256 = ( n19253 & n19254 ) | ( n19253 & n19255 ) | ( n19254 & n19255 ) ;
  assign n19257 = n41 & n19177 ;
  assign n19258 = ( x2 & ~n19256 ) | ( x2 & n19257 ) | ( ~n19256 & n19257 ) ;
  assign n19259 = ~x2 & n19256 ;
  assign n19260 = n9600 & n18730 ;
  assign n19261 = ( x2 & n19257 ) | ( x2 & n19260 ) | ( n19257 & n19260 ) ;
  assign n19262 = ( n19258 & n19259 ) | ( n19258 & ~n19261 ) | ( n19259 & ~n19261 ) ;
  assign n19263 = ( n18273 & ~n18377 ) | ( n18273 & n18529 ) | ( ~n18377 & n18529 ) ;
  assign n19264 = ( ~n18273 & n18530 ) | ( ~n18273 & n19263 ) | ( n18530 & n19263 ) ;
  assign n19265 = ( n19194 & n19262 ) | ( n19194 & ~n19264 ) | ( n19262 & ~n19264 ) ;
  assign n19266 = n101 & ~n13475 ;
  assign n19267 = ( x23 & ~x24 ) | ( x23 & x25 ) | ( ~x24 & x25 ) ;
  assign n19268 = ( x24 & ~x26 ) | ( x24 & n19267 ) | ( ~x26 & n19267 ) ;
  assign n19269 = ~n19266 & n19268 ;
  assign n19270 = n187 & ~n13475 ;
  assign n19271 = n19269 | n19270 ;
  assign n19272 = n3501 & ~n13280 ;
  assign n19273 = x29 & n19272 ;
  assign n19274 = n4039 & ~n13473 ;
  assign n19275 = n3536 & ~n10235 ;
  assign n19276 = n19274 | n19275 ;
  assign n19277 = n3541 | n19276 ;
  assign n19278 = ( ~n13480 & n19276 ) | ( ~n13480 & n19277 ) | ( n19276 & n19277 ) ;
  assign n19279 = x29 & ~n19278 ;
  assign n19280 = ( ~x29 & n19272 ) | ( ~x29 & n19278 ) | ( n19272 & n19278 ) ;
  assign n19281 = ( ~n19273 & n19279 ) | ( ~n19273 & n19280 ) | ( n19279 & n19280 ) ;
  assign n19282 = n285 | n1041 ;
  assign n19283 = n268 | n19282 ;
  assign n19284 = n317 | n3448 ;
  assign n19285 = n19283 | n19284 ;
  assign n19286 = n1437 | n2357 ;
  assign n19287 = n19285 | n19286 ;
  assign n19288 = n6034 | n19287 ;
  assign n19289 = n398 | n565 ;
  assign n19290 = n976 | n2658 ;
  assign n19291 = n19289 | n19290 ;
  assign n19292 = n1846 | n19291 ;
  assign n19293 = n19288 | n19292 ;
  assign n19294 = n561 | n19293 ;
  assign n19295 = n654 & ~n19294 ;
  assign n19296 = ~n10189 & n19295 ;
  assign n19297 = n3273 & ~n10332 ;
  assign n19298 = n3270 | n19297 ;
  assign n19299 = ( n10214 & n19297 ) | ( n10214 & n19298 ) | ( n19297 & n19298 ) ;
  assign n19300 = n390 | n19299 ;
  assign n19301 = ( n12953 & n19299 ) | ( n12953 & n19300 ) | ( n19299 & n19300 ) ;
  assign n19302 = n3274 & ~n10237 ;
  assign n19303 = n19301 | n19302 ;
  assign n19304 = ( n19234 & ~n19296 ) | ( n19234 & n19303 ) | ( ~n19296 & n19303 ) ;
  assign n19305 = ( n19234 & n19296 ) | ( n19234 & n19303 ) | ( n19296 & n19303 ) ;
  assign n19306 = ( n19296 & n19304 ) | ( n19296 & ~n19305 ) | ( n19304 & ~n19305 ) ;
  assign n19307 = ( ~n19237 & n19281 ) | ( ~n19237 & n19306 ) | ( n19281 & n19306 ) ;
  assign n19308 = ( n19237 & n19281 ) | ( n19237 & n19306 ) | ( n19281 & n19306 ) ;
  assign n19309 = ( n19237 & n19307 ) | ( n19237 & ~n19308 ) | ( n19307 & ~n19308 ) ;
  assign n19310 = ( ~n19240 & n19271 ) | ( ~n19240 & n19309 ) | ( n19271 & n19309 ) ;
  assign n19311 = ( n19240 & n19271 ) | ( n19240 & ~n19309 ) | ( n19271 & ~n19309 ) ;
  assign n19312 = ( ~n19271 & n19310 ) | ( ~n19271 & n19311 ) | ( n19310 & n19311 ) ;
  assign n19313 = ( ~n19244 & n19247 ) | ( ~n19244 & n19312 ) | ( n19247 & n19312 ) ;
  assign n19314 = ( n19244 & n19247 ) | ( n19244 & ~n19312 ) | ( n19247 & ~n19312 ) ;
  assign n19315 = ( ~n19247 & n19313 ) | ( ~n19247 & n19314 ) | ( n19313 & n19314 ) ;
  assign n19316 = n19251 & n19315 ;
  assign n19317 = n19248 | n19249 ;
  assign n19318 = ( ~n19251 & n19315 ) | ( ~n19251 & n19317 ) | ( n19315 & n19317 ) ;
  assign n19319 = n19315 & n19317 ;
  assign n19320 = ( n19316 & n19318 ) | ( n19316 & ~n19319 ) | ( n19318 & ~n19319 ) ;
  assign n19321 = n9593 & ~n19315 ;
  assign n19322 = n9592 | n19321 ;
  assign n19323 = ( ~n19320 & n19321 ) | ( ~n19320 & n19322 ) | ( n19321 & n19322 ) ;
  assign n19324 = n41 & n19248 ;
  assign n19325 = ( x2 & ~n19323 ) | ( x2 & n19324 ) | ( ~n19323 & n19324 ) ;
  assign n19326 = ~x2 & n19323 ;
  assign n19327 = n9600 & n19177 ;
  assign n19328 = ( x2 & n19324 ) | ( x2 & n19327 ) | ( n19324 & n19327 ) ;
  assign n19329 = ( n19325 & n19326 ) | ( n19325 & ~n19328 ) | ( n19326 & ~n19328 ) ;
  assign n19330 = ( ~n18748 & n19265 ) | ( ~n18748 & n19329 ) | ( n19265 & n19329 ) ;
  assign n19331 = n3273 & ~n10237 ;
  assign n19332 = n3270 | n19331 ;
  assign n19333 = ( ~n10235 & n19331 ) | ( ~n10235 & n19332 ) | ( n19331 & n19332 ) ;
  assign n19334 = n390 | n19333 ;
  assign n19335 = ( n10371 & n19333 ) | ( n10371 & n19334 ) | ( n19333 & n19334 ) ;
  assign n19336 = n3274 & n10214 ;
  assign n19337 = n19335 | n19336 ;
  assign n19338 = n751 | n977 ;
  assign n19339 = n677 | n19338 ;
  assign n19340 = n2201 | n12866 ;
  assign n19341 = n19339 | n19340 ;
  assign n19342 = n1631 | n19341 ;
  assign n19343 = n3596 | n19342 ;
  assign n19344 = n1248 | n2260 ;
  assign n19345 = n19343 | n19344 ;
  assign n19346 = n514 | n19345 ;
  assign n19347 = ( n19295 & n19337 ) | ( n19295 & n19346 ) | ( n19337 & n19346 ) ;
  assign n19348 = ( ~n19295 & n19337 ) | ( ~n19295 & n19346 ) | ( n19337 & n19346 ) ;
  assign n19349 = ( n19295 & ~n19347 ) | ( n19295 & n19348 ) | ( ~n19347 & n19348 ) ;
  assign n19350 = ( n19305 & ~n19307 ) | ( n19305 & n19349 ) | ( ~n19307 & n19349 ) ;
  assign n19351 = ( n19305 & n19307 ) | ( n19305 & n19349 ) | ( n19307 & n19349 ) ;
  assign n19352 = ( n19307 & n19350 ) | ( n19307 & ~n19351 ) | ( n19350 & ~n19351 ) ;
  assign n19353 = n3536 & ~n13280 ;
  assign n19354 = n4039 | n19353 ;
  assign n19355 = ( n13475 & n19353 ) | ( n13475 & n19354 ) | ( n19353 & n19354 ) ;
  assign n19356 = n3501 & ~n13473 ;
  assign n19357 = n19355 | n19356 ;
  assign n19358 = x29 & n19357 ;
  assign n19359 = n3541 & n13671 ;
  assign n19360 = ( ~x29 & n19357 ) | ( ~x29 & n19359 ) | ( n19357 & n19359 ) ;
  assign n19361 = x29 & ~n19359 ;
  assign n19362 = ( ~n19358 & n19360 ) | ( ~n19358 & n19361 ) | ( n19360 & n19361 ) ;
  assign n19363 = ( ~n19268 & n19352 ) | ( ~n19268 & n19362 ) | ( n19352 & n19362 ) ;
  assign n19364 = ( n19268 & n19352 ) | ( n19268 & n19362 ) | ( n19352 & n19362 ) ;
  assign n19365 = ( n19268 & n19363 ) | ( n19268 & ~n19364 ) | ( n19363 & ~n19364 ) ;
  assign n19366 = ( n19311 & n19314 ) | ( n19311 & n19365 ) | ( n19314 & n19365 ) ;
  assign n19367 = ( n19311 & ~n19314 ) | ( n19311 & n19365 ) | ( ~n19314 & n19365 ) ;
  assign n19368 = ( n19314 & ~n19366 ) | ( n19314 & n19367 ) | ( ~n19366 & n19367 ) ;
  assign n19369 = ~n19315 & n19317 ;
  assign n19370 = n19368 & n19369 ;
  assign n19371 = ~n19251 & n19315 ;
  assign n19372 = n19368 & ~n19371 ;
  assign n19373 = ( ~n19368 & n19369 ) | ( ~n19368 & n19371 ) | ( n19369 & n19371 ) ;
  assign n19374 = ( ~n19370 & n19372 ) | ( ~n19370 & n19373 ) | ( n19372 & n19373 ) ;
  assign n19375 = n9592 & ~n19374 ;
  assign n19376 = n9593 & n19368 ;
  assign n19377 = n41 & ~n19315 ;
  assign n19378 = n19376 | n19377 ;
  assign n19379 = x2 | n19378 ;
  assign n19380 = ( ~n19375 & n19378 ) | ( ~n19375 & n19379 ) | ( n19378 & n19379 ) ;
  assign n19381 = n9591 & ~n19374 ;
  assign n19382 = n19380 | n19381 ;
  assign n19383 = n9600 & n19248 ;
  assign n19384 = ( x2 & n19378 ) | ( x2 & n19383 ) | ( n19378 & n19383 ) ;
  assign n19385 = n19382 & ~n19384 ;
  assign n19386 = n40 & n19177 ;
  assign n19387 = n8721 & n18730 ;
  assign n19388 = n8340 & ~n18362 ;
  assign n19389 = n19387 | n19388 ;
  assign n19390 = n19386 | n19389 ;
  assign n19391 = x5 & n19390 ;
  assign n19392 = n8341 & ~n19182 ;
  assign n19393 = ( ~x5 & n19390 ) | ( ~x5 & n19392 ) | ( n19390 & n19392 ) ;
  assign n19394 = x5 & ~n19392 ;
  assign n19395 = ( ~n19391 & n19393 ) | ( ~n19391 & n19394 ) | ( n19393 & n19394 ) ;
  assign n19396 = n6796 & n17346 ;
  assign n19397 = x11 & n19396 ;
  assign n19398 = n6567 & ~n17126 ;
  assign n19399 = n6570 | n19398 ;
  assign n19400 = ( ~n17635 & n19398 ) | ( ~n17635 & n19399 ) | ( n19398 & n19399 ) ;
  assign n19401 = n6571 | n19400 ;
  assign n19402 = ( ~n17646 & n19400 ) | ( ~n17646 & n19401 ) | ( n19400 & n19401 ) ;
  assign n19403 = x11 & ~n19402 ;
  assign n19404 = ( ~x11 & n19396 ) | ( ~x11 & n19402 ) | ( n19396 & n19402 ) ;
  assign n19405 = ( ~n19397 & n19403 ) | ( ~n19397 & n19404 ) | ( n19403 & n19404 ) ;
  assign n19406 = n6332 & n16724 ;
  assign n19407 = x14 & n19406 ;
  assign n19408 = n5909 & ~n16531 ;
  assign n19409 = n5914 | n19408 ;
  assign n19410 = ( n16925 & n19408 ) | ( n16925 & n19409 ) | ( n19408 & n19409 ) ;
  assign n19411 = n5915 | n19410 ;
  assign n19412 = ( ~n16936 & n19410 ) | ( ~n16936 & n19411 ) | ( n19410 & n19411 ) ;
  assign n19413 = x14 & ~n19412 ;
  assign n19414 = ( ~x14 & n19406 ) | ( ~x14 & n19412 ) | ( n19406 & n19412 ) ;
  assign n19415 = ( ~n19407 & n19413 ) | ( ~n19407 & n19414 ) | ( n19413 & n19414 ) ;
  assign n19416 = n4637 & n14942 ;
  assign n19417 = x23 & n19416 ;
  assign n19418 = n4584 & ~n14723 ;
  assign n19419 = n4649 | n19418 ;
  assign n19420 = ( ~n15184 & n19418 ) | ( ~n15184 & n19419 ) | ( n19418 & n19419 ) ;
  assign n19421 = n4591 | n19420 ;
  assign n19422 = ( ~n15195 & n19420 ) | ( ~n15195 & n19421 ) | ( n19420 & n19421 ) ;
  assign n19423 = x23 & ~n19422 ;
  assign n19424 = ( ~x23 & n19416 ) | ( ~x23 & n19422 ) | ( n19416 & n19422 ) ;
  assign n19425 = ( ~n19417 & n19423 ) | ( ~n19417 & n19424 ) | ( n19423 & n19424 ) ;
  assign n19426 = n4215 & n14520 ;
  assign n19427 = n4200 & n14352 ;
  assign n19428 = n2083 & n13992 ;
  assign n19429 = n19427 | n19428 ;
  assign n19430 = n19426 | n19429 ;
  assign n19431 = x26 & n19430 ;
  assign n19432 = n4203 & n14531 ;
  assign n19433 = ( ~x26 & n19430 ) | ( ~x26 & n19432 ) | ( n19430 & n19432 ) ;
  assign n19434 = x26 & ~n19432 ;
  assign n19435 = ( ~n19431 & n19433 ) | ( ~n19431 & n19434 ) | ( n19433 & n19434 ) ;
  assign n19436 = n3541 & ~n14130 ;
  assign n19437 = x29 & n19436 ;
  assign n19438 = n3536 & ~n14000 ;
  assign n19439 = n4039 | n19438 ;
  assign n19440 = ( n13996 & n19438 ) | ( n13996 & n19439 ) | ( n19438 & n19439 ) ;
  assign n19441 = n3501 & n13998 ;
  assign n19442 = n19440 | n19441 ;
  assign n19443 = x29 & ~n19442 ;
  assign n19444 = ( ~x29 & n19436 ) | ( ~x29 & n19442 ) | ( n19436 & n19442 ) ;
  assign n19445 = ( ~n19437 & n19443 ) | ( ~n19437 & n19444 ) | ( n19443 & n19444 ) ;
  assign n19446 = n1276 | n3355 ;
  assign n19447 = n581 | n2762 ;
  assign n19448 = n18332 | n19447 ;
  assign n19449 = n19446 | n19448 ;
  assign n19450 = n4137 | n19449 ;
  assign n19451 = n613 | n1081 ;
  assign n19452 = n3623 | n19451 ;
  assign n19453 = n1302 | n2449 ;
  assign n19454 = n19452 | n19453 ;
  assign n19455 = n2177 | n19454 ;
  assign n19456 = n133 | n781 ;
  assign n19457 = n358 | n19456 ;
  assign n19458 = n19455 | n19457 ;
  assign n19459 = n19450 | n19458 ;
  assign n19460 = n5090 | n19459 ;
  assign n19461 = n1553 | n19460 ;
  assign n19462 = n2466 | n19461 ;
  assign n19463 = n3273 & ~n14004 ;
  assign n19464 = n3270 | n19463 ;
  assign n19465 = ( ~n14007 & n19463 ) | ( ~n14007 & n19464 ) | ( n19463 & n19464 ) ;
  assign n19466 = n390 | n19465 ;
  assign n19467 = ( n14066 & n19465 ) | ( n14066 & n19466 ) | ( n19465 & n19466 ) ;
  assign n19468 = n3274 & n14002 ;
  assign n19469 = n19467 | n19468 ;
  assign n19470 = ( n18617 & n19462 ) | ( n18617 & n19469 ) | ( n19462 & n19469 ) ;
  assign n19471 = ( ~n18617 & n19462 ) | ( ~n18617 & n19469 ) | ( n19462 & n19469 ) ;
  assign n19472 = ( n18617 & ~n19470 ) | ( n18617 & n19471 ) | ( ~n19470 & n19471 ) ;
  assign n19473 = ( ~n18621 & n19445 ) | ( ~n18621 & n19472 ) | ( n19445 & n19472 ) ;
  assign n19474 = ( n18621 & n19445 ) | ( n18621 & n19472 ) | ( n19445 & n19472 ) ;
  assign n19475 = ( n18621 & n19473 ) | ( n18621 & ~n19474 ) | ( n19473 & ~n19474 ) ;
  assign n19476 = ( n18624 & n19435 ) | ( n18624 & n19475 ) | ( n19435 & n19475 ) ;
  assign n19477 = ( ~n18624 & n19435 ) | ( ~n18624 & n19475 ) | ( n19435 & n19475 ) ;
  assign n19478 = ( n18624 & ~n19476 ) | ( n18624 & n19477 ) | ( ~n19476 & n19477 ) ;
  assign n19479 = ( ~n18626 & n19425 ) | ( ~n18626 & n19478 ) | ( n19425 & n19478 ) ;
  assign n19480 = ( n18626 & n19425 ) | ( n18626 & n19478 ) | ( n19425 & n19478 ) ;
  assign n19481 = ( n18626 & n19479 ) | ( n18626 & ~n19480 ) | ( n19479 & ~n19480 ) ;
  assign n19482 = n5232 & n15561 ;
  assign n19483 = x20 & n19482 ;
  assign n19484 = n4874 & ~n15394 ;
  assign n19485 = n4878 | n19484 ;
  assign n19486 = ( ~n15806 & n19484 ) | ( ~n15806 & n19485 ) | ( n19484 & n19485 ) ;
  assign n19487 = n4879 | n19486 ;
  assign n19488 = ( n15817 & n19486 ) | ( n15817 & n19487 ) | ( n19486 & n19487 ) ;
  assign n19489 = x20 & ~n19488 ;
  assign n19490 = ( ~x20 & n19482 ) | ( ~x20 & n19488 ) | ( n19482 & n19488 ) ;
  assign n19491 = ( ~n19483 & n19489 ) | ( ~n19483 & n19490 ) | ( n19489 & n19490 ) ;
  assign n19492 = ( ~n18629 & n19481 ) | ( ~n18629 & n19491 ) | ( n19481 & n19491 ) ;
  assign n19493 = ( n18629 & n19481 ) | ( n18629 & n19491 ) | ( n19481 & n19491 ) ;
  assign n19494 = ( n18629 & n19492 ) | ( n18629 & ~n19493 ) | ( n19492 & ~n19493 ) ;
  assign n19495 = n5584 & ~n16150 ;
  assign n19496 = x17 & n19495 ;
  assign n19497 = n5413 & ~n15954 ;
  assign n19498 = n5417 | n19497 ;
  assign n19499 = ( ~n16338 & n19497 ) | ( ~n16338 & n19498 ) | ( n19497 & n19498 ) ;
  assign n19500 = n5418 | n19499 ;
  assign n19501 = ( ~n16349 & n19499 ) | ( ~n16349 & n19500 ) | ( n19499 & n19500 ) ;
  assign n19502 = x17 & ~n19501 ;
  assign n19503 = ( ~x17 & n19495 ) | ( ~x17 & n19501 ) | ( n19495 & n19501 ) ;
  assign n19504 = ( ~n19496 & n19502 ) | ( ~n19496 & n19503 ) | ( n19502 & n19503 ) ;
  assign n19505 = ( ~n18633 & n19494 ) | ( ~n18633 & n19504 ) | ( n19494 & n19504 ) ;
  assign n19506 = ( n18633 & n19494 ) | ( n18633 & n19504 ) | ( n19494 & n19504 ) ;
  assign n19507 = ( n18633 & n19505 ) | ( n18633 & ~n19506 ) | ( n19505 & ~n19506 ) ;
  assign n19508 = ( ~n18646 & n19415 ) | ( ~n18646 & n19507 ) | ( n19415 & n19507 ) ;
  assign n19509 = ( n18646 & n19415 ) | ( n18646 & n19507 ) | ( n19415 & n19507 ) ;
  assign n19510 = ( n18646 & n19508 ) | ( n18646 & ~n19509 ) | ( n19508 & ~n19509 ) ;
  assign n19511 = ( ~n18649 & n19405 ) | ( ~n18649 & n19510 ) | ( n19405 & n19510 ) ;
  assign n19512 = ( n18649 & n19405 ) | ( n18649 & n19510 ) | ( n19405 & n19510 ) ;
  assign n19513 = ( n18649 & n19511 ) | ( n18649 & ~n19512 ) | ( n19511 & ~n19512 ) ;
  assign n19514 = n7644 & ~n17963 ;
  assign n19515 = x8 & n19514 ;
  assign n19516 = n7341 & n17742 ;
  assign n19517 = n7345 | n19516 ;
  assign n19518 = ( ~n18258 & n19516 ) | ( ~n18258 & n19517 ) | ( n19516 & n19517 ) ;
  assign n19519 = n7346 | n19518 ;
  assign n19520 = ( n18268 & n19518 ) | ( n18268 & n19519 ) | ( n19518 & n19519 ) ;
  assign n19521 = x8 & ~n19520 ;
  assign n19522 = ( ~x8 & n19514 ) | ( ~x8 & n19520 ) | ( n19514 & n19520 ) ;
  assign n19523 = ( ~n19515 & n19521 ) | ( ~n19515 & n19522 ) | ( n19521 & n19522 ) ;
  assign n19524 = ( ~n18661 & n19513 ) | ( ~n18661 & n19523 ) | ( n19513 & n19523 ) ;
  assign n19525 = ( n18661 & n19513 ) | ( n18661 & n19523 ) | ( n19513 & n19523 ) ;
  assign n19526 = ( n18661 & n19524 ) | ( n18661 & ~n19525 ) | ( n19524 & ~n19525 ) ;
  assign n19527 = ( ~n18746 & n19395 ) | ( ~n18746 & n19526 ) | ( n19395 & n19526 ) ;
  assign n19528 = ( n18746 & n19395 ) | ( n18746 & n19526 ) | ( n19395 & n19526 ) ;
  assign n19529 = ( n18746 & n19527 ) | ( n18746 & ~n19528 ) | ( n19527 & ~n19528 ) ;
  assign n19530 = ( n19330 & n19385 ) | ( n19330 & n19529 ) | ( n19385 & n19529 ) ;
  assign n19531 = n40 & n19248 ;
  assign n19532 = n8721 & n19177 ;
  assign n19533 = n8340 & n18730 ;
  assign n19534 = n19532 | n19533 ;
  assign n19535 = n19531 | n19534 ;
  assign n19536 = x5 & n19535 ;
  assign n19537 = n8341 & n19253 ;
  assign n19538 = ( ~x5 & n19535 ) | ( ~x5 & n19537 ) | ( n19535 & n19537 ) ;
  assign n19539 = x5 & ~n19537 ;
  assign n19540 = ( ~n19536 & n19538 ) | ( ~n19536 & n19539 ) | ( n19538 & n19539 ) ;
  assign n19541 = n7346 & ~n18373 ;
  assign n19542 = x8 & n19541 ;
  assign n19543 = n7341 & ~n17963 ;
  assign n19544 = n7345 | n19543 ;
  assign n19545 = ( ~n18362 & n19543 ) | ( ~n18362 & n19544 ) | ( n19543 & n19544 ) ;
  assign n19546 = n7644 & ~n18258 ;
  assign n19547 = n19545 | n19546 ;
  assign n19548 = x8 & ~n19547 ;
  assign n19549 = ( ~x8 & n19541 ) | ( ~x8 & n19547 ) | ( n19541 & n19547 ) ;
  assign n19550 = ( ~n19542 & n19548 ) | ( ~n19542 & n19549 ) | ( n19548 & n19549 ) ;
  assign n19551 = n6570 & n17742 ;
  assign n19552 = x11 & n19551 ;
  assign n19553 = n6796 & ~n17635 ;
  assign n19554 = n6567 & n17346 ;
  assign n19555 = n19553 | n19554 ;
  assign n19556 = n6571 | n19555 ;
  assign n19557 = ( ~n17749 & n19555 ) | ( ~n17749 & n19556 ) | ( n19555 & n19556 ) ;
  assign n19558 = x11 & ~n19557 ;
  assign n19559 = ( ~x11 & n19551 ) | ( ~x11 & n19557 ) | ( n19551 & n19557 ) ;
  assign n19560 = ( ~n19552 & n19558 ) | ( ~n19552 & n19559 ) | ( n19558 & n19559 ) ;
  assign n19561 = n5915 & ~n17139 ;
  assign n19562 = x14 & n19561 ;
  assign n19563 = n5909 & n16724 ;
  assign n19564 = n5914 | n19563 ;
  assign n19565 = ( ~n17126 & n19563 ) | ( ~n17126 & n19564 ) | ( n19563 & n19564 ) ;
  assign n19566 = n6332 & n16925 ;
  assign n19567 = n19565 | n19566 ;
  assign n19568 = x14 & ~n19567 ;
  assign n19569 = ( ~x14 & n19561 ) | ( ~x14 & n19567 ) | ( n19561 & n19567 ) ;
  assign n19570 = ( ~n19562 & n19568 ) | ( ~n19562 & n19569 ) | ( n19568 & n19569 ) ;
  assign n19571 = n5584 & ~n16338 ;
  assign n19572 = x17 & n19571 ;
  assign n19573 = n5413 & ~n16150 ;
  assign n19574 = n5417 | n19573 ;
  assign n19575 = ( ~n16531 & n19573 ) | ( ~n16531 & n19574 ) | ( n19573 & n19574 ) ;
  assign n19576 = n5418 | n19575 ;
  assign n19577 = ( ~n16542 & n19575 ) | ( ~n16542 & n19576 ) | ( n19575 & n19576 ) ;
  assign n19578 = x17 & ~n19577 ;
  assign n19579 = ( ~x17 & n19571 ) | ( ~x17 & n19577 ) | ( n19571 & n19577 ) ;
  assign n19580 = ( ~n19572 & n19578 ) | ( ~n19572 & n19579 ) | ( n19578 & n19579 ) ;
  assign n19581 = n5232 & ~n15806 ;
  assign n19582 = x20 & n19581 ;
  assign n19583 = n4874 & n15561 ;
  assign n19584 = n4878 | n19583 ;
  assign n19585 = ( ~n15954 & n19583 ) | ( ~n15954 & n19584 ) | ( n19583 & n19584 ) ;
  assign n19586 = n4879 | n19585 ;
  assign n19587 = ( ~n15965 & n19585 ) | ( ~n15965 & n19586 ) | ( n19585 & n19586 ) ;
  assign n19588 = x20 & ~n19587 ;
  assign n19589 = ( ~x20 & n19581 ) | ( ~x20 & n19587 ) | ( n19581 & n19587 ) ;
  assign n19590 = ( ~n19582 & n19588 ) | ( ~n19582 & n19589 ) | ( n19588 & n19589 ) ;
  assign n19591 = n4637 & ~n15184 ;
  assign n19592 = x23 & n19591 ;
  assign n19593 = n4584 & n14942 ;
  assign n19594 = n4649 | n19593 ;
  assign n19595 = ( ~n15394 & n19593 ) | ( ~n15394 & n19594 ) | ( n19593 & n19594 ) ;
  assign n19596 = n4591 | n19595 ;
  assign n19597 = ( n15405 & n19595 ) | ( n15405 & n19596 ) | ( n19595 & n19596 ) ;
  assign n19598 = x23 & ~n19597 ;
  assign n19599 = ( ~x23 & n19591 ) | ( ~x23 & n19597 ) | ( n19591 & n19597 ) ;
  assign n19600 = ( ~n19592 & n19598 ) | ( ~n19592 & n19599 ) | ( n19598 & n19599 ) ;
  assign n19601 = n4039 & n13992 ;
  assign n19602 = x29 & n19601 ;
  assign n19603 = n3501 & n13996 ;
  assign n19604 = n3536 & n13998 ;
  assign n19605 = n19603 | n19604 ;
  assign n19606 = n3541 | n19605 ;
  assign n19607 = ( n14024 & n19605 ) | ( n14024 & n19606 ) | ( n19605 & n19606 ) ;
  assign n19608 = x29 & ~n19607 ;
  assign n19609 = ( ~x29 & n19601 ) | ( ~x29 & n19607 ) | ( n19601 & n19607 ) ;
  assign n19610 = ( ~n19602 & n19608 ) | ( ~n19602 & n19609 ) | ( n19608 & n19609 ) ;
  assign n19611 = n3273 & n14002 ;
  assign n19612 = n3270 | n19611 ;
  assign n19613 = ( ~n14000 & n19611 ) | ( ~n14000 & n19612 ) | ( n19611 & n19612 ) ;
  assign n19614 = n390 | n19613 ;
  assign n19615 = ( ~n14042 & n19613 ) | ( ~n14042 & n19614 ) | ( n19613 & n19614 ) ;
  assign n19616 = n3274 & ~n14007 ;
  assign n19617 = n19615 | n19616 ;
  assign n19618 = n17909 | n19132 ;
  assign n19619 = n586 | n1094 ;
  assign n19620 = n589 | n712 ;
  assign n19621 = n19619 | n19620 ;
  assign n19622 = n5466 | n19621 ;
  assign n19623 = n12668 | n19622 ;
  assign n19624 = n404 | n611 ;
  assign n19625 = n339 | n19624 ;
  assign n19626 = n19623 | n19625 ;
  assign n19627 = n759 | n17940 ;
  assign n19628 = n19626 | n19627 ;
  assign n19629 = n19618 | n19628 ;
  assign n19630 = n13403 & ~n19629 ;
  assign n19631 = ( n19470 & n19617 ) | ( n19470 & ~n19630 ) | ( n19617 & ~n19630 ) ;
  assign n19632 = ( n19470 & ~n19617 ) | ( n19470 & n19630 ) | ( ~n19617 & n19630 ) ;
  assign n19633 = ( ~n19470 & n19631 ) | ( ~n19470 & n19632 ) | ( n19631 & n19632 ) ;
  assign n19634 = ( n19474 & n19610 ) | ( n19474 & ~n19633 ) | ( n19610 & ~n19633 ) ;
  assign n19635 = ( n19474 & ~n19610 ) | ( n19474 & n19633 ) | ( ~n19610 & n19633 ) ;
  assign n19636 = ( ~n19474 & n19634 ) | ( ~n19474 & n19635 ) | ( n19634 & n19635 ) ;
  assign n19637 = n4215 & ~n14723 ;
  assign n19638 = n4200 & n14520 ;
  assign n19639 = n2083 & n14352 ;
  assign n19640 = n19638 | n19639 ;
  assign n19641 = n19637 | n19640 ;
  assign n19642 = x26 & n19641 ;
  assign n19643 = n4203 & ~n14734 ;
  assign n19644 = ( ~x26 & n19641 ) | ( ~x26 & n19643 ) | ( n19641 & n19643 ) ;
  assign n19645 = x26 & ~n19643 ;
  assign n19646 = ( ~n19642 & n19644 ) | ( ~n19642 & n19645 ) | ( n19644 & n19645 ) ;
  assign n19647 = ( n19476 & n19636 ) | ( n19476 & n19646 ) | ( n19636 & n19646 ) ;
  assign n19648 = ( n19476 & ~n19636 ) | ( n19476 & n19646 ) | ( ~n19636 & n19646 ) ;
  assign n19649 = ( n19636 & ~n19647 ) | ( n19636 & n19648 ) | ( ~n19647 & n19648 ) ;
  assign n19650 = ( n19480 & ~n19600 ) | ( n19480 & n19649 ) | ( ~n19600 & n19649 ) ;
  assign n19651 = ( n19480 & n19600 ) | ( n19480 & ~n19649 ) | ( n19600 & ~n19649 ) ;
  assign n19652 = ( ~n19480 & n19650 ) | ( ~n19480 & n19651 ) | ( n19650 & n19651 ) ;
  assign n19653 = ( n19493 & ~n19590 ) | ( n19493 & n19652 ) | ( ~n19590 & n19652 ) ;
  assign n19654 = ( n19493 & n19590 ) | ( n19493 & ~n19652 ) | ( n19590 & ~n19652 ) ;
  assign n19655 = ( ~n19493 & n19653 ) | ( ~n19493 & n19654 ) | ( n19653 & n19654 ) ;
  assign n19656 = ( n19506 & n19580 ) | ( n19506 & ~n19655 ) | ( n19580 & ~n19655 ) ;
  assign n19657 = ( n19506 & ~n19580 ) | ( n19506 & n19655 ) | ( ~n19580 & n19655 ) ;
  assign n19658 = ( ~n19506 & n19656 ) | ( ~n19506 & n19657 ) | ( n19656 & n19657 ) ;
  assign n19659 = ( n19509 & ~n19570 ) | ( n19509 & n19658 ) | ( ~n19570 & n19658 ) ;
  assign n19660 = ( n19509 & n19570 ) | ( n19509 & ~n19658 ) | ( n19570 & ~n19658 ) ;
  assign n19661 = ( ~n19509 & n19659 ) | ( ~n19509 & n19660 ) | ( n19659 & n19660 ) ;
  assign n19662 = ( n19512 & n19560 ) | ( n19512 & ~n19661 ) | ( n19560 & ~n19661 ) ;
  assign n19663 = ( n19512 & ~n19560 ) | ( n19512 & n19661 ) | ( ~n19560 & n19661 ) ;
  assign n19664 = ( ~n19512 & n19662 ) | ( ~n19512 & n19663 ) | ( n19662 & n19663 ) ;
  assign n19665 = ( n19525 & n19550 ) | ( n19525 & ~n19664 ) | ( n19550 & ~n19664 ) ;
  assign n19666 = ( n19525 & ~n19550 ) | ( n19525 & n19664 ) | ( ~n19550 & n19664 ) ;
  assign n19667 = ( ~n19525 & n19665 ) | ( ~n19525 & n19666 ) | ( n19665 & n19666 ) ;
  assign n19668 = ( n19528 & n19540 ) | ( n19528 & ~n19667 ) | ( n19540 & ~n19667 ) ;
  assign n19669 = ( n19528 & ~n19540 ) | ( n19528 & n19667 ) | ( ~n19540 & n19667 ) ;
  assign n19670 = ( ~n19528 & n19668 ) | ( ~n19528 & n19669 ) | ( n19668 & n19669 ) ;
  assign n19671 = n3272 & ~n10235 ;
  assign n19672 = ~n49 & n13280 ;
  assign n19673 = x29 & ~x31 ;
  assign n19674 = n13280 | n19673 ;
  assign n19675 = ( n19671 & ~n19672 ) | ( n19671 & n19674 ) | ( ~n19672 & n19674 ) ;
  assign n19676 = x30 & ~x31 ;
  assign n19677 = n10235 & n19676 ;
  assign n19678 = n19675 & ~n19677 ;
  assign n19679 = n390 & ~n13285 ;
  assign n19680 = n19678 | n19679 ;
  assign n19681 = ~n3416 & n3585 ;
  assign n19682 = ( ~n19268 & n19296 ) | ( ~n19268 & n19681 ) | ( n19296 & n19681 ) ;
  assign n19683 = ( n19268 & n19296 ) | ( n19268 & n19681 ) | ( n19296 & n19681 ) ;
  assign n19684 = ( n19268 & n19682 ) | ( n19268 & ~n19683 ) | ( n19682 & ~n19683 ) ;
  assign n19685 = ( n19347 & n19680 ) | ( n19347 & ~n19684 ) | ( n19680 & ~n19684 ) ;
  assign n19686 = ( n19347 & ~n19680 ) | ( n19347 & n19684 ) | ( ~n19680 & n19684 ) ;
  assign n19687 = ( ~n19347 & n19685 ) | ( ~n19347 & n19686 ) | ( n19685 & n19686 ) ;
  assign n19688 = n3501 | n4039 ;
  assign n19689 = n3536 | n19688 ;
  assign n19690 = ( ~n13473 & n19688 ) | ( ~n13473 & n19689 ) | ( n19688 & n19689 ) ;
  assign n19691 = n3541 | n19690 ;
  assign n19692 = ( n13477 & n19690 ) | ( n13477 & n19691 ) | ( n19690 & n19691 ) ;
  assign n19693 = x29 & ~n19692 ;
  assign n19694 = ~x29 & n19692 ;
  assign n19695 = n19693 | n19694 ;
  assign n19696 = ( n19351 & n19687 ) | ( n19351 & n19695 ) | ( n19687 & n19695 ) ;
  assign n19697 = ( n19351 & ~n19687 ) | ( n19351 & n19695 ) | ( ~n19687 & n19695 ) ;
  assign n19698 = ( n19687 & ~n19696 ) | ( n19687 & n19697 ) | ( ~n19696 & n19697 ) ;
  assign n19699 = ( ~n19364 & n19366 ) | ( ~n19364 & n19698 ) | ( n19366 & n19698 ) ;
  assign n19700 = ( n19364 & n19366 ) | ( n19364 & ~n19698 ) | ( n19366 & ~n19698 ) ;
  assign n19701 = ( ~n19366 & n19699 ) | ( ~n19366 & n19700 ) | ( n19699 & n19700 ) ;
  assign n19702 = n19372 & n19701 ;
  assign n19703 = n19368 | n19369 ;
  assign n19704 = ( ~n19372 & n19701 ) | ( ~n19372 & n19703 ) | ( n19701 & n19703 ) ;
  assign n19705 = n19701 & n19703 ;
  assign n19706 = ( n19702 & n19704 ) | ( n19702 & ~n19705 ) | ( n19704 & ~n19705 ) ;
  assign n19707 = n9592 & ~n19706 ;
  assign n19708 = n9593 & ~n19701 ;
  assign n19709 = n41 & n19368 ;
  assign n19710 = n19708 | n19709 ;
  assign n19711 = x2 | n19710 ;
  assign n19712 = ( ~n19707 & n19710 ) | ( ~n19707 & n19711 ) | ( n19710 & n19711 ) ;
  assign n19713 = n9591 & ~n19706 ;
  assign n19714 = n19712 | n19713 ;
  assign n19715 = n9600 & ~n19315 ;
  assign n19716 = ( x2 & n19710 ) | ( x2 & n19715 ) | ( n19710 & n19715 ) ;
  assign n19717 = n19714 & ~n19716 ;
  assign n19718 = ( n19530 & ~n19670 ) | ( n19530 & n19717 ) | ( ~n19670 & n19717 ) ;
  assign n19719 = ( n19530 & n19670 ) | ( n19530 & ~n19717 ) | ( n19670 & ~n19717 ) ;
  assign n19720 = ( ~n19530 & n19718 ) | ( ~n19530 & n19719 ) | ( n19718 & n19719 ) ;
  assign n19721 = n7644 & ~n18362 ;
  assign n19722 = x8 & n19721 ;
  assign n19723 = n7341 & ~n18258 ;
  assign n19724 = n7345 | n19723 ;
  assign n19725 = ( n18730 & n19723 ) | ( n18730 & n19724 ) | ( n19723 & n19724 ) ;
  assign n19726 = n7346 | n19725 ;
  assign n19727 = ( n18735 & n19725 ) | ( n18735 & n19726 ) | ( n19725 & n19726 ) ;
  assign n19728 = x8 & ~n19727 ;
  assign n19729 = ( ~x8 & n19721 ) | ( ~x8 & n19727 ) | ( n19721 & n19727 ) ;
  assign n19730 = ( ~n19722 & n19728 ) | ( ~n19722 & n19729 ) | ( n19728 & n19729 ) ;
  assign n19731 = n6571 & ~n17976 ;
  assign n19732 = x11 & n19731 ;
  assign n19733 = n6570 & ~n17963 ;
  assign n19734 = n6796 & n17742 ;
  assign n19735 = n6567 & ~n17635 ;
  assign n19736 = n19734 | n19735 ;
  assign n19737 = n19733 | n19736 ;
  assign n19738 = x11 & ~n19737 ;
  assign n19739 = ( ~x11 & n19731 ) | ( ~x11 & n19737 ) | ( n19731 & n19737 ) ;
  assign n19740 = ( ~n19732 & n19738 ) | ( ~n19732 & n19739 ) | ( n19738 & n19739 ) ;
  assign n19741 = n6332 & ~n17126 ;
  assign n19742 = x14 & n19741 ;
  assign n19743 = n5909 & n16925 ;
  assign n19744 = n5914 | n19743 ;
  assign n19745 = ( n17346 & n19743 ) | ( n17346 & n19744 ) | ( n19743 & n19744 ) ;
  assign n19746 = n5915 | n19745 ;
  assign n19747 = ( ~n17356 & n19745 ) | ( ~n17356 & n19746 ) | ( n19745 & n19746 ) ;
  assign n19748 = x14 & ~n19747 ;
  assign n19749 = ( ~x14 & n19741 ) | ( ~x14 & n19747 ) | ( n19741 & n19747 ) ;
  assign n19750 = ( ~n19742 & n19748 ) | ( ~n19742 & n19749 ) | ( n19748 & n19749 ) ;
  assign n19751 = n5584 & ~n16531 ;
  assign n19752 = x17 & n19751 ;
  assign n19753 = n5413 & ~n16338 ;
  assign n19754 = n5417 | n19753 ;
  assign n19755 = ( n16724 & n19753 ) | ( n16724 & n19754 ) | ( n19753 & n19754 ) ;
  assign n19756 = n5418 | n19755 ;
  assign n19757 = ( n16735 & n19755 ) | ( n16735 & n19756 ) | ( n19755 & n19756 ) ;
  assign n19758 = x17 & ~n19757 ;
  assign n19759 = ( ~x17 & n19751 ) | ( ~x17 & n19757 ) | ( n19751 & n19757 ) ;
  assign n19760 = ( ~n19752 & n19758 ) | ( ~n19752 & n19759 ) | ( n19758 & n19759 ) ;
  assign n19761 = n4879 & ~n16161 ;
  assign n19762 = x20 & n19761 ;
  assign n19763 = n4874 & ~n15806 ;
  assign n19764 = n4878 | n19763 ;
  assign n19765 = ( ~n16150 & n19763 ) | ( ~n16150 & n19764 ) | ( n19763 & n19764 ) ;
  assign n19766 = n5232 & ~n15954 ;
  assign n19767 = n19765 | n19766 ;
  assign n19768 = x20 & ~n19767 ;
  assign n19769 = ( ~x20 & n19761 ) | ( ~x20 & n19767 ) | ( n19761 & n19767 ) ;
  assign n19770 = ( ~n19762 & n19768 ) | ( ~n19762 & n19769 ) | ( n19768 & n19769 ) ;
  assign n19771 = n4203 & ~n14953 ;
  assign n19772 = x26 & n19771 ;
  assign n19773 = n4215 & n14942 ;
  assign n19774 = n4200 & ~n14723 ;
  assign n19775 = n2083 & n14520 ;
  assign n19776 = n19774 | n19775 ;
  assign n19777 = n19773 | n19776 ;
  assign n19778 = x26 & ~n19777 ;
  assign n19779 = ( ~x26 & n19771 ) | ( ~x26 & n19777 ) | ( n19771 & n19777 ) ;
  assign n19780 = ( ~n19772 & n19778 ) | ( ~n19772 & n19779 ) | ( n19778 & n19779 ) ;
  assign n19781 = n3501 & n13992 ;
  assign n19782 = x29 & n19781 ;
  assign n19783 = n3536 & n13996 ;
  assign n19784 = n4039 | n19783 ;
  assign n19785 = ( n14352 & n19783 ) | ( n14352 & n19784 ) | ( n19783 & n19784 ) ;
  assign n19786 = n3541 | n19785 ;
  assign n19787 = ( n14363 & n19785 ) | ( n14363 & n19786 ) | ( n19785 & n19786 ) ;
  assign n19788 = x29 & ~n19787 ;
  assign n19789 = ( ~x29 & n19781 ) | ( ~x29 & n19787 ) | ( n19781 & n19787 ) ;
  assign n19790 = ( ~n19782 & n19788 ) | ( ~n19782 & n19789 ) | ( n19788 & n19789 ) ;
  assign n19791 = n3273 & ~n14007 ;
  assign n19792 = n3270 | n19791 ;
  assign n19793 = ( n13998 & n19791 ) | ( n13998 & n19792 ) | ( n19791 & n19792 ) ;
  assign n19794 = n390 | n19793 ;
  assign n19795 = ( n14115 & n19793 ) | ( n14115 & n19794 ) | ( n19793 & n19794 ) ;
  assign n19796 = n3274 & ~n14000 ;
  assign n19797 = n19795 | n19796 ;
  assign n19798 = ~n3977 & n17599 ;
  assign n19799 = n2195 | n17936 ;
  assign n19800 = n358 | n762 ;
  assign n19801 = n19799 | n19800 ;
  assign n19802 = n4805 | n19801 ;
  assign n19803 = n83 | n2386 ;
  assign n19804 = n159 | n3811 ;
  assign n19805 = n1586 | n19804 ;
  assign n19806 = n19803 | n19805 ;
  assign n19807 = n19802 | n19806 ;
  assign n19808 = n19798 & ~n19807 ;
  assign n19809 = ~n4387 & n19808 ;
  assign n19810 = ~n17291 & n19809 ;
  assign n19811 = ( n19631 & ~n19797 ) | ( n19631 & n19810 ) | ( ~n19797 & n19810 ) ;
  assign n19812 = ( n19631 & n19797 ) | ( n19631 & ~n19810 ) | ( n19797 & ~n19810 ) ;
  assign n19813 = ( ~n19631 & n19811 ) | ( ~n19631 & n19812 ) | ( n19811 & n19812 ) ;
  assign n19814 = ( n19634 & ~n19790 ) | ( n19634 & n19813 ) | ( ~n19790 & n19813 ) ;
  assign n19815 = ( n19634 & n19790 ) | ( n19634 & ~n19813 ) | ( n19790 & ~n19813 ) ;
  assign n19816 = ( ~n19634 & n19814 ) | ( ~n19634 & n19815 ) | ( n19814 & n19815 ) ;
  assign n19817 = ( n19648 & n19780 ) | ( n19648 & ~n19816 ) | ( n19780 & ~n19816 ) ;
  assign n19818 = ( n19648 & ~n19780 ) | ( n19648 & n19816 ) | ( ~n19780 & n19816 ) ;
  assign n19819 = ( ~n19648 & n19817 ) | ( ~n19648 & n19818 ) | ( n19817 & n19818 ) ;
  assign n19820 = n4637 & ~n15394 ;
  assign n19821 = x23 & n19820 ;
  assign n19822 = n4584 & ~n15184 ;
  assign n19823 = n4649 | n19822 ;
  assign n19824 = ( n15561 & n19822 ) | ( n15561 & n19823 ) | ( n19822 & n19823 ) ;
  assign n19825 = n4591 | n19824 ;
  assign n19826 = ( n15573 & n19824 ) | ( n15573 & n19825 ) | ( n19824 & n19825 ) ;
  assign n19827 = x23 & ~n19826 ;
  assign n19828 = ( ~x23 & n19820 ) | ( ~x23 & n19826 ) | ( n19820 & n19826 ) ;
  assign n19829 = ( ~n19821 & n19827 ) | ( ~n19821 & n19828 ) | ( n19827 & n19828 ) ;
  assign n19830 = ( n19651 & ~n19819 ) | ( n19651 & n19829 ) | ( ~n19819 & n19829 ) ;
  assign n19831 = ( n19651 & n19819 ) | ( n19651 & ~n19829 ) | ( n19819 & ~n19829 ) ;
  assign n19832 = ( ~n19651 & n19830 ) | ( ~n19651 & n19831 ) | ( n19830 & n19831 ) ;
  assign n19833 = ( n19654 & n19770 ) | ( n19654 & ~n19832 ) | ( n19770 & ~n19832 ) ;
  assign n19834 = ( n19654 & ~n19770 ) | ( n19654 & n19832 ) | ( ~n19770 & n19832 ) ;
  assign n19835 = ( ~n19654 & n19833 ) | ( ~n19654 & n19834 ) | ( n19833 & n19834 ) ;
  assign n19836 = ( n19656 & n19760 ) | ( n19656 & ~n19835 ) | ( n19760 & ~n19835 ) ;
  assign n19837 = ( n19656 & ~n19760 ) | ( n19656 & n19835 ) | ( ~n19760 & n19835 ) ;
  assign n19838 = ( ~n19656 & n19836 ) | ( ~n19656 & n19837 ) | ( n19836 & n19837 ) ;
  assign n19839 = ( n19660 & ~n19750 ) | ( n19660 & n19838 ) | ( ~n19750 & n19838 ) ;
  assign n19840 = ( n19660 & n19750 ) | ( n19660 & ~n19838 ) | ( n19750 & ~n19838 ) ;
  assign n19841 = ( ~n19660 & n19839 ) | ( ~n19660 & n19840 ) | ( n19839 & n19840 ) ;
  assign n19842 = ( n19662 & n19740 ) | ( n19662 & ~n19841 ) | ( n19740 & ~n19841 ) ;
  assign n19843 = ( n19662 & ~n19740 ) | ( n19662 & n19841 ) | ( ~n19740 & n19841 ) ;
  assign n19844 = ( ~n19662 & n19842 ) | ( ~n19662 & n19843 ) | ( n19842 & n19843 ) ;
  assign n19845 = ( n19665 & ~n19730 ) | ( n19665 & n19844 ) | ( ~n19730 & n19844 ) ;
  assign n19846 = ( n19665 & n19730 ) | ( n19665 & ~n19844 ) | ( n19730 & ~n19844 ) ;
  assign n19847 = ( ~n19665 & n19845 ) | ( ~n19665 & n19846 ) | ( n19845 & n19846 ) ;
  assign n19848 = n40 & ~n19315 ;
  assign n19849 = n8721 & n19248 ;
  assign n19850 = n8340 & n19177 ;
  assign n19851 = n19849 | n19850 ;
  assign n19852 = n19848 | n19851 ;
  assign n19853 = x5 & n19852 ;
  assign n19854 = n8341 & ~n19320 ;
  assign n19855 = ( ~x5 & n19852 ) | ( ~x5 & n19854 ) | ( n19852 & n19854 ) ;
  assign n19856 = x5 & ~n19854 ;
  assign n19857 = ( ~n19853 & n19855 ) | ( ~n19853 & n19856 ) | ( n19855 & n19856 ) ;
  assign n19858 = ( n19668 & n19847 ) | ( n19668 & ~n19857 ) | ( n19847 & ~n19857 ) ;
  assign n19859 = ( n19668 & ~n19847 ) | ( n19668 & n19857 ) | ( ~n19847 & n19857 ) ;
  assign n19860 = ( ~n19668 & n19858 ) | ( ~n19668 & n19859 ) | ( n19858 & n19859 ) ;
  assign n19861 = n41 & ~n19701 ;
  assign n19862 = x2 & n19861 ;
  assign n19863 = ( x26 & ~x27 ) | ( x26 & x28 ) | ( ~x27 & x28 ) ;
  assign n19864 = ( x27 & ~x29 ) | ( x27 & n19863 ) | ( ~x29 & n19863 ) ;
  assign n19865 = n3414 | n3513 ;
  assign n19866 = n3554 | n19865 ;
  assign n19867 = n3270 & ~n13473 ;
  assign n19868 = n3274 & ~n13280 ;
  assign n19869 = n19867 | n19868 ;
  assign n19870 = n390 | n19869 ;
  assign n19871 = ( ~n13480 & n19869 ) | ( ~n13480 & n19870 ) | ( n19869 & n19870 ) ;
  assign n19872 = n3273 & n13280 ;
  assign n19873 = n19871 | n19872 ;
  assign n19874 = ( n19683 & n19866 ) | ( n19683 & n19873 ) | ( n19866 & n19873 ) ;
  assign n19875 = ( n19683 & ~n19866 ) | ( n19683 & n19873 ) | ( ~n19866 & n19873 ) ;
  assign n19876 = ( n19866 & ~n19874 ) | ( n19866 & n19875 ) | ( ~n19874 & n19875 ) ;
  assign n19877 = ( ~n19685 & n19864 ) | ( ~n19685 & n19876 ) | ( n19864 & n19876 ) ;
  assign n19878 = ( n19685 & n19864 ) | ( n19685 & n19876 ) | ( n19864 & n19876 ) ;
  assign n19879 = ( n19685 & n19877 ) | ( n19685 & ~n19878 ) | ( n19877 & ~n19878 ) ;
  assign n19880 = ( n19697 & ~n19700 ) | ( n19697 & n19879 ) | ( ~n19700 & n19879 ) ;
  assign n19881 = ( n19697 & n19700 ) | ( n19697 & n19879 ) | ( n19700 & n19879 ) ;
  assign n19882 = ( n19700 & n19880 ) | ( n19700 & ~n19881 ) | ( n19880 & ~n19881 ) ;
  assign n19883 = n9600 & n19368 ;
  assign n19884 = n9593 | n19883 ;
  assign n19885 = ( n19882 & n19883 ) | ( n19882 & n19884 ) | ( n19883 & n19884 ) ;
  assign n19886 = n9592 | n19885 ;
  assign n19887 = ~n19701 & n19703 ;
  assign n19888 = ~n19372 & n19701 ;
  assign n19889 = n19882 & ~n19888 ;
  assign n19890 = ~n19887 & n19889 ;
  assign n19891 = n19882 | n19887 ;
  assign n19892 = ( n19701 & ~n19702 ) | ( n19701 & n19891 ) | ( ~n19702 & n19891 ) ;
  assign n19893 = ( ~n19882 & n19890 ) | ( ~n19882 & n19892 ) | ( n19890 & n19892 ) ;
  assign n19894 = ( n19885 & n19886 ) | ( n19885 & ~n19893 ) | ( n19886 & ~n19893 ) ;
  assign n19895 = x2 & ~n19894 ;
  assign n19896 = ( ~x2 & n19861 ) | ( ~x2 & n19894 ) | ( n19861 & n19894 ) ;
  assign n19897 = ( ~n19862 & n19895 ) | ( ~n19862 & n19896 ) | ( n19895 & n19896 ) ;
  assign n19898 = ( n19718 & ~n19860 ) | ( n19718 & n19897 ) | ( ~n19860 & n19897 ) ;
  assign n19899 = ( n19718 & n19860 ) | ( n19718 & ~n19897 ) | ( n19860 & ~n19897 ) ;
  assign n19900 = ( ~n19718 & n19898 ) | ( ~n19718 & n19899 ) | ( n19898 & n19899 ) ;
  assign n19901 = n19720 & n19900 ;
  assign n19902 = n19720 | n19900 ;
  assign n19903 = ~n19901 & n19902 ;
  assign n19904 = n3515 | n3529 ;
  assign n19905 = ( n19873 & n19875 ) | ( n19873 & n19904 ) | ( n19875 & n19904 ) ;
  assign n19906 = ( n19683 & ~n19874 ) | ( n19683 & n19904 ) | ( ~n19874 & n19904 ) ;
  assign n19907 = ( n19873 & ~n19905 ) | ( n19873 & n19906 ) | ( ~n19905 & n19906 ) ;
  assign n19908 = n66 & ~n19872 ;
  assign n19909 = n3270 & n19908 ;
  assign n19910 = ( n13671 & n19908 ) | ( n13671 & n19909 ) | ( n19908 & n19909 ) ;
  assign n19911 = ( ~n19864 & n19907 ) | ( ~n19864 & n19910 ) | ( n19907 & n19910 ) ;
  assign n19912 = ( n19864 & n19907 ) | ( n19864 & n19910 ) | ( n19907 & n19910 ) ;
  assign n19913 = ( n19864 & n19911 ) | ( n19864 & ~n19912 ) | ( n19911 & ~n19912 ) ;
  assign n19914 = ( ~n19878 & n19881 ) | ( ~n19878 & n19913 ) | ( n19881 & n19913 ) ;
  assign n19915 = ( n19878 & n19881 ) | ( n19878 & n19913 ) | ( n19881 & n19913 ) ;
  assign n19916 = ( n19878 & n19914 ) | ( n19878 & ~n19915 ) | ( n19914 & ~n19915 ) ;
  assign n19917 = ~n19891 & n19916 ;
  assign n19918 = ( ~n19889 & n19891 ) | ( ~n19889 & n19916 ) | ( n19891 & n19916 ) ;
  assign n19919 = ~n19889 & n19916 ;
  assign n19920 = ( n19917 & n19918 ) | ( n19917 & ~n19919 ) | ( n19918 & ~n19919 ) ;
  assign n19921 = n9592 & n19920 ;
  assign n19922 = n9593 & n19916 ;
  assign n19923 = n41 & n19882 ;
  assign n19924 = n19922 | n19923 ;
  assign n19925 = x2 | n19924 ;
  assign n19926 = ( ~n19921 & n19924 ) | ( ~n19921 & n19925 ) | ( n19924 & n19925 ) ;
  assign n19927 = n9591 & n19920 ;
  assign n19928 = n19926 | n19927 ;
  assign n19929 = n9600 & ~n19701 ;
  assign n19930 = ( x2 & n19924 ) | ( x2 & n19929 ) | ( n19924 & n19929 ) ;
  assign n19931 = n19928 & ~n19930 ;
  assign n19932 = n7346 & ~n19182 ;
  assign n19933 = x8 & n19932 ;
  assign n19934 = n7341 & ~n18362 ;
  assign n19935 = n7345 | n19934 ;
  assign n19936 = ( n19177 & n19934 ) | ( n19177 & n19935 ) | ( n19934 & n19935 ) ;
  assign n19937 = n7644 & n18730 ;
  assign n19938 = n19936 | n19937 ;
  assign n19939 = x8 & ~n19938 ;
  assign n19940 = ( ~x8 & n19932 ) | ( ~x8 & n19938 ) | ( n19932 & n19938 ) ;
  assign n19941 = ( ~n19933 & n19939 ) | ( ~n19933 & n19940 ) | ( n19939 & n19940 ) ;
  assign n19942 = n6796 & ~n17963 ;
  assign n19943 = x11 & n19942 ;
  assign n19944 = n6567 & n17742 ;
  assign n19945 = n6570 | n19944 ;
  assign n19946 = ( ~n18258 & n19944 ) | ( ~n18258 & n19945 ) | ( n19944 & n19945 ) ;
  assign n19947 = n6571 | n19946 ;
  assign n19948 = ( n18268 & n19946 ) | ( n18268 & n19947 ) | ( n19946 & n19947 ) ;
  assign n19949 = x11 & ~n19948 ;
  assign n19950 = ( ~x11 & n19942 ) | ( ~x11 & n19948 ) | ( n19942 & n19948 ) ;
  assign n19951 = ( ~n19943 & n19949 ) | ( ~n19943 & n19950 ) | ( n19949 & n19950 ) ;
  assign n19952 = n6332 & n17346 ;
  assign n19953 = x14 & n19952 ;
  assign n19954 = n5909 & ~n17126 ;
  assign n19955 = n5914 | n19954 ;
  assign n19956 = ( ~n17635 & n19954 ) | ( ~n17635 & n19955 ) | ( n19954 & n19955 ) ;
  assign n19957 = n5915 | n19956 ;
  assign n19958 = ( ~n17646 & n19956 ) | ( ~n17646 & n19957 ) | ( n19956 & n19957 ) ;
  assign n19959 = x14 & ~n19958 ;
  assign n19960 = ( ~x14 & n19952 ) | ( ~x14 & n19958 ) | ( n19952 & n19958 ) ;
  assign n19961 = ( ~n19953 & n19959 ) | ( ~n19953 & n19960 ) | ( n19959 & n19960 ) ;
  assign n19962 = n5584 & n16724 ;
  assign n19963 = x17 & n19962 ;
  assign n19964 = n5413 & ~n16531 ;
  assign n19965 = n5417 | n19964 ;
  assign n19966 = ( n16925 & n19964 ) | ( n16925 & n19965 ) | ( n19964 & n19965 ) ;
  assign n19967 = n5418 | n19966 ;
  assign n19968 = ( ~n16936 & n19966 ) | ( ~n16936 & n19967 ) | ( n19966 & n19967 ) ;
  assign n19969 = x17 & ~n19968 ;
  assign n19970 = ( ~x17 & n19962 ) | ( ~x17 & n19968 ) | ( n19962 & n19968 ) ;
  assign n19971 = ( ~n19963 & n19969 ) | ( ~n19963 & n19970 ) | ( n19969 & n19970 ) ;
  assign n19972 = n5232 & ~n16150 ;
  assign n19973 = x20 & n19972 ;
  assign n19974 = n4874 & ~n15954 ;
  assign n19975 = n4878 | n19974 ;
  assign n19976 = ( ~n16338 & n19974 ) | ( ~n16338 & n19975 ) | ( n19974 & n19975 ) ;
  assign n19977 = n4879 | n19976 ;
  assign n19978 = ( ~n16349 & n19976 ) | ( ~n16349 & n19977 ) | ( n19976 & n19977 ) ;
  assign n19979 = x20 & ~n19978 ;
  assign n19980 = ( ~x20 & n19972 ) | ( ~x20 & n19978 ) | ( n19972 & n19978 ) ;
  assign n19981 = ( ~n19973 & n19979 ) | ( ~n19973 & n19980 ) | ( n19979 & n19980 ) ;
  assign n19982 = n4215 & ~n15184 ;
  assign n19983 = n4200 & n14942 ;
  assign n19984 = n2083 & ~n14723 ;
  assign n19985 = n19983 | n19984 ;
  assign n19986 = n19982 | n19985 ;
  assign n19987 = x26 & n19986 ;
  assign n19988 = n4203 & ~n15195 ;
  assign n19989 = ( ~x26 & n19986 ) | ( ~x26 & n19988 ) | ( n19986 & n19988 ) ;
  assign n19990 = x26 & ~n19988 ;
  assign n19991 = ( ~n19987 & n19989 ) | ( ~n19987 & n19990 ) | ( n19989 & n19990 ) ;
  assign n19992 = n4039 & n14520 ;
  assign n19993 = n3541 | n19992 ;
  assign n19994 = ( n14531 & n19992 ) | ( n14531 & n19993 ) | ( n19992 & n19993 ) ;
  assign n19995 = n3536 & n13992 ;
  assign n19996 = ( ~x29 & n19994 ) | ( ~x29 & n19995 ) | ( n19994 & n19995 ) ;
  assign n19997 = n3501 & n14352 ;
  assign n19998 = x29 & ~n19995 ;
  assign n19999 = n19997 | n19998 ;
  assign n20000 = ( n19994 & n19997 ) | ( n19994 & n19998 ) | ( n19997 & n19998 ) ;
  assign n20001 = ( n19996 & n19999 ) | ( n19996 & ~n20000 ) | ( n19999 & ~n20000 ) ;
  assign n20002 = n83 | n1859 ;
  assign n20003 = ~n2105 & n2283 ;
  assign n20004 = ~n20002 & n20003 ;
  assign n20005 = n5986 | n6065 ;
  assign n20006 = n20004 & ~n20005 ;
  assign n20007 = n854 | n907 ;
  assign n20008 = n3037 | n3465 ;
  assign n20009 = n20007 | n20008 ;
  assign n20010 = n199 | n347 ;
  assign n20011 = n2158 | n20010 ;
  assign n20012 = n2480 | n20011 ;
  assign n20013 = n20009 | n20012 ;
  assign n20014 = n15523 | n20013 ;
  assign n20015 = n20006 & ~n20014 ;
  assign n20016 = n1117 | n2886 ;
  assign n20017 = n20015 & ~n20016 ;
  assign n20018 = n3273 & ~n14000 ;
  assign n20019 = n3270 | n20018 ;
  assign n20020 = ( n13996 & n20018 ) | ( n13996 & n20019 ) | ( n20018 & n20019 ) ;
  assign n20021 = n390 | n20020 ;
  assign n20022 = ( ~n14130 & n20020 ) | ( ~n14130 & n20021 ) | ( n20020 & n20021 ) ;
  assign n20023 = n3274 & n13998 ;
  assign n20024 = n20022 | n20023 ;
  assign n20025 = ( n19812 & ~n20017 ) | ( n19812 & n20024 ) | ( ~n20017 & n20024 ) ;
  assign n20026 = ( n19812 & n20017 ) | ( n19812 & ~n20024 ) | ( n20017 & ~n20024 ) ;
  assign n20027 = ( ~n19812 & n20025 ) | ( ~n19812 & n20026 ) | ( n20025 & n20026 ) ;
  assign n20028 = ( n19815 & n20001 ) | ( n19815 & ~n20027 ) | ( n20001 & ~n20027 ) ;
  assign n20029 = ( n19815 & ~n20001 ) | ( n19815 & n20027 ) | ( ~n20001 & n20027 ) ;
  assign n20030 = ( ~n19815 & n20028 ) | ( ~n19815 & n20029 ) | ( n20028 & n20029 ) ;
  assign n20031 = ( n19817 & n19991 ) | ( n19817 & ~n20030 ) | ( n19991 & ~n20030 ) ;
  assign n20032 = ( n19817 & ~n19991 ) | ( n19817 & n20030 ) | ( ~n19991 & n20030 ) ;
  assign n20033 = ( ~n19817 & n20031 ) | ( ~n19817 & n20032 ) | ( n20031 & n20032 ) ;
  assign n20034 = n4637 & n15561 ;
  assign n20035 = x23 & n20034 ;
  assign n20036 = n4584 & ~n15394 ;
  assign n20037 = n4649 | n20036 ;
  assign n20038 = ( ~n15806 & n20036 ) | ( ~n15806 & n20037 ) | ( n20036 & n20037 ) ;
  assign n20039 = n4591 | n20038 ;
  assign n20040 = ( n15817 & n20038 ) | ( n15817 & n20039 ) | ( n20038 & n20039 ) ;
  assign n20041 = x23 & ~n20040 ;
  assign n20042 = ( ~x23 & n20034 ) | ( ~x23 & n20040 ) | ( n20034 & n20040 ) ;
  assign n20043 = ( ~n20035 & n20041 ) | ( ~n20035 & n20042 ) | ( n20041 & n20042 ) ;
  assign n20044 = ( n19830 & n20033 ) | ( n19830 & ~n20043 ) | ( n20033 & ~n20043 ) ;
  assign n20045 = ( n19830 & ~n20033 ) | ( n19830 & n20043 ) | ( ~n20033 & n20043 ) ;
  assign n20046 = ( ~n19830 & n20044 ) | ( ~n19830 & n20045 ) | ( n20044 & n20045 ) ;
  assign n20047 = ( n19833 & ~n19981 ) | ( n19833 & n20046 ) | ( ~n19981 & n20046 ) ;
  assign n20048 = ( n19833 & n19981 ) | ( n19833 & ~n20046 ) | ( n19981 & ~n20046 ) ;
  assign n20049 = ( ~n19833 & n20047 ) | ( ~n19833 & n20048 ) | ( n20047 & n20048 ) ;
  assign n20050 = ( n19836 & n19971 ) | ( n19836 & ~n20049 ) | ( n19971 & ~n20049 ) ;
  assign n20051 = ( n19836 & ~n19971 ) | ( n19836 & n20049 ) | ( ~n19971 & n20049 ) ;
  assign n20052 = ( ~n19836 & n20050 ) | ( ~n19836 & n20051 ) | ( n20050 & n20051 ) ;
  assign n20053 = ( n19840 & n19961 ) | ( n19840 & ~n20052 ) | ( n19961 & ~n20052 ) ;
  assign n20054 = ( n19840 & ~n19961 ) | ( n19840 & n20052 ) | ( ~n19961 & n20052 ) ;
  assign n20055 = ( ~n19840 & n20053 ) | ( ~n19840 & n20054 ) | ( n20053 & n20054 ) ;
  assign n20056 = ( n19842 & n19951 ) | ( n19842 & ~n20055 ) | ( n19951 & ~n20055 ) ;
  assign n20057 = ( n19842 & ~n19951 ) | ( n19842 & n20055 ) | ( ~n19951 & n20055 ) ;
  assign n20058 = ( ~n19842 & n20056 ) | ( ~n19842 & n20057 ) | ( n20056 & n20057 ) ;
  assign n20059 = ( n19846 & n19941 ) | ( n19846 & ~n20058 ) | ( n19941 & ~n20058 ) ;
  assign n20060 = ( n19846 & ~n19941 ) | ( n19846 & n20058 ) | ( ~n19941 & n20058 ) ;
  assign n20061 = ( ~n19846 & n20059 ) | ( ~n19846 & n20060 ) | ( n20059 & n20060 ) ;
  assign n20062 = n40 & n19368 ;
  assign n20063 = n8721 & ~n19315 ;
  assign n20064 = n8340 & n19248 ;
  assign n20065 = n20063 | n20064 ;
  assign n20066 = n20062 | n20065 ;
  assign n20067 = x5 & n20066 ;
  assign n20068 = n8341 & ~n19374 ;
  assign n20069 = ( ~x5 & n20066 ) | ( ~x5 & n20068 ) | ( n20066 & n20068 ) ;
  assign n20070 = x5 & ~n20068 ;
  assign n20071 = ( ~n20067 & n20069 ) | ( ~n20067 & n20070 ) | ( n20069 & n20070 ) ;
  assign n20072 = ( n19859 & n20061 ) | ( n19859 & n20071 ) | ( n20061 & n20071 ) ;
  assign n20073 = ( n19859 & ~n20061 ) | ( n19859 & n20071 ) | ( ~n20061 & n20071 ) ;
  assign n20074 = ( n20061 & ~n20072 ) | ( n20061 & n20073 ) | ( ~n20072 & n20073 ) ;
  assign n20075 = ( n19898 & n19931 ) | ( n19898 & ~n20074 ) | ( n19931 & ~n20074 ) ;
  assign n20076 = ( n19898 & ~n19931 ) | ( n19898 & n20074 ) | ( ~n19931 & n20074 ) ;
  assign n20077 = ( ~n19898 & n20075 ) | ( ~n19898 & n20076 ) | ( n20075 & n20076 ) ;
  assign n20078 = n19902 | n20077 ;
  assign n20079 = n19902 & n20077 ;
  assign n20080 = n20078 & ~n20079 ;
  assign n20081 = x31 | n66 ;
  assign n20082 = ( n3272 & n3529 ) | ( n3272 & n20081 ) | ( n3529 & n20081 ) ;
  assign n20083 = n19864 | n20082 ;
  assign n20084 = n19864 & n20082 ;
  assign n20085 = n20083 & ~n20084 ;
  assign n20086 = ( n19906 & ~n19912 ) | ( n19906 & n20085 ) | ( ~n19912 & n20085 ) ;
  assign n20087 = ( n19906 & n19912 ) | ( n19906 & n20085 ) | ( n19912 & n20085 ) ;
  assign n20088 = ( n19912 & n20086 ) | ( n19912 & ~n20087 ) | ( n20086 & ~n20087 ) ;
  assign n20089 = n19915 | n20088 ;
  assign n20090 = n19915 & n20088 ;
  assign n20091 = n20089 & ~n20090 ;
  assign n20092 = n9593 & n20091 ;
  assign n20093 = n9592 | n20092 ;
  assign n20094 = n19889 | n19916 ;
  assign n20095 = n20091 | n20094 ;
  assign n20096 = n20091 & n20094 ;
  assign n20097 = n20095 & ~n20096 ;
  assign n20098 = n19891 & n19916 ;
  assign n20099 = ( n20091 & ~n20094 ) | ( n20091 & n20098 ) | ( ~n20094 & n20098 ) ;
  assign n20100 = ( n20094 & n20096 ) | ( n20094 & ~n20098 ) | ( n20096 & ~n20098 ) ;
  assign n20101 = ( n20097 & n20099 ) | ( n20097 & n20100 ) | ( n20099 & n20100 ) ;
  assign n20102 = ( n20092 & n20093 ) | ( n20092 & n20101 ) | ( n20093 & n20101 ) ;
  assign n20103 = n41 & n19916 ;
  assign n20104 = ( x2 & ~n20102 ) | ( x2 & n20103 ) | ( ~n20102 & n20103 ) ;
  assign n20105 = ~x2 & n20102 ;
  assign n20106 = n9600 & n19882 ;
  assign n20107 = ( x2 & n20103 ) | ( x2 & n20106 ) | ( n20103 & n20106 ) ;
  assign n20108 = ( n20104 & n20105 ) | ( n20104 & ~n20107 ) | ( n20105 & ~n20107 ) ;
  assign n20109 = n40 & ~n19701 ;
  assign n20110 = n8721 & n19368 ;
  assign n20111 = n8340 & ~n19315 ;
  assign n20112 = n20110 | n20111 ;
  assign n20113 = n20109 | n20112 ;
  assign n20114 = x5 & n20113 ;
  assign n20115 = n8341 & ~n19706 ;
  assign n20116 = ( ~x5 & n20113 ) | ( ~x5 & n20115 ) | ( n20113 & n20115 ) ;
  assign n20117 = x5 & ~n20115 ;
  assign n20118 = ( ~n20114 & n20116 ) | ( ~n20114 & n20117 ) | ( n20116 & n20117 ) ;
  assign n20119 = n7644 & n19177 ;
  assign n20120 = x8 & n20119 ;
  assign n20121 = n7341 & n18730 ;
  assign n20122 = n7345 | n20121 ;
  assign n20123 = ( n19248 & n20121 ) | ( n19248 & n20122 ) | ( n20121 & n20122 ) ;
  assign n20124 = n7346 | n20123 ;
  assign n20125 = ( n19253 & n20123 ) | ( n19253 & n20124 ) | ( n20123 & n20124 ) ;
  assign n20126 = x8 & ~n20125 ;
  assign n20127 = ( ~x8 & n20119 ) | ( ~x8 & n20125 ) | ( n20119 & n20125 ) ;
  assign n20128 = ( ~n20120 & n20126 ) | ( ~n20120 & n20127 ) | ( n20126 & n20127 ) ;
  assign n20129 = n3501 & n14520 ;
  assign n20130 = x29 & n20129 ;
  assign n20131 = n3536 & n14352 ;
  assign n20132 = n4039 | n20131 ;
  assign n20133 = ( ~n14723 & n20131 ) | ( ~n14723 & n20132 ) | ( n20131 & n20132 ) ;
  assign n20134 = n3541 | n20133 ;
  assign n20135 = ( ~n14734 & n20133 ) | ( ~n14734 & n20134 ) | ( n20133 & n20134 ) ;
  assign n20136 = x29 & ~n20135 ;
  assign n20137 = ( ~x29 & n20129 ) | ( ~x29 & n20135 ) | ( n20129 & n20135 ) ;
  assign n20138 = ( ~n20130 & n20136 ) | ( ~n20130 & n20137 ) | ( n20136 & n20137 ) ;
  assign n20139 = n3274 & n13996 ;
  assign n20140 = n3273 & n13998 ;
  assign n20141 = n20139 | n20140 ;
  assign n20142 = n390 | n20141 ;
  assign n20143 = ( n14024 & n20141 ) | ( n14024 & n20142 ) | ( n20141 & n20142 ) ;
  assign n20144 = n3270 & n13992 ;
  assign n20145 = n20143 | n20144 ;
  assign n20146 = n2152 | n3927 ;
  assign n20147 = n2841 | n15901 ;
  assign n20148 = n864 | n2706 ;
  assign n20149 = n20147 | n20148 ;
  assign n20150 = n404 | n772 ;
  assign n20151 = n265 | n851 ;
  assign n20152 = n20150 | n20151 ;
  assign n20153 = n20149 | n20152 ;
  assign n20154 = n1338 | n6045 ;
  assign n20155 = n20153 | n20154 ;
  assign n20156 = n2276 | n5086 ;
  assign n20157 = n14844 | n20156 ;
  assign n20158 = n2347 | n20157 ;
  assign n20159 = n20155 | n20158 ;
  assign n20160 = n3949 | n20159 ;
  assign n20161 = n20146 | n20160 ;
  assign n20162 = ( ~n20025 & n20145 ) | ( ~n20025 & n20161 ) | ( n20145 & n20161 ) ;
  assign n20163 = ( n20025 & n20145 ) | ( n20025 & n20161 ) | ( n20145 & n20161 ) ;
  assign n20164 = ( n20025 & n20162 ) | ( n20025 & ~n20163 ) | ( n20162 & ~n20163 ) ;
  assign n20165 = ( ~n20028 & n20138 ) | ( ~n20028 & n20164 ) | ( n20138 & n20164 ) ;
  assign n20166 = ( n20028 & n20138 ) | ( n20028 & n20164 ) | ( n20138 & n20164 ) ;
  assign n20167 = ( n20028 & n20165 ) | ( n20028 & ~n20166 ) | ( n20165 & ~n20166 ) ;
  assign n20168 = n4215 & ~n15394 ;
  assign n20169 = n4200 & ~n15184 ;
  assign n20170 = n2083 & n14942 ;
  assign n20171 = n20169 | n20170 ;
  assign n20172 = n20168 | n20171 ;
  assign n20173 = x26 & n20172 ;
  assign n20174 = n4203 & n15405 ;
  assign n20175 = ( ~x26 & n20172 ) | ( ~x26 & n20174 ) | ( n20172 & n20174 ) ;
  assign n20176 = x26 & ~n20174 ;
  assign n20177 = ( ~n20173 & n20175 ) | ( ~n20173 & n20176 ) | ( n20175 & n20176 ) ;
  assign n20178 = ( ~n20031 & n20167 ) | ( ~n20031 & n20177 ) | ( n20167 & n20177 ) ;
  assign n20179 = ( n20031 & n20167 ) | ( n20031 & n20177 ) | ( n20167 & n20177 ) ;
  assign n20180 = ( n20031 & n20178 ) | ( n20031 & ~n20179 ) | ( n20178 & ~n20179 ) ;
  assign n20181 = n4637 & ~n15806 ;
  assign n20182 = x23 & n20181 ;
  assign n20183 = n4584 & n15561 ;
  assign n20184 = n4649 | n20183 ;
  assign n20185 = ( ~n15954 & n20183 ) | ( ~n15954 & n20184 ) | ( n20183 & n20184 ) ;
  assign n20186 = n4591 | n20185 ;
  assign n20187 = ( ~n15965 & n20185 ) | ( ~n15965 & n20186 ) | ( n20185 & n20186 ) ;
  assign n20188 = x23 & ~n20187 ;
  assign n20189 = ( ~x23 & n20181 ) | ( ~x23 & n20187 ) | ( n20181 & n20187 ) ;
  assign n20190 = ( ~n20182 & n20188 ) | ( ~n20182 & n20189 ) | ( n20188 & n20189 ) ;
  assign n20191 = ( n20045 & n20180 ) | ( n20045 & n20190 ) | ( n20180 & n20190 ) ;
  assign n20192 = ( ~n20045 & n20180 ) | ( ~n20045 & n20190 ) | ( n20180 & n20190 ) ;
  assign n20193 = ( n20045 & ~n20191 ) | ( n20045 & n20192 ) | ( ~n20191 & n20192 ) ;
  assign n20194 = n4879 & ~n16542 ;
  assign n20195 = x20 & n20194 ;
  assign n20196 = n4874 & ~n16150 ;
  assign n20197 = n4878 | n20196 ;
  assign n20198 = ( ~n16531 & n20196 ) | ( ~n16531 & n20197 ) | ( n20196 & n20197 ) ;
  assign n20199 = n5232 & ~n16338 ;
  assign n20200 = n20198 | n20199 ;
  assign n20201 = x20 & ~n20200 ;
  assign n20202 = ( ~x20 & n20194 ) | ( ~x20 & n20200 ) | ( n20194 & n20200 ) ;
  assign n20203 = ( ~n20195 & n20201 ) | ( ~n20195 & n20202 ) | ( n20201 & n20202 ) ;
  assign n20204 = ( ~n20048 & n20193 ) | ( ~n20048 & n20203 ) | ( n20193 & n20203 ) ;
  assign n20205 = ( n20048 & n20193 ) | ( n20048 & n20203 ) | ( n20193 & n20203 ) ;
  assign n20206 = ( n20048 & n20204 ) | ( n20048 & ~n20205 ) | ( n20204 & ~n20205 ) ;
  assign n20207 = n5584 & n16925 ;
  assign n20208 = x17 & n20207 ;
  assign n20209 = n5413 & n16724 ;
  assign n20210 = n5417 | n20209 ;
  assign n20211 = ( ~n17126 & n20209 ) | ( ~n17126 & n20210 ) | ( n20209 & n20210 ) ;
  assign n20212 = n5418 | n20211 ;
  assign n20213 = ( ~n17139 & n20211 ) | ( ~n17139 & n20212 ) | ( n20211 & n20212 ) ;
  assign n20214 = x17 & ~n20213 ;
  assign n20215 = ( ~x17 & n20207 ) | ( ~x17 & n20213 ) | ( n20207 & n20213 ) ;
  assign n20216 = ( ~n20208 & n20214 ) | ( ~n20208 & n20215 ) | ( n20214 & n20215 ) ;
  assign n20217 = ( n20050 & n20206 ) | ( n20050 & n20216 ) | ( n20206 & n20216 ) ;
  assign n20218 = ( ~n20050 & n20206 ) | ( ~n20050 & n20216 ) | ( n20206 & n20216 ) ;
  assign n20219 = ( n20050 & ~n20217 ) | ( n20050 & n20218 ) | ( ~n20217 & n20218 ) ;
  assign n20220 = n5914 & n17742 ;
  assign n20221 = x14 & n20220 ;
  assign n20222 = n6332 & ~n17635 ;
  assign n20223 = n5909 & n17346 ;
  assign n20224 = n20222 | n20223 ;
  assign n20225 = n5915 | n20224 ;
  assign n20226 = ( ~n17749 & n20224 ) | ( ~n17749 & n20225 ) | ( n20224 & n20225 ) ;
  assign n20227 = x14 & ~n20226 ;
  assign n20228 = ( ~x14 & n20220 ) | ( ~x14 & n20226 ) | ( n20220 & n20226 ) ;
  assign n20229 = ( ~n20221 & n20227 ) | ( ~n20221 & n20228 ) | ( n20227 & n20228 ) ;
  assign n20230 = ( ~n20053 & n20219 ) | ( ~n20053 & n20229 ) | ( n20219 & n20229 ) ;
  assign n20231 = ( n20053 & n20219 ) | ( n20053 & n20229 ) | ( n20219 & n20229 ) ;
  assign n20232 = ( n20053 & n20230 ) | ( n20053 & ~n20231 ) | ( n20230 & ~n20231 ) ;
  assign n20233 = n6796 & ~n18258 ;
  assign n20234 = x11 & n20233 ;
  assign n20235 = n6567 & ~n17963 ;
  assign n20236 = n6570 | n20235 ;
  assign n20237 = ( ~n18362 & n20235 ) | ( ~n18362 & n20236 ) | ( n20235 & n20236 ) ;
  assign n20238 = n6571 | n20237 ;
  assign n20239 = ( ~n18373 & n20237 ) | ( ~n18373 & n20238 ) | ( n20237 & n20238 ) ;
  assign n20240 = x11 & ~n20239 ;
  assign n20241 = ( ~x11 & n20233 ) | ( ~x11 & n20239 ) | ( n20233 & n20239 ) ;
  assign n20242 = ( ~n20234 & n20240 ) | ( ~n20234 & n20241 ) | ( n20240 & n20241 ) ;
  assign n20243 = ( n20056 & n20232 ) | ( n20056 & n20242 ) | ( n20232 & n20242 ) ;
  assign n20244 = ( ~n20056 & n20232 ) | ( ~n20056 & n20242 ) | ( n20232 & n20242 ) ;
  assign n20245 = ( n20056 & ~n20243 ) | ( n20056 & n20244 ) | ( ~n20243 & n20244 ) ;
  assign n20246 = ( ~n20059 & n20128 ) | ( ~n20059 & n20245 ) | ( n20128 & n20245 ) ;
  assign n20247 = ( n20059 & n20128 ) | ( n20059 & n20245 ) | ( n20128 & n20245 ) ;
  assign n20248 = ( n20059 & n20246 ) | ( n20059 & ~n20247 ) | ( n20246 & ~n20247 ) ;
  assign n20249 = ( n20073 & n20118 ) | ( n20073 & n20248 ) | ( n20118 & n20248 ) ;
  assign n20250 = ( ~n20073 & n20118 ) | ( ~n20073 & n20248 ) | ( n20118 & n20248 ) ;
  assign n20251 = ( n20073 & ~n20249 ) | ( n20073 & n20250 ) | ( ~n20249 & n20250 ) ;
  assign n20252 = ( ~n20075 & n20108 ) | ( ~n20075 & n20251 ) | ( n20108 & n20251 ) ;
  assign n20253 = ( n20075 & n20108 ) | ( n20075 & n20251 ) | ( n20108 & n20251 ) ;
  assign n20254 = ( n20075 & n20252 ) | ( n20075 & ~n20253 ) | ( n20252 & ~n20253 ) ;
  assign n20255 = n20078 | n20254 ;
  assign n20256 = n20078 & n20254 ;
  assign n20257 = n20255 & ~n20256 ;
  assign n20258 = ~n20078 & n20254 ;
  assign n20259 = n6570 & n18730 ;
  assign n20260 = n6571 | n20259 ;
  assign n20261 = ( n18735 & n20259 ) | ( n18735 & n20260 ) | ( n20259 & n20260 ) ;
  assign n20262 = n6567 & ~n18258 ;
  assign n20263 = ( ~x11 & n20261 ) | ( ~x11 & n20262 ) | ( n20261 & n20262 ) ;
  assign n20264 = n6796 & ~n18362 ;
  assign n20265 = x11 & ~n20262 ;
  assign n20266 = n20264 | n20265 ;
  assign n20267 = ( n20261 & n20264 ) | ( n20261 & n20265 ) | ( n20264 & n20265 ) ;
  assign n20268 = ( n20263 & n20266 ) | ( n20263 & ~n20267 ) | ( n20266 & ~n20267 ) ;
  assign n20269 = n5915 & ~n17976 ;
  assign n20270 = x14 & n20269 ;
  assign n20271 = n5909 & ~n17635 ;
  assign n20272 = n5914 | n20271 ;
  assign n20273 = ( ~n17963 & n20271 ) | ( ~n17963 & n20272 ) | ( n20271 & n20272 ) ;
  assign n20274 = n6332 & n17742 ;
  assign n20275 = n20273 | n20274 ;
  assign n20276 = x14 & ~n20275 ;
  assign n20277 = ( ~x14 & n20269 ) | ( ~x14 & n20275 ) | ( n20269 & n20275 ) ;
  assign n20278 = ( ~n20270 & n20276 ) | ( ~n20270 & n20277 ) | ( n20276 & n20277 ) ;
  assign n20279 = n4878 & n16724 ;
  assign n20280 = n5232 & ~n16531 ;
  assign n20281 = n4874 & ~n16338 ;
  assign n20282 = n20280 | n20281 ;
  assign n20283 = n20279 | n20282 ;
  assign n20284 = x20 & n20283 ;
  assign n20285 = n4879 & n16735 ;
  assign n20286 = ( ~x20 & n20283 ) | ( ~x20 & n20285 ) | ( n20283 & n20285 ) ;
  assign n20287 = x20 & ~n20285 ;
  assign n20288 = ( ~n20284 & n20286 ) | ( ~n20284 & n20287 ) | ( n20286 & n20287 ) ;
  assign n20289 = n4215 & n15561 ;
  assign n20290 = n4200 & ~n15394 ;
  assign n20291 = n2083 & ~n15184 ;
  assign n20292 = n20290 | n20291 ;
  assign n20293 = n20289 | n20292 ;
  assign n20294 = x26 & n20293 ;
  assign n20295 = n4203 & n15573 ;
  assign n20296 = ( ~x26 & n20293 ) | ( ~x26 & n20295 ) | ( n20293 & n20295 ) ;
  assign n20297 = x26 & ~n20295 ;
  assign n20298 = ( ~n20294 & n20296 ) | ( ~n20294 & n20297 ) | ( n20296 & n20297 ) ;
  assign n20299 = n390 & n14363 ;
  assign n20300 = n3270 & n14352 ;
  assign n20301 = n3274 & n13992 ;
  assign n20302 = n3273 & n13996 ;
  assign n20303 = n20301 | n20302 ;
  assign n20304 = n20300 | n20303 ;
  assign n20305 = n20299 | n20304 ;
  assign n20306 = n2714 | n3769 ;
  assign n20307 = n788 | n2841 ;
  assign n20308 = n5936 | n20307 ;
  assign n20309 = n2267 | n20308 ;
  assign n20310 = n1019 | n2131 ;
  assign n20311 = n1106 | n20310 ;
  assign n20312 = n2247 | n20311 ;
  assign n20313 = n20309 | n20312 ;
  assign n20314 = n227 | n1294 ;
  assign n20315 = n4807 | n20314 ;
  assign n20316 = n14460 | n20315 ;
  assign n20317 = n20313 | n20316 ;
  assign n20318 = n20306 | n20317 ;
  assign n20319 = n6048 & ~n20318 ;
  assign n20320 = ( n20163 & n20305 ) | ( n20163 & ~n20319 ) | ( n20305 & ~n20319 ) ;
  assign n20321 = ( n20163 & ~n20305 ) | ( n20163 & n20319 ) | ( ~n20305 & n20319 ) ;
  assign n20322 = ( ~n20163 & n20320 ) | ( ~n20163 & n20321 ) | ( n20320 & n20321 ) ;
  assign n20323 = n3501 & ~n14723 ;
  assign n20324 = x29 & n20323 ;
  assign n20325 = n3536 & n14520 ;
  assign n20326 = n4039 | n20325 ;
  assign n20327 = ( n14942 & n20325 ) | ( n14942 & n20326 ) | ( n20325 & n20326 ) ;
  assign n20328 = n3541 | n20327 ;
  assign n20329 = ( ~n14953 & n20327 ) | ( ~n14953 & n20328 ) | ( n20327 & n20328 ) ;
  assign n20330 = x29 & ~n20329 ;
  assign n20331 = ( ~x29 & n20323 ) | ( ~x29 & n20329 ) | ( n20323 & n20329 ) ;
  assign n20332 = ( ~n20324 & n20330 ) | ( ~n20324 & n20331 ) | ( n20330 & n20331 ) ;
  assign n20333 = ( n20166 & ~n20322 ) | ( n20166 & n20332 ) | ( ~n20322 & n20332 ) ;
  assign n20334 = ( n20166 & n20322 ) | ( n20166 & ~n20332 ) | ( n20322 & ~n20332 ) ;
  assign n20335 = ( ~n20166 & n20333 ) | ( ~n20166 & n20334 ) | ( n20333 & n20334 ) ;
  assign n20336 = ( n20179 & ~n20298 ) | ( n20179 & n20335 ) | ( ~n20298 & n20335 ) ;
  assign n20337 = ( n20179 & n20298 ) | ( n20179 & ~n20335 ) | ( n20298 & ~n20335 ) ;
  assign n20338 = ( ~n20179 & n20336 ) | ( ~n20179 & n20337 ) | ( n20336 & n20337 ) ;
  assign n20339 = n4591 & ~n16161 ;
  assign n20340 = x23 & n20339 ;
  assign n20341 = n4649 & ~n16150 ;
  assign n20342 = n4637 & ~n15954 ;
  assign n20343 = n4584 & ~n15806 ;
  assign n20344 = n20342 | n20343 ;
  assign n20345 = n20341 | n20344 ;
  assign n20346 = x23 & ~n20345 ;
  assign n20347 = ( ~x23 & n20339 ) | ( ~x23 & n20345 ) | ( n20339 & n20345 ) ;
  assign n20348 = ( ~n20340 & n20346 ) | ( ~n20340 & n20347 ) | ( n20346 & n20347 ) ;
  assign n20349 = ( n20191 & ~n20338 ) | ( n20191 & n20348 ) | ( ~n20338 & n20348 ) ;
  assign n20350 = ( n20191 & n20338 ) | ( n20191 & ~n20348 ) | ( n20338 & ~n20348 ) ;
  assign n20351 = ( ~n20191 & n20349 ) | ( ~n20191 & n20350 ) | ( n20349 & n20350 ) ;
  assign n20352 = ( n20205 & n20288 ) | ( n20205 & ~n20351 ) | ( n20288 & ~n20351 ) ;
  assign n20353 = ( n20205 & ~n20288 ) | ( n20205 & n20351 ) | ( ~n20288 & n20351 ) ;
  assign n20354 = ( ~n20205 & n20352 ) | ( ~n20205 & n20353 ) | ( n20352 & n20353 ) ;
  assign n20355 = n5584 & ~n17126 ;
  assign n20356 = x17 & n20355 ;
  assign n20357 = n5413 & n16925 ;
  assign n20358 = n5417 | n20357 ;
  assign n20359 = ( n17346 & n20357 ) | ( n17346 & n20358 ) | ( n20357 & n20358 ) ;
  assign n20360 = n5418 | n20359 ;
  assign n20361 = ( ~n17356 & n20359 ) | ( ~n17356 & n20360 ) | ( n20359 & n20360 ) ;
  assign n20362 = x17 & ~n20361 ;
  assign n20363 = ( ~x17 & n20355 ) | ( ~x17 & n20361 ) | ( n20355 & n20361 ) ;
  assign n20364 = ( ~n20356 & n20362 ) | ( ~n20356 & n20363 ) | ( n20362 & n20363 ) ;
  assign n20365 = ( n20217 & ~n20354 ) | ( n20217 & n20364 ) | ( ~n20354 & n20364 ) ;
  assign n20366 = ( n20217 & n20354 ) | ( n20217 & ~n20364 ) | ( n20354 & ~n20364 ) ;
  assign n20367 = ( ~n20217 & n20365 ) | ( ~n20217 & n20366 ) | ( n20365 & n20366 ) ;
  assign n20368 = ( n20231 & n20278 ) | ( n20231 & ~n20367 ) | ( n20278 & ~n20367 ) ;
  assign n20369 = ( n20231 & ~n20278 ) | ( n20231 & n20367 ) | ( ~n20278 & n20367 ) ;
  assign n20370 = ( ~n20231 & n20368 ) | ( ~n20231 & n20369 ) | ( n20368 & n20369 ) ;
  assign n20371 = ( n20243 & ~n20268 ) | ( n20243 & n20370 ) | ( ~n20268 & n20370 ) ;
  assign n20372 = ( n20243 & n20268 ) | ( n20243 & ~n20370 ) | ( n20268 & ~n20370 ) ;
  assign n20373 = ( ~n20243 & n20371 ) | ( ~n20243 & n20372 ) | ( n20371 & n20372 ) ;
  assign n20374 = n7644 & n19248 ;
  assign n20375 = n7346 | n20374 ;
  assign n20376 = ( ~n19320 & n20374 ) | ( ~n19320 & n20375 ) | ( n20374 & n20375 ) ;
  assign n20377 = n7341 & n19177 ;
  assign n20378 = ( ~x8 & n20376 ) | ( ~x8 & n20377 ) | ( n20376 & n20377 ) ;
  assign n20379 = n7345 & ~n19315 ;
  assign n20380 = x8 & ~n20377 ;
  assign n20381 = n20379 | n20380 ;
  assign n20382 = ( n20376 & n20379 ) | ( n20376 & n20380 ) | ( n20379 & n20380 ) ;
  assign n20383 = ( n20378 & n20381 ) | ( n20378 & ~n20382 ) | ( n20381 & ~n20382 ) ;
  assign n20384 = ( n20247 & ~n20373 ) | ( n20247 & n20383 ) | ( ~n20373 & n20383 ) ;
  assign n20385 = ( n20247 & n20373 ) | ( n20247 & ~n20383 ) | ( n20373 & ~n20383 ) ;
  assign n20386 = ( ~n20247 & n20384 ) | ( ~n20247 & n20385 ) | ( n20384 & n20385 ) ;
  assign n20387 = n40 & n19882 ;
  assign n20388 = n8721 & ~n19701 ;
  assign n20389 = n8340 & n19368 ;
  assign n20390 = n20388 | n20389 ;
  assign n20391 = n20387 | n20390 ;
  assign n20392 = x5 & n20391 ;
  assign n20393 = n8341 & ~n19893 ;
  assign n20394 = ( ~x5 & n20391 ) | ( ~x5 & n20393 ) | ( n20391 & n20393 ) ;
  assign n20395 = x5 & ~n20393 ;
  assign n20396 = ( ~n20392 & n20394 ) | ( ~n20392 & n20395 ) | ( n20394 & n20395 ) ;
  assign n20397 = ( n20249 & n20386 ) | ( n20249 & ~n20396 ) | ( n20386 & ~n20396 ) ;
  assign n20398 = ( n20249 & ~n20386 ) | ( n20249 & n20396 ) | ( ~n20386 & n20396 ) ;
  assign n20399 = ( ~n20249 & n20397 ) | ( ~n20249 & n20398 ) | ( n20397 & n20398 ) ;
  assign n20400 = n9593 & ~n20095 ;
  assign n20401 = n41 & n20091 ;
  assign n20402 = n20400 | n20401 ;
  assign n20403 = n9158 & ~n20100 ;
  assign n20404 = n20402 | n20403 ;
  assign n20405 = ~x2 & n20404 ;
  assign n20406 = ( x2 & n9155 ) | ( x2 & ~n19916 ) | ( n9155 & ~n19916 ) ;
  assign n20407 = ~n9592 & n20406 ;
  assign n20408 = ( n20100 & n20406 ) | ( n20100 & n20407 ) | ( n20406 & n20407 ) ;
  assign n20409 = ~n20402 & n20408 ;
  assign n20410 = n20405 | n20409 ;
  assign n20411 = ( n20253 & ~n20399 ) | ( n20253 & n20410 ) | ( ~n20399 & n20410 ) ;
  assign n20412 = ( n20253 & n20399 ) | ( n20253 & ~n20410 ) | ( n20399 & ~n20410 ) ;
  assign n20413 = ( ~n20253 & n20411 ) | ( ~n20253 & n20412 ) | ( n20411 & n20412 ) ;
  assign n20414 = n20258 & ~n20413 ;
  assign n20415 = ~n20258 & n20413 ;
  assign n20416 = n20414 | n20415 ;
  assign n20417 = n7644 & ~n19315 ;
  assign n20418 = x8 & n20417 ;
  assign n20419 = n7341 & n19248 ;
  assign n20420 = n7345 | n20419 ;
  assign n20421 = ( n19368 & n20419 ) | ( n19368 & n20420 ) | ( n20419 & n20420 ) ;
  assign n20422 = n7346 | n20421 ;
  assign n20423 = ( ~n19374 & n20421 ) | ( ~n19374 & n20422 ) | ( n20421 & n20422 ) ;
  assign n20424 = x8 & ~n20423 ;
  assign n20425 = ( ~x8 & n20417 ) | ( ~x8 & n20423 ) | ( n20417 & n20423 ) ;
  assign n20426 = ( ~n20418 & n20424 ) | ( ~n20418 & n20425 ) | ( n20424 & n20425 ) ;
  assign n20427 = n6570 & n19177 ;
  assign n20428 = n6796 & n18730 ;
  assign n20429 = n6567 & ~n18362 ;
  assign n20430 = n20428 | n20429 ;
  assign n20431 = n20427 | n20430 ;
  assign n20432 = x11 & n20431 ;
  assign n20433 = n6571 & ~n19182 ;
  assign n20434 = ( ~x11 & n20431 ) | ( ~x11 & n20433 ) | ( n20431 & n20433 ) ;
  assign n20435 = x11 & ~n20433 ;
  assign n20436 = ( ~n20432 & n20434 ) | ( ~n20432 & n20435 ) | ( n20434 & n20435 ) ;
  assign n20437 = n5232 & n16724 ;
  assign n20438 = x20 & n20437 ;
  assign n20439 = n4874 & ~n16531 ;
  assign n20440 = n4878 | n20439 ;
  assign n20441 = ( n16925 & n20439 ) | ( n16925 & n20440 ) | ( n20439 & n20440 ) ;
  assign n20442 = n4879 | n20441 ;
  assign n20443 = ( ~n16936 & n20441 ) | ( ~n16936 & n20442 ) | ( n20441 & n20442 ) ;
  assign n20444 = x20 & ~n20443 ;
  assign n20445 = ( ~x20 & n20437 ) | ( ~x20 & n20443 ) | ( n20437 & n20443 ) ;
  assign n20446 = ( ~n20438 & n20444 ) | ( ~n20438 & n20445 ) | ( n20444 & n20445 ) ;
  assign n20447 = n4215 & ~n15806 ;
  assign n20448 = n4200 & n15561 ;
  assign n20449 = n2083 & ~n15394 ;
  assign n20450 = n20448 | n20449 ;
  assign n20451 = n20447 | n20450 ;
  assign n20452 = x26 & n20451 ;
  assign n20453 = n4203 & n15817 ;
  assign n20454 = ( ~x26 & n20451 ) | ( ~x26 & n20453 ) | ( n20451 & n20453 ) ;
  assign n20455 = x26 & ~n20453 ;
  assign n20456 = ( ~n20452 & n20454 ) | ( ~n20452 & n20455 ) | ( n20454 & n20455 ) ;
  assign n20457 = n3541 & ~n15195 ;
  assign n20458 = x29 & n20457 ;
  assign n20459 = n3536 & ~n14723 ;
  assign n20460 = n4039 | n20459 ;
  assign n20461 = ( ~n15184 & n20459 ) | ( ~n15184 & n20460 ) | ( n20459 & n20460 ) ;
  assign n20462 = n3501 & n14942 ;
  assign n20463 = n20461 | n20462 ;
  assign n20464 = x29 & ~n20463 ;
  assign n20465 = ( ~x29 & n20457 ) | ( ~x29 & n20463 ) | ( n20457 & n20463 ) ;
  assign n20466 = ( ~n20458 & n20464 ) | ( ~n20458 & n20465 ) | ( n20464 & n20465 ) ;
  assign n20467 = n3273 & n13992 ;
  assign n20468 = n3270 | n20467 ;
  assign n20469 = ( n14520 & n20467 ) | ( n14520 & n20468 ) | ( n20467 & n20468 ) ;
  assign n20470 = n390 | n20469 ;
  assign n20471 = ( n14531 & n20469 ) | ( n14531 & n20470 ) | ( n20469 & n20470 ) ;
  assign n20472 = n3274 & n14352 ;
  assign n20473 = n20471 | n20472 ;
  assign n20474 = n1610 | n5638 ;
  assign n20475 = n2549 | n20474 ;
  assign n20476 = n599 | n1241 ;
  assign n20477 = n2105 | n20476 ;
  assign n20478 = n20475 | n20477 ;
  assign n20479 = n148 | n318 ;
  assign n20480 = n1092 | n20479 ;
  assign n20481 = n20478 | n20480 ;
  assign n20482 = n2222 | n5093 ;
  assign n20483 = n1292 | n20482 ;
  assign n20484 = n711 | n2544 ;
  assign n20485 = n20483 | n20484 ;
  assign n20486 = n364 | n871 ;
  assign n20487 = n4001 | n20486 ;
  assign n20488 = n20485 | n20487 ;
  assign n20489 = n2500 & ~n20488 ;
  assign n20490 = ~n20481 & n20489 ;
  assign n20491 = n765 | n988 ;
  assign n20492 = n1746 | n1937 ;
  assign n20493 = n20491 | n20492 ;
  assign n20494 = n20490 & ~n20493 ;
  assign n20495 = ~n3881 & n20494 ;
  assign n20496 = ~n4438 & n20495 ;
  assign n20497 = ( n20320 & ~n20473 ) | ( n20320 & n20496 ) | ( ~n20473 & n20496 ) ;
  assign n20498 = ( n20320 & n20473 ) | ( n20320 & ~n20496 ) | ( n20473 & ~n20496 ) ;
  assign n20499 = ( ~n20320 & n20497 ) | ( ~n20320 & n20498 ) | ( n20497 & n20498 ) ;
  assign n20500 = ( n20333 & n20466 ) | ( n20333 & ~n20499 ) | ( n20466 & ~n20499 ) ;
  assign n20501 = ( n20333 & ~n20466 ) | ( n20333 & n20499 ) | ( ~n20466 & n20499 ) ;
  assign n20502 = ( ~n20333 & n20500 ) | ( ~n20333 & n20501 ) | ( n20500 & n20501 ) ;
  assign n20503 = ( n20337 & n20456 ) | ( n20337 & ~n20502 ) | ( n20456 & ~n20502 ) ;
  assign n20504 = ( n20337 & ~n20456 ) | ( n20337 & n20502 ) | ( ~n20456 & n20502 ) ;
  assign n20505 = ( ~n20337 & n20503 ) | ( ~n20337 & n20504 ) | ( n20503 & n20504 ) ;
  assign n20506 = n4637 & ~n16150 ;
  assign n20507 = x23 & n20506 ;
  assign n20508 = n4584 & ~n15954 ;
  assign n20509 = n4649 | n20508 ;
  assign n20510 = ( ~n16338 & n20508 ) | ( ~n16338 & n20509 ) | ( n20508 & n20509 ) ;
  assign n20511 = n4591 | n20510 ;
  assign n20512 = ( ~n16349 & n20510 ) | ( ~n16349 & n20511 ) | ( n20510 & n20511 ) ;
  assign n20513 = x23 & ~n20512 ;
  assign n20514 = ( ~x23 & n20506 ) | ( ~x23 & n20512 ) | ( n20506 & n20512 ) ;
  assign n20515 = ( ~n20507 & n20513 ) | ( ~n20507 & n20514 ) | ( n20513 & n20514 ) ;
  assign n20516 = ( n20349 & ~n20505 ) | ( n20349 & n20515 ) | ( ~n20505 & n20515 ) ;
  assign n20517 = ( n20349 & n20505 ) | ( n20349 & ~n20515 ) | ( n20505 & ~n20515 ) ;
  assign n20518 = ( ~n20349 & n20516 ) | ( ~n20349 & n20517 ) | ( n20516 & n20517 ) ;
  assign n20519 = ( n20352 & n20446 ) | ( n20352 & ~n20518 ) | ( n20446 & ~n20518 ) ;
  assign n20520 = ( n20352 & ~n20446 ) | ( n20352 & n20518 ) | ( ~n20446 & n20518 ) ;
  assign n20521 = ( ~n20352 & n20519 ) | ( ~n20352 & n20520 ) | ( n20519 & n20520 ) ;
  assign n20522 = n5584 & n17346 ;
  assign n20523 = x17 & n20522 ;
  assign n20524 = n5413 & ~n17126 ;
  assign n20525 = n5417 | n20524 ;
  assign n20526 = ( ~n17635 & n20524 ) | ( ~n17635 & n20525 ) | ( n20524 & n20525 ) ;
  assign n20527 = n5418 | n20526 ;
  assign n20528 = ( ~n17646 & n20526 ) | ( ~n17646 & n20527 ) | ( n20526 & n20527 ) ;
  assign n20529 = x17 & ~n20528 ;
  assign n20530 = ( ~x17 & n20522 ) | ( ~x17 & n20528 ) | ( n20522 & n20528 ) ;
  assign n20531 = ( ~n20523 & n20529 ) | ( ~n20523 & n20530 ) | ( n20529 & n20530 ) ;
  assign n20532 = ( n20365 & ~n20521 ) | ( n20365 & n20531 ) | ( ~n20521 & n20531 ) ;
  assign n20533 = ( n20365 & n20521 ) | ( n20365 & ~n20531 ) | ( n20521 & ~n20531 ) ;
  assign n20534 = ( ~n20365 & n20532 ) | ( ~n20365 & n20533 ) | ( n20532 & n20533 ) ;
  assign n20535 = n6332 & ~n17963 ;
  assign n20536 = x14 & n20535 ;
  assign n20537 = n5909 & n17742 ;
  assign n20538 = n5914 | n20537 ;
  assign n20539 = ( ~n18258 & n20537 ) | ( ~n18258 & n20538 ) | ( n20537 & n20538 ) ;
  assign n20540 = n5915 | n20539 ;
  assign n20541 = ( n18268 & n20539 ) | ( n18268 & n20540 ) | ( n20539 & n20540 ) ;
  assign n20542 = x14 & ~n20541 ;
  assign n20543 = ( ~x14 & n20535 ) | ( ~x14 & n20541 ) | ( n20535 & n20541 ) ;
  assign n20544 = ( ~n20536 & n20542 ) | ( ~n20536 & n20543 ) | ( n20542 & n20543 ) ;
  assign n20545 = ( n20368 & ~n20534 ) | ( n20368 & n20544 ) | ( ~n20534 & n20544 ) ;
  assign n20546 = ( n20368 & n20534 ) | ( n20368 & ~n20544 ) | ( n20534 & ~n20544 ) ;
  assign n20547 = ( ~n20368 & n20545 ) | ( ~n20368 & n20546 ) | ( n20545 & n20546 ) ;
  assign n20548 = ( n20372 & n20436 ) | ( n20372 & ~n20547 ) | ( n20436 & ~n20547 ) ;
  assign n20549 = ( n20372 & ~n20436 ) | ( n20372 & n20547 ) | ( ~n20436 & n20547 ) ;
  assign n20550 = ( ~n20372 & n20548 ) | ( ~n20372 & n20549 ) | ( n20548 & n20549 ) ;
  assign n20551 = ( n20384 & n20426 ) | ( n20384 & ~n20550 ) | ( n20426 & ~n20550 ) ;
  assign n20552 = ( n20384 & ~n20426 ) | ( n20384 & n20550 ) | ( ~n20426 & n20550 ) ;
  assign n20553 = ( ~n20384 & n20551 ) | ( ~n20384 & n20552 ) | ( n20551 & n20552 ) ;
  assign n20554 = n40 & n19916 ;
  assign n20555 = n8721 & n19882 ;
  assign n20556 = n8340 & ~n19701 ;
  assign n20557 = n20555 | n20556 ;
  assign n20558 = n20554 | n20557 ;
  assign n20559 = x5 & n20558 ;
  assign n20560 = n8341 & n19920 ;
  assign n20561 = ( ~x5 & n20558 ) | ( ~x5 & n20560 ) | ( n20558 & n20560 ) ;
  assign n20562 = x5 & ~n20560 ;
  assign n20563 = ( ~n20559 & n20561 ) | ( ~n20559 & n20562 ) | ( n20561 & n20562 ) ;
  assign n20564 = ( n20398 & n20553 ) | ( n20398 & ~n20563 ) | ( n20553 & ~n20563 ) ;
  assign n20565 = ( n20398 & ~n20553 ) | ( n20398 & n20563 ) | ( ~n20553 & n20563 ) ;
  assign n20566 = ( ~n20398 & n20564 ) | ( ~n20398 & n20565 ) | ( n20564 & n20565 ) ;
  assign n20567 = ( x2 & n9590 ) | ( x2 & n20097 ) | ( n9590 & n20097 ) ;
  assign n20568 = n41 & ~n20095 ;
  assign n20569 = ( n9591 & ~n20097 ) | ( n9591 & n20568 ) | ( ~n20097 & n20568 ) ;
  assign n20570 = n20567 | n20569 ;
  assign n20571 = ~n9154 & n20091 ;
  assign n20572 = ( x2 & n20568 ) | ( x2 & n20571 ) | ( n20568 & n20571 ) ;
  assign n20573 = n20570 & ~n20572 ;
  assign n20574 = ( n20411 & ~n20566 ) | ( n20411 & n20573 ) | ( ~n20566 & n20573 ) ;
  assign n20575 = ( n20411 & n20566 ) | ( n20411 & ~n20573 ) | ( n20566 & ~n20573 ) ;
  assign n20576 = ( ~n20411 & n20574 ) | ( ~n20411 & n20575 ) | ( n20574 & n20575 ) ;
  assign n20577 = n20414 & ~n20576 ;
  assign n20578 = ~n20414 & n20576 ;
  assign n20579 = n20577 | n20578 ;
  assign n20580 = n8340 & n19882 ;
  assign n20581 = x5 & n20580 ;
  assign n20582 = n40 & n20091 ;
  assign n20583 = n8721 & n19916 ;
  assign n20584 = n20582 | n20583 ;
  assign n20585 = n8341 | n20584 ;
  assign n20586 = ( n20101 & n20584 ) | ( n20101 & n20585 ) | ( n20584 & n20585 ) ;
  assign n20587 = x5 & ~n20586 ;
  assign n20588 = ( ~x5 & n20580 ) | ( ~x5 & n20586 ) | ( n20580 & n20586 ) ;
  assign n20589 = ( ~n20581 & n20587 ) | ( ~n20581 & n20588 ) | ( n20587 & n20588 ) ;
  assign n20590 = n7341 & ~n19315 ;
  assign n20591 = n7345 | n20590 ;
  assign n20592 = ( ~n19701 & n20590 ) | ( ~n19701 & n20591 ) | ( n20590 & n20591 ) ;
  assign n20593 = n7644 & n19368 ;
  assign n20594 = n20592 | n20593 ;
  assign n20595 = x8 & n20594 ;
  assign n20596 = n7346 & ~n19706 ;
  assign n20597 = x8 & ~n20596 ;
  assign n20598 = ( ~x8 & n20594 ) | ( ~x8 & n20596 ) | ( n20594 & n20596 ) ;
  assign n20599 = ( ~n20595 & n20597 ) | ( ~n20595 & n20598 ) | ( n20597 & n20598 ) ;
  assign n20600 = n6796 & n19177 ;
  assign n20601 = x11 & n20600 ;
  assign n20602 = n6567 & n18730 ;
  assign n20603 = n6570 | n20602 ;
  assign n20604 = ( n19248 & n20602 ) | ( n19248 & n20603 ) | ( n20602 & n20603 ) ;
  assign n20605 = n6571 | n20604 ;
  assign n20606 = ( n19253 & n20604 ) | ( n19253 & n20605 ) | ( n20604 & n20605 ) ;
  assign n20607 = x11 & ~n20606 ;
  assign n20608 = ( ~x11 & n20600 ) | ( ~x11 & n20606 ) | ( n20600 & n20606 ) ;
  assign n20609 = ( ~n20601 & n20607 ) | ( ~n20601 & n20608 ) | ( n20607 & n20608 ) ;
  assign n20610 = n4215 & ~n15954 ;
  assign n20611 = n4200 & ~n15806 ;
  assign n20612 = n2083 & n15561 ;
  assign n20613 = n20611 | n20612 ;
  assign n20614 = n20610 | n20613 ;
  assign n20615 = x26 & n20614 ;
  assign n20616 = n4203 & ~n15965 ;
  assign n20617 = ( ~x26 & n20614 ) | ( ~x26 & n20616 ) | ( n20614 & n20616 ) ;
  assign n20618 = x26 & ~n20616 ;
  assign n20619 = ( ~n20615 & n20617 ) | ( ~n20615 & n20618 ) | ( n20617 & n20618 ) ;
  assign n20620 = n3501 & ~n15184 ;
  assign n20621 = x29 & n20620 ;
  assign n20622 = n3536 & n14942 ;
  assign n20623 = n4039 | n20622 ;
  assign n20624 = ( ~n15394 & n20622 ) | ( ~n15394 & n20623 ) | ( n20622 & n20623 ) ;
  assign n20625 = n3541 | n20624 ;
  assign n20626 = ( n15405 & n20624 ) | ( n15405 & n20625 ) | ( n20624 & n20625 ) ;
  assign n20627 = x29 & ~n20626 ;
  assign n20628 = ( ~x29 & n20620 ) | ( ~x29 & n20626 ) | ( n20620 & n20626 ) ;
  assign n20629 = ( ~n20621 & n20627 ) | ( ~n20621 & n20628 ) | ( n20627 & n20628 ) ;
  assign n20630 = n3273 & n14352 ;
  assign n20631 = n3270 | n20630 ;
  assign n20632 = ( ~n14723 & n20630 ) | ( ~n14723 & n20631 ) | ( n20630 & n20631 ) ;
  assign n20633 = n390 | n20632 ;
  assign n20634 = ( ~n14734 & n20632 ) | ( ~n14734 & n20633 ) | ( n20632 & n20633 ) ;
  assign n20635 = n3274 & n14520 ;
  assign n20636 = n20634 | n20635 ;
  assign n20637 = n791 | n3719 ;
  assign n20638 = n1331 | n12844 ;
  assign n20639 = n1224 | n20638 ;
  assign n20640 = n3546 | n3755 ;
  assign n20641 = n20639 | n20640 ;
  assign n20642 = n218 | n733 ;
  assign n20643 = n526 | n678 ;
  assign n20644 = n153 | n260 ;
  assign n20645 = n20643 | n20644 ;
  assign n20646 = n20642 | n20645 ;
  assign n20647 = n20641 | n20646 ;
  assign n20648 = n20637 | n20647 ;
  assign n20649 = n3780 | n20648 ;
  assign n20650 = n5126 | n20649 ;
  assign n20651 = n13224 & ~n20650 ;
  assign n20652 = ( n20498 & ~n20636 ) | ( n20498 & n20651 ) | ( ~n20636 & n20651 ) ;
  assign n20653 = ( n20498 & n20636 ) | ( n20498 & ~n20651 ) | ( n20636 & ~n20651 ) ;
  assign n20654 = ( ~n20498 & n20652 ) | ( ~n20498 & n20653 ) | ( n20652 & n20653 ) ;
  assign n20655 = ( n20500 & n20629 ) | ( n20500 & ~n20654 ) | ( n20629 & ~n20654 ) ;
  assign n20656 = ( n20500 & ~n20629 ) | ( n20500 & n20654 ) | ( ~n20629 & n20654 ) ;
  assign n20657 = ( ~n20500 & n20655 ) | ( ~n20500 & n20656 ) | ( n20655 & n20656 ) ;
  assign n20658 = ( n20503 & n20619 ) | ( n20503 & ~n20657 ) | ( n20619 & ~n20657 ) ;
  assign n20659 = ( n20503 & ~n20619 ) | ( n20503 & n20657 ) | ( ~n20619 & n20657 ) ;
  assign n20660 = ( ~n20503 & n20658 ) | ( ~n20503 & n20659 ) | ( n20658 & n20659 ) ;
  assign n20661 = n4637 & ~n16338 ;
  assign n20662 = x23 & n20661 ;
  assign n20663 = n4584 & ~n16150 ;
  assign n20664 = n4649 | n20663 ;
  assign n20665 = ( ~n16531 & n20663 ) | ( ~n16531 & n20664 ) | ( n20663 & n20664 ) ;
  assign n20666 = n4591 | n20665 ;
  assign n20667 = ( ~n16542 & n20665 ) | ( ~n16542 & n20666 ) | ( n20665 & n20666 ) ;
  assign n20668 = x23 & ~n20667 ;
  assign n20669 = ( ~x23 & n20661 ) | ( ~x23 & n20667 ) | ( n20661 & n20667 ) ;
  assign n20670 = ( ~n20662 & n20668 ) | ( ~n20662 & n20669 ) | ( n20668 & n20669 ) ;
  assign n20671 = ( n20516 & ~n20660 ) | ( n20516 & n20670 ) | ( ~n20660 & n20670 ) ;
  assign n20672 = ( n20516 & n20660 ) | ( n20516 & ~n20670 ) | ( n20660 & ~n20670 ) ;
  assign n20673 = ( ~n20516 & n20671 ) | ( ~n20516 & n20672 ) | ( n20671 & n20672 ) ;
  assign n20674 = n4879 & ~n17139 ;
  assign n20675 = x20 & n20674 ;
  assign n20676 = n4874 & n16724 ;
  assign n20677 = n4878 | n20676 ;
  assign n20678 = ( ~n17126 & n20676 ) | ( ~n17126 & n20677 ) | ( n20676 & n20677 ) ;
  assign n20679 = n5232 & n16925 ;
  assign n20680 = n20678 | n20679 ;
  assign n20681 = x20 & ~n20680 ;
  assign n20682 = ( ~x20 & n20674 ) | ( ~x20 & n20680 ) | ( n20674 & n20680 ) ;
  assign n20683 = ( ~n20675 & n20681 ) | ( ~n20675 & n20682 ) | ( n20681 & n20682 ) ;
  assign n20684 = ( n20519 & ~n20673 ) | ( n20519 & n20683 ) | ( ~n20673 & n20683 ) ;
  assign n20685 = ( n20519 & n20673 ) | ( n20519 & ~n20683 ) | ( n20673 & ~n20683 ) ;
  assign n20686 = ( ~n20519 & n20684 ) | ( ~n20519 & n20685 ) | ( n20684 & n20685 ) ;
  assign n20687 = n5418 & ~n17749 ;
  assign n20688 = x17 & n20687 ;
  assign n20689 = n5417 & n17742 ;
  assign n20690 = n5584 & ~n17635 ;
  assign n20691 = n5413 & n17346 ;
  assign n20692 = n20690 | n20691 ;
  assign n20693 = n20689 | n20692 ;
  assign n20694 = x17 & ~n20693 ;
  assign n20695 = ( ~x17 & n20687 ) | ( ~x17 & n20693 ) | ( n20687 & n20693 ) ;
  assign n20696 = ( ~n20688 & n20694 ) | ( ~n20688 & n20695 ) | ( n20694 & n20695 ) ;
  assign n20697 = ( n20532 & ~n20686 ) | ( n20532 & n20696 ) | ( ~n20686 & n20696 ) ;
  assign n20698 = ( n20532 & n20686 ) | ( n20532 & ~n20696 ) | ( n20686 & ~n20696 ) ;
  assign n20699 = ( ~n20532 & n20697 ) | ( ~n20532 & n20698 ) | ( n20697 & n20698 ) ;
  assign n20700 = n6332 & ~n18258 ;
  assign n20701 = x14 & n20700 ;
  assign n20702 = n5909 & ~n17963 ;
  assign n20703 = n5914 | n20702 ;
  assign n20704 = ( ~n18362 & n20702 ) | ( ~n18362 & n20703 ) | ( n20702 & n20703 ) ;
  assign n20705 = n5915 | n20704 ;
  assign n20706 = ( ~n18373 & n20704 ) | ( ~n18373 & n20705 ) | ( n20704 & n20705 ) ;
  assign n20707 = x14 & ~n20706 ;
  assign n20708 = ( ~x14 & n20700 ) | ( ~x14 & n20706 ) | ( n20700 & n20706 ) ;
  assign n20709 = ( ~n20701 & n20707 ) | ( ~n20701 & n20708 ) | ( n20707 & n20708 ) ;
  assign n20710 = ( n20545 & n20699 ) | ( n20545 & ~n20709 ) | ( n20699 & ~n20709 ) ;
  assign n20711 = ( n20545 & ~n20699 ) | ( n20545 & n20709 ) | ( ~n20699 & n20709 ) ;
  assign n20712 = ( ~n20545 & n20710 ) | ( ~n20545 & n20711 ) | ( n20710 & n20711 ) ;
  assign n20713 = ( n20548 & n20609 ) | ( n20548 & ~n20712 ) | ( n20609 & ~n20712 ) ;
  assign n20714 = ( n20548 & ~n20609 ) | ( n20548 & n20712 ) | ( ~n20609 & n20712 ) ;
  assign n20715 = ( ~n20548 & n20713 ) | ( ~n20548 & n20714 ) | ( n20713 & n20714 ) ;
  assign n20716 = ( n20551 & n20599 ) | ( n20551 & ~n20715 ) | ( n20599 & ~n20715 ) ;
  assign n20717 = ( n20551 & ~n20599 ) | ( n20551 & n20715 ) | ( ~n20599 & n20715 ) ;
  assign n20718 = ( ~n20551 & n20716 ) | ( ~n20551 & n20717 ) | ( n20716 & n20717 ) ;
  assign n20719 = ( n20565 & n20589 ) | ( n20565 & ~n20718 ) | ( n20589 & ~n20718 ) ;
  assign n20720 = ( n20565 & ~n20589 ) | ( n20565 & n20718 ) | ( ~n20589 & n20718 ) ;
  assign n20721 = ( ~n20565 & n20719 ) | ( ~n20565 & n20720 ) | ( n20719 & n20720 ) ;
  assign n20722 = ( x2 & n9155 ) | ( x2 & n20095 ) | ( n9155 & n20095 ) ;
  assign n20723 = ( n20574 & n20721 ) | ( n20574 & ~n20722 ) | ( n20721 & ~n20722 ) ;
  assign n20724 = ( n20574 & ~n20721 ) | ( n20574 & n20722 ) | ( ~n20721 & n20722 ) ;
  assign n20725 = ( ~n20574 & n20723 ) | ( ~n20574 & n20724 ) | ( n20723 & n20724 ) ;
  assign n20726 = n20577 & ~n20725 ;
  assign n20727 = ~n20577 & n20725 ;
  assign n20728 = n20726 | n20727 ;
  assign n20729 = n7644 & ~n19701 ;
  assign n20730 = x8 & n20729 ;
  assign n20731 = n7341 & n19368 ;
  assign n20732 = n7345 | n20731 ;
  assign n20733 = ( n19882 & n20731 ) | ( n19882 & n20732 ) | ( n20731 & n20732 ) ;
  assign n20734 = n7346 | n20733 ;
  assign n20735 = ( ~n19893 & n20733 ) | ( ~n19893 & n20734 ) | ( n20733 & n20734 ) ;
  assign n20736 = x8 & ~n20735 ;
  assign n20737 = ( ~x8 & n20729 ) | ( ~x8 & n20735 ) | ( n20729 & n20735 ) ;
  assign n20738 = ( ~n20730 & n20736 ) | ( ~n20730 & n20737 ) | ( n20736 & n20737 ) ;
  assign n20739 = n6796 & n19248 ;
  assign n20740 = x11 & n20739 ;
  assign n20741 = n6567 & n19177 ;
  assign n20742 = n6570 | n20741 ;
  assign n20743 = ( ~n19315 & n20741 ) | ( ~n19315 & n20742 ) | ( n20741 & n20742 ) ;
  assign n20744 = n6571 | n20743 ;
  assign n20745 = ( ~n19320 & n20743 ) | ( ~n19320 & n20744 ) | ( n20743 & n20744 ) ;
  assign n20746 = x11 & ~n20745 ;
  assign n20747 = ( ~x11 & n20739 ) | ( ~x11 & n20745 ) | ( n20739 & n20745 ) ;
  assign n20748 = ( ~n20740 & n20746 ) | ( ~n20740 & n20747 ) | ( n20746 & n20747 ) ;
  assign n20749 = n5914 & n18730 ;
  assign n20750 = n5915 | n20749 ;
  assign n20751 = ( n18735 & n20749 ) | ( n18735 & n20750 ) | ( n20749 & n20750 ) ;
  assign n20752 = n6332 & ~n18362 ;
  assign n20753 = n20751 | n20752 ;
  assign n20754 = n5908 & ~n18258 ;
  assign n20755 = n5909 & ~n18258 ;
  assign n20756 = x14 & ~n20755 ;
  assign n20757 = ( ~n20753 & n20754 ) | ( ~n20753 & n20756 ) | ( n20754 & n20756 ) ;
  assign n20758 = n20753 | n20756 ;
  assign n20759 = ( ~x14 & n20757 ) | ( ~x14 & n20758 ) | ( n20757 & n20758 ) ;
  assign n20760 = n5418 & ~n17976 ;
  assign n20761 = x17 & n20760 ;
  assign n20762 = n5417 & ~n17963 ;
  assign n20763 = n5584 & n17742 ;
  assign n20764 = n5413 & ~n17635 ;
  assign n20765 = n20763 | n20764 ;
  assign n20766 = n20762 | n20765 ;
  assign n20767 = x17 & ~n20766 ;
  assign n20768 = ( ~x17 & n20760 ) | ( ~x17 & n20766 ) | ( n20760 & n20766 ) ;
  assign n20769 = ( ~n20761 & n20767 ) | ( ~n20761 & n20768 ) | ( n20767 & n20768 ) ;
  assign n20770 = n4649 & n16724 ;
  assign n20771 = n4637 & ~n16531 ;
  assign n20772 = n4584 & ~n16338 ;
  assign n20773 = n20771 | n20772 ;
  assign n20774 = n20770 | n20773 ;
  assign n20775 = x23 & n20774 ;
  assign n20776 = n4591 & n16735 ;
  assign n20777 = ( ~x23 & n20774 ) | ( ~x23 & n20776 ) | ( n20774 & n20776 ) ;
  assign n20778 = x23 & ~n20776 ;
  assign n20779 = ( ~n20775 & n20777 ) | ( ~n20775 & n20778 ) | ( n20777 & n20778 ) ;
  assign n20780 = n3501 & ~n15394 ;
  assign n20781 = x29 & n20780 ;
  assign n20782 = n3536 & ~n15184 ;
  assign n20783 = n4039 | n20782 ;
  assign n20784 = ( n15561 & n20782 ) | ( n15561 & n20783 ) | ( n20782 & n20783 ) ;
  assign n20785 = n3541 | n20784 ;
  assign n20786 = ( n15573 & n20784 ) | ( n15573 & n20785 ) | ( n20784 & n20785 ) ;
  assign n20787 = x29 & ~n20786 ;
  assign n20788 = ( ~x29 & n20780 ) | ( ~x29 & n20786 ) | ( n20780 & n20786 ) ;
  assign n20789 = ( ~n20781 & n20787 ) | ( ~n20781 & n20788 ) | ( n20787 & n20788 ) ;
  assign n20790 = n3273 & n14520 ;
  assign n20791 = n3270 | n20790 ;
  assign n20792 = ( n14942 & n20790 ) | ( n14942 & n20791 ) | ( n20790 & n20791 ) ;
  assign n20793 = n390 | n20792 ;
  assign n20794 = ( ~n14953 & n20792 ) | ( ~n14953 & n20793 ) | ( n20792 & n20793 ) ;
  assign n20795 = n3274 & ~n14723 ;
  assign n20796 = n20794 | n20795 ;
  assign n20797 = n2886 | n14865 ;
  assign n20798 = n242 | n261 ;
  assign n20799 = n618 & ~n20798 ;
  assign n20800 = ~n1194 & n20799 ;
  assign n20801 = ~n15904 & n20800 ;
  assign n20802 = n2051 | n2214 ;
  assign n20803 = n4927 | n20802 ;
  assign n20804 = n420 | n3061 ;
  assign n20805 = n20803 | n20804 ;
  assign n20806 = n20801 & ~n20805 ;
  assign n20807 = n2792 | n4001 ;
  assign n20808 = n20806 & ~n20807 ;
  assign n20809 = ~n20797 & n20808 ;
  assign n20810 = n358 | n2003 ;
  assign n20811 = n786 | n1291 ;
  assign n20812 = n20810 | n20811 ;
  assign n20813 = n1675 | n20311 ;
  assign n20814 = n20812 | n20813 ;
  assign n20815 = n4912 | n20814 ;
  assign n20816 = n20809 & ~n20815 ;
  assign n20817 = ( n20653 & ~n20796 ) | ( n20653 & n20816 ) | ( ~n20796 & n20816 ) ;
  assign n20818 = ( n20653 & n20796 ) | ( n20653 & ~n20816 ) | ( n20796 & ~n20816 ) ;
  assign n20819 = ( ~n20653 & n20817 ) | ( ~n20653 & n20818 ) | ( n20817 & n20818 ) ;
  assign n20820 = ( n20655 & ~n20789 ) | ( n20655 & n20819 ) | ( ~n20789 & n20819 ) ;
  assign n20821 = ( n20655 & n20789 ) | ( n20655 & ~n20819 ) | ( n20789 & ~n20819 ) ;
  assign n20822 = ( ~n20655 & n20820 ) | ( ~n20655 & n20821 ) | ( n20820 & n20821 ) ;
  assign n20823 = n4215 & ~n16150 ;
  assign n20824 = n4200 & ~n15954 ;
  assign n20825 = n2083 & ~n15806 ;
  assign n20826 = n20824 | n20825 ;
  assign n20827 = n20823 | n20826 ;
  assign n20828 = x26 & n20827 ;
  assign n20829 = n4203 & ~n16161 ;
  assign n20830 = ( ~x26 & n20827 ) | ( ~x26 & n20829 ) | ( n20827 & n20829 ) ;
  assign n20831 = x26 & ~n20829 ;
  assign n20832 = ( ~n20828 & n20830 ) | ( ~n20828 & n20831 ) | ( n20830 & n20831 ) ;
  assign n20833 = ( n20658 & ~n20822 ) | ( n20658 & n20832 ) | ( ~n20822 & n20832 ) ;
  assign n20834 = ( n20658 & n20822 ) | ( n20658 & ~n20832 ) | ( n20822 & ~n20832 ) ;
  assign n20835 = ( ~n20658 & n20833 ) | ( ~n20658 & n20834 ) | ( n20833 & n20834 ) ;
  assign n20836 = ( n20671 & n20779 ) | ( n20671 & ~n20835 ) | ( n20779 & ~n20835 ) ;
  assign n20837 = ( n20671 & ~n20779 ) | ( n20671 & n20835 ) | ( ~n20779 & n20835 ) ;
  assign n20838 = ( ~n20671 & n20836 ) | ( ~n20671 & n20837 ) | ( n20836 & n20837 ) ;
  assign n20839 = n5232 & ~n17126 ;
  assign n20840 = x20 & n20839 ;
  assign n20841 = n4874 & n16925 ;
  assign n20842 = n4878 | n20841 ;
  assign n20843 = ( n17346 & n20841 ) | ( n17346 & n20842 ) | ( n20841 & n20842 ) ;
  assign n20844 = n4879 | n20843 ;
  assign n20845 = ( ~n17356 & n20843 ) | ( ~n17356 & n20844 ) | ( n20843 & n20844 ) ;
  assign n20846 = x20 & ~n20845 ;
  assign n20847 = ( ~x20 & n20839 ) | ( ~x20 & n20845 ) | ( n20839 & n20845 ) ;
  assign n20848 = ( ~n20840 & n20846 ) | ( ~n20840 & n20847 ) | ( n20846 & n20847 ) ;
  assign n20849 = ( n20684 & ~n20838 ) | ( n20684 & n20848 ) | ( ~n20838 & n20848 ) ;
  assign n20850 = ( n20684 & n20838 ) | ( n20684 & ~n20848 ) | ( n20838 & ~n20848 ) ;
  assign n20851 = ( ~n20684 & n20849 ) | ( ~n20684 & n20850 ) | ( n20849 & n20850 ) ;
  assign n20852 = ( n20697 & n20769 ) | ( n20697 & ~n20851 ) | ( n20769 & ~n20851 ) ;
  assign n20853 = ( n20697 & ~n20769 ) | ( n20697 & n20851 ) | ( ~n20769 & n20851 ) ;
  assign n20854 = ( ~n20697 & n20852 ) | ( ~n20697 & n20853 ) | ( n20852 & n20853 ) ;
  assign n20855 = ( n20711 & n20759 ) | ( n20711 & ~n20854 ) | ( n20759 & ~n20854 ) ;
  assign n20856 = ( n20711 & ~n20759 ) | ( n20711 & n20854 ) | ( ~n20759 & n20854 ) ;
  assign n20857 = ( ~n20711 & n20855 ) | ( ~n20711 & n20856 ) | ( n20855 & n20856 ) ;
  assign n20858 = ( n20713 & n20748 ) | ( n20713 & ~n20857 ) | ( n20748 & ~n20857 ) ;
  assign n20859 = ( n20713 & ~n20748 ) | ( n20713 & n20857 ) | ( ~n20748 & n20857 ) ;
  assign n20860 = ( ~n20713 & n20858 ) | ( ~n20713 & n20859 ) | ( n20858 & n20859 ) ;
  assign n20861 = ( n20716 & n20738 ) | ( n20716 & ~n20860 ) | ( n20738 & ~n20860 ) ;
  assign n20862 = ( n20716 & ~n20738 ) | ( n20716 & n20860 ) | ( ~n20738 & n20860 ) ;
  assign n20863 = ( ~n20716 & n20861 ) | ( ~n20716 & n20862 ) | ( n20861 & n20862 ) ;
  assign n20864 = n8340 & n19916 ;
  assign n20865 = x5 & n20864 ;
  assign n20866 = n40 & ~n20095 ;
  assign n20867 = n8721 & n20091 ;
  assign n20868 = n20866 | n20867 ;
  assign n20869 = n8341 & ~n20100 ;
  assign n20870 = n20868 | n20869 ;
  assign n20871 = x5 & ~n20870 ;
  assign n20872 = ( ~x5 & n20864 ) | ( ~x5 & n20870 ) | ( n20864 & n20870 ) ;
  assign n20873 = ( ~n20865 & n20871 ) | ( ~n20865 & n20872 ) | ( n20871 & n20872 ) ;
  assign n20874 = x2 | n20873 ;
  assign n20875 = x2 & n20873 ;
  assign n20876 = n20874 & ~n20875 ;
  assign n20877 = ( n20719 & n20863 ) | ( n20719 & ~n20876 ) | ( n20863 & ~n20876 ) ;
  assign n20878 = ( ~n20719 & n20863 ) | ( ~n20719 & n20876 ) | ( n20863 & n20876 ) ;
  assign n20879 = ( ~n20863 & n20877 ) | ( ~n20863 & n20878 ) | ( n20877 & n20878 ) ;
  assign n20880 = n20724 | n20879 ;
  assign n20881 = n20724 & n20879 ;
  assign n20882 = n20880 & ~n20881 ;
  assign n20883 = n20726 & ~n20882 ;
  assign n20884 = ~n20726 & n20882 ;
  assign n20885 = n20883 | n20884 ;
  assign n20886 = n8721 & ~n20095 ;
  assign n20887 = x5 & n20886 ;
  assign n20888 = n8340 & n20091 ;
  assign n20889 = n8341 | n20888 ;
  assign n20890 = ( ~n20097 & n20888 ) | ( ~n20097 & n20889 ) | ( n20888 & n20889 ) ;
  assign n20891 = x5 & ~n20890 ;
  assign n20892 = ( ~x5 & n20886 ) | ( ~x5 & n20890 ) | ( n20886 & n20890 ) ;
  assign n20893 = ( ~n20887 & n20891 ) | ( ~n20887 & n20892 ) | ( n20891 & n20892 ) ;
  assign n20894 = n7346 & n19920 ;
  assign n20895 = x8 & n20894 ;
  assign n20896 = n7341 & ~n19701 ;
  assign n20897 = n7345 | n20896 ;
  assign n20898 = ( n19916 & n20896 ) | ( n19916 & n20897 ) | ( n20896 & n20897 ) ;
  assign n20899 = n7644 & n19882 ;
  assign n20900 = n20898 | n20899 ;
  assign n20901 = x8 & ~n20900 ;
  assign n20902 = ( ~x8 & n20894 ) | ( ~x8 & n20900 ) | ( n20894 & n20900 ) ;
  assign n20903 = ( ~n20895 & n20901 ) | ( ~n20895 & n20902 ) | ( n20901 & n20902 ) ;
  assign n20904 = n6796 & ~n19315 ;
  assign n20905 = x11 & n20904 ;
  assign n20906 = n6567 & n19248 ;
  assign n20907 = n6570 | n20906 ;
  assign n20908 = ( n19368 & n20906 ) | ( n19368 & n20907 ) | ( n20906 & n20907 ) ;
  assign n20909 = n6571 | n20908 ;
  assign n20910 = ( ~n19374 & n20908 ) | ( ~n19374 & n20909 ) | ( n20908 & n20909 ) ;
  assign n20911 = x11 & ~n20910 ;
  assign n20912 = ( ~x11 & n20904 ) | ( ~x11 & n20910 ) | ( n20904 & n20910 ) ;
  assign n20913 = ( ~n20905 & n20911 ) | ( ~n20905 & n20912 ) | ( n20911 & n20912 ) ;
  assign n20914 = n5914 & n19177 ;
  assign n20915 = n6332 & n18730 ;
  assign n20916 = n5909 & ~n18362 ;
  assign n20917 = n20915 | n20916 ;
  assign n20918 = n20914 | n20917 ;
  assign n20919 = x14 & n20918 ;
  assign n20920 = n5915 & ~n19182 ;
  assign n20921 = ( ~x14 & n20918 ) | ( ~x14 & n20920 ) | ( n20918 & n20920 ) ;
  assign n20922 = x14 & ~n20920 ;
  assign n20923 = ( ~n20919 & n20921 ) | ( ~n20919 & n20922 ) | ( n20921 & n20922 ) ;
  assign n20924 = n5418 & n18268 ;
  assign n20925 = x17 & n20924 ;
  assign n20926 = n5413 & n17742 ;
  assign n20927 = n5417 | n20926 ;
  assign n20928 = ( ~n18258 & n20926 ) | ( ~n18258 & n20927 ) | ( n20926 & n20927 ) ;
  assign n20929 = n5584 & ~n17963 ;
  assign n20930 = n20928 | n20929 ;
  assign n20931 = x17 & ~n20930 ;
  assign n20932 = ( ~x17 & n20924 ) | ( ~x17 & n20930 ) | ( n20924 & n20930 ) ;
  assign n20933 = ( ~n20925 & n20931 ) | ( ~n20925 & n20932 ) | ( n20931 & n20932 ) ;
  assign n20934 = n4878 & ~n17635 ;
  assign n20935 = n5232 & n17346 ;
  assign n20936 = n4874 & ~n17126 ;
  assign n20937 = n20935 | n20936 ;
  assign n20938 = n20934 | n20937 ;
  assign n20939 = x20 & n20938 ;
  assign n20940 = n4879 & ~n17646 ;
  assign n20941 = ( ~x20 & n20938 ) | ( ~x20 & n20940 ) | ( n20938 & n20940 ) ;
  assign n20942 = x20 & ~n20940 ;
  assign n20943 = ( ~n20939 & n20941 ) | ( ~n20939 & n20942 ) | ( n20941 & n20942 ) ;
  assign n20944 = n4637 & n16724 ;
  assign n20945 = x23 & n20944 ;
  assign n20946 = n4584 & ~n16531 ;
  assign n20947 = n4649 | n20946 ;
  assign n20948 = ( n16925 & n20946 ) | ( n16925 & n20947 ) | ( n20946 & n20947 ) ;
  assign n20949 = n4591 | n20948 ;
  assign n20950 = ( ~n16936 & n20948 ) | ( ~n16936 & n20949 ) | ( n20948 & n20949 ) ;
  assign n20951 = x23 & ~n20950 ;
  assign n20952 = ( ~x23 & n20944 ) | ( ~x23 & n20950 ) | ( n20944 & n20950 ) ;
  assign n20953 = ( ~n20945 & n20951 ) | ( ~n20945 & n20952 ) | ( n20951 & n20952 ) ;
  assign n20954 = n3501 & n15561 ;
  assign n20955 = x29 & n20954 ;
  assign n20956 = n3536 & ~n15394 ;
  assign n20957 = n4039 | n20956 ;
  assign n20958 = ( ~n15806 & n20956 ) | ( ~n15806 & n20957 ) | ( n20956 & n20957 ) ;
  assign n20959 = n3541 | n20958 ;
  assign n20960 = ( n15817 & n20958 ) | ( n15817 & n20959 ) | ( n20958 & n20959 ) ;
  assign n20961 = x29 & ~n20960 ;
  assign n20962 = ( ~x29 & n20954 ) | ( ~x29 & n20960 ) | ( n20954 & n20960 ) ;
  assign n20963 = ( ~n20955 & n20961 ) | ( ~n20955 & n20962 ) | ( n20961 & n20962 ) ;
  assign n20964 = ~n6014 & n17933 ;
  assign n20965 = ~n3589 & n20964 ;
  assign n20966 = n842 | n999 ;
  assign n20967 = n5483 | n20966 ;
  assign n20968 = n2375 | n20967 ;
  assign n20969 = n876 | n2834 ;
  assign n20970 = n546 | n734 ;
  assign n20971 = n20969 | n20970 ;
  assign n20972 = n20968 | n20971 ;
  assign n20973 = n20965 & ~n20972 ;
  assign n20974 = n2482 | n17695 ;
  assign n20975 = n2529 | n20974 ;
  assign n20976 = n20973 & ~n20975 ;
  assign n20977 = ~n2904 & n20976 ;
  assign n20978 = ~n462 & n20977 ;
  assign n20979 = n390 & ~n15195 ;
  assign n20980 = n3270 & ~n15184 ;
  assign n20981 = n3274 & n14942 ;
  assign n20982 = n3273 & ~n14723 ;
  assign n20983 = n20981 | n20982 ;
  assign n20984 = n20980 | n20983 ;
  assign n20985 = n20979 | n20984 ;
  assign n20986 = ( x2 & n20978 ) | ( x2 & ~n20985 ) | ( n20978 & ~n20985 ) ;
  assign n20987 = ( ~x2 & n20978 ) | ( ~x2 & n20985 ) | ( n20978 & n20985 ) ;
  assign n20988 = ( ~n20978 & n20986 ) | ( ~n20978 & n20987 ) | ( n20986 & n20987 ) ;
  assign n20989 = ( ~n20818 & n20963 ) | ( ~n20818 & n20988 ) | ( n20963 & n20988 ) ;
  assign n20990 = ( n20818 & n20963 ) | ( n20818 & ~n20988 ) | ( n20963 & ~n20988 ) ;
  assign n20991 = ( ~n20963 & n20989 ) | ( ~n20963 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = n4215 & ~n16338 ;
  assign n20993 = n4200 & ~n16150 ;
  assign n20994 = n2083 & ~n15954 ;
  assign n20995 = n20993 | n20994 ;
  assign n20996 = n20992 | n20995 ;
  assign n20997 = x26 & n20996 ;
  assign n20998 = n4203 & ~n16349 ;
  assign n20999 = ( ~x26 & n20996 ) | ( ~x26 & n20998 ) | ( n20996 & n20998 ) ;
  assign n21000 = x26 & ~n20998 ;
  assign n21001 = ( ~n20997 & n20999 ) | ( ~n20997 & n21000 ) | ( n20999 & n21000 ) ;
  assign n21002 = ( n20821 & n20991 ) | ( n20821 & n21001 ) | ( n20991 & n21001 ) ;
  assign n21003 = ( n20821 & ~n20991 ) | ( n20821 & n21001 ) | ( ~n20991 & n21001 ) ;
  assign n21004 = ( n20991 & ~n21002 ) | ( n20991 & n21003 ) | ( ~n21002 & n21003 ) ;
  assign n21005 = ( ~n20833 & n20953 ) | ( ~n20833 & n21004 ) | ( n20953 & n21004 ) ;
  assign n21006 = ( n20833 & n20953 ) | ( n20833 & ~n21004 ) | ( n20953 & ~n21004 ) ;
  assign n21007 = ( ~n20953 & n21005 ) | ( ~n20953 & n21006 ) | ( n21005 & n21006 ) ;
  assign n21008 = ( ~n20836 & n20943 ) | ( ~n20836 & n21007 ) | ( n20943 & n21007 ) ;
  assign n21009 = ( n20836 & n20943 ) | ( n20836 & ~n21007 ) | ( n20943 & ~n21007 ) ;
  assign n21010 = ( ~n20943 & n21008 ) | ( ~n20943 & n21009 ) | ( n21008 & n21009 ) ;
  assign n21011 = ( n20849 & n20933 ) | ( n20849 & ~n21010 ) | ( n20933 & ~n21010 ) ;
  assign n21012 = ( n20849 & ~n20933 ) | ( n20849 & n21010 ) | ( ~n20933 & n21010 ) ;
  assign n21013 = ( ~n20849 & n21011 ) | ( ~n20849 & n21012 ) | ( n21011 & n21012 ) ;
  assign n21014 = ( n20852 & ~n20923 ) | ( n20852 & n21013 ) | ( ~n20923 & n21013 ) ;
  assign n21015 = ( n20852 & n20923 ) | ( n20852 & ~n21013 ) | ( n20923 & ~n21013 ) ;
  assign n21016 = ( ~n20852 & n21014 ) | ( ~n20852 & n21015 ) | ( n21014 & n21015 ) ;
  assign n21017 = ( n20855 & ~n20913 ) | ( n20855 & n21016 ) | ( ~n20913 & n21016 ) ;
  assign n21018 = ( n20855 & n20913 ) | ( n20855 & ~n21016 ) | ( n20913 & ~n21016 ) ;
  assign n21019 = ( ~n20855 & n21017 ) | ( ~n20855 & n21018 ) | ( n21017 & n21018 ) ;
  assign n21020 = ( ~n20858 & n20903 ) | ( ~n20858 & n21019 ) | ( n20903 & n21019 ) ;
  assign n21021 = ( n20858 & n20903 ) | ( n20858 & ~n21019 ) | ( n20903 & ~n21019 ) ;
  assign n21022 = ( ~n20903 & n21020 ) | ( ~n20903 & n21021 ) | ( n21020 & n21021 ) ;
  assign n21023 = ( n20861 & ~n20893 ) | ( n20861 & n21022 ) | ( ~n20893 & n21022 ) ;
  assign n21024 = ( n20861 & n20893 ) | ( n20861 & ~n21022 ) | ( n20893 & ~n21022 ) ;
  assign n21025 = ( ~n20861 & n21023 ) | ( ~n20861 & n21024 ) | ( n21023 & n21024 ) ;
  assign n21026 = ~n20863 & n20875 ;
  assign n21027 = ( x2 & ~n20863 ) | ( x2 & n20873 ) | ( ~n20863 & n20873 ) ;
  assign n21028 = n20724 & n21027 ;
  assign n21029 = ( n20719 & n21026 ) | ( n20719 & n21028 ) | ( n21026 & n21028 ) ;
  assign n21030 = n20863 & ~n20874 ;
  assign n21031 = n20724 | n21027 ;
  assign n21032 = ( n20719 & ~n21030 ) | ( n20719 & n21031 ) | ( ~n21030 & n21031 ) ;
  assign n21033 = ~n21025 & n21032 ;
  assign n21034 = n21029 | n21033 ;
  assign n21035 = ( n21029 & n21032 ) | ( n21029 & ~n21033 ) | ( n21032 & ~n21033 ) ;
  assign n21036 = ( n21025 & n21034 ) | ( n21025 & ~n21035 ) | ( n21034 & ~n21035 ) ;
  assign n21037 = n20883 & ~n21036 ;
  assign n21038 = ~n20883 & n21036 ;
  assign n21039 = n21037 | n21038 ;
  assign n21040 = n8336 | n20095 ;
  assign n21041 = x5 & ~n8338 ;
  assign n21042 = n20095 | n21041 ;
  assign n21043 = ( x5 & n21040 ) | ( x5 & ~n21042 ) | ( n21040 & ~n21042 ) ;
  assign n21044 = n7345 & n20091 ;
  assign n21045 = n7346 | n21044 ;
  assign n21046 = ( n20101 & n21044 ) | ( n20101 & n21045 ) | ( n21044 & n21045 ) ;
  assign n21047 = n7341 & n19882 ;
  assign n21048 = ( ~x8 & n21046 ) | ( ~x8 & n21047 ) | ( n21046 & n21047 ) ;
  assign n21049 = n7644 & n19916 ;
  assign n21050 = x8 & ~n21047 ;
  assign n21051 = n21049 | n21050 ;
  assign n21052 = ( n21046 & n21049 ) | ( n21046 & n21050 ) | ( n21049 & n21050 ) ;
  assign n21053 = ( n21048 & n21051 ) | ( n21048 & ~n21052 ) | ( n21051 & ~n21052 ) ;
  assign n21054 = n6796 & n19368 ;
  assign n21055 = x11 & n21054 ;
  assign n21056 = n6567 & ~n19315 ;
  assign n21057 = n6570 | n21056 ;
  assign n21058 = ( ~n19701 & n21056 ) | ( ~n19701 & n21057 ) | ( n21056 & n21057 ) ;
  assign n21059 = n6571 | n21058 ;
  assign n21060 = ( ~n19706 & n21058 ) | ( ~n19706 & n21059 ) | ( n21058 & n21059 ) ;
  assign n21061 = x11 & ~n21060 ;
  assign n21062 = ( ~x11 & n21054 ) | ( ~x11 & n21060 ) | ( n21054 & n21060 ) ;
  assign n21063 = ( ~n21055 & n21061 ) | ( ~n21055 & n21062 ) | ( n21061 & n21062 ) ;
  assign n21064 = n5915 & n19253 ;
  assign n21065 = x14 & n21064 ;
  assign n21066 = n5909 & n18730 ;
  assign n21067 = n5914 | n21066 ;
  assign n21068 = ( n19248 & n21066 ) | ( n19248 & n21067 ) | ( n21066 & n21067 ) ;
  assign n21069 = n6332 & n19177 ;
  assign n21070 = n21068 | n21069 ;
  assign n21071 = x14 & ~n21070 ;
  assign n21072 = ( ~x14 & n21064 ) | ( ~x14 & n21070 ) | ( n21064 & n21070 ) ;
  assign n21073 = ( ~n21065 & n21071 ) | ( ~n21065 & n21072 ) | ( n21071 & n21072 ) ;
  assign n21074 = n5584 & ~n18258 ;
  assign n21075 = x17 & n21074 ;
  assign n21076 = n5413 & ~n17963 ;
  assign n21077 = n5417 | n21076 ;
  assign n21078 = ( ~n18362 & n21076 ) | ( ~n18362 & n21077 ) | ( n21076 & n21077 ) ;
  assign n21079 = n5418 | n21078 ;
  assign n21080 = ( ~n18373 & n21078 ) | ( ~n18373 & n21079 ) | ( n21078 & n21079 ) ;
  assign n21081 = x17 & ~n21080 ;
  assign n21082 = ( ~x17 & n21074 ) | ( ~x17 & n21080 ) | ( n21074 & n21080 ) ;
  assign n21083 = ( ~n21075 & n21081 ) | ( ~n21075 & n21082 ) | ( n21081 & n21082 ) ;
  assign n21084 = n4879 & ~n17749 ;
  assign n21085 = x20 & n21084 ;
  assign n21086 = n4878 & n17742 ;
  assign n21087 = n5232 & ~n17635 ;
  assign n21088 = n4874 & n17346 ;
  assign n21089 = n21087 | n21088 ;
  assign n21090 = n21086 | n21089 ;
  assign n21091 = x20 & ~n21090 ;
  assign n21092 = ( ~x20 & n21084 ) | ( ~x20 & n21090 ) | ( n21084 & n21090 ) ;
  assign n21093 = ( ~n21085 & n21091 ) | ( ~n21085 & n21092 ) | ( n21091 & n21092 ) ;
  assign n21094 = n4637 & n16925 ;
  assign n21095 = x23 & n21094 ;
  assign n21096 = n4584 & n16724 ;
  assign n21097 = n4649 | n21096 ;
  assign n21098 = ( ~n17126 & n21096 ) | ( ~n17126 & n21097 ) | ( n21096 & n21097 ) ;
  assign n21099 = n4591 | n21098 ;
  assign n21100 = ( ~n17139 & n21098 ) | ( ~n17139 & n21099 ) | ( n21098 & n21099 ) ;
  assign n21101 = x23 & ~n21100 ;
  assign n21102 = ( ~x23 & n21094 ) | ( ~x23 & n21100 ) | ( n21094 & n21100 ) ;
  assign n21103 = ( ~n21095 & n21101 ) | ( ~n21095 & n21102 ) | ( n21101 & n21102 ) ;
  assign n21104 = n4215 & ~n16531 ;
  assign n21105 = n4200 & ~n16338 ;
  assign n21106 = n2083 & ~n16150 ;
  assign n21107 = n21105 | n21106 ;
  assign n21108 = n21104 | n21107 ;
  assign n21109 = x26 & n21108 ;
  assign n21110 = n4203 & ~n16542 ;
  assign n21111 = ( ~x26 & n21108 ) | ( ~x26 & n21110 ) | ( n21108 & n21110 ) ;
  assign n21112 = x26 & ~n21110 ;
  assign n21113 = ( ~n21109 & n21111 ) | ( ~n21109 & n21112 ) | ( n21111 & n21112 ) ;
  assign n21114 = n3037 | n6041 ;
  assign n21115 = n1971 | n18599 ;
  assign n21116 = n21114 | n21115 ;
  assign n21117 = n99 | n123 ;
  assign n21118 = n2321 | n21117 ;
  assign n21119 = n21116 | n21118 ;
  assign n21120 = n1130 | n1543 ;
  assign n21121 = n1658 | n21120 ;
  assign n21122 = n21119 | n21121 ;
  assign n21123 = n1199 | n2841 ;
  assign n21124 = n3563 | n3791 ;
  assign n21125 = n21123 | n21124 ;
  assign n21126 = n1916 | n21125 ;
  assign n21127 = n21122 | n21126 ;
  assign n21128 = n4806 | n12882 ;
  assign n21129 = n635 | n1332 ;
  assign n21130 = n408 | n21129 ;
  assign n21131 = n21128 | n21130 ;
  assign n21132 = n21127 | n21131 ;
  assign n21133 = n2600 | n12686 ;
  assign n21134 = n21132 | n21133 ;
  assign n21135 = ( n20978 & ~n20987 ) | ( n20978 & n21134 ) | ( ~n20987 & n21134 ) ;
  assign n21136 = ( n20978 & n20987 ) | ( n20978 & ~n21134 ) | ( n20987 & ~n21134 ) ;
  assign n21137 = ( ~n20978 & n21135 ) | ( ~n20978 & n21136 ) | ( n21135 & n21136 ) ;
  assign n21138 = n3273 & n14942 ;
  assign n21139 = n3270 | n21138 ;
  assign n21140 = ( ~n15394 & n21138 ) | ( ~n15394 & n21139 ) | ( n21138 & n21139 ) ;
  assign n21141 = n390 | n21140 ;
  assign n21142 = ( n15405 & n21140 ) | ( n15405 & n21141 ) | ( n21140 & n21141 ) ;
  assign n21143 = n3274 & ~n15184 ;
  assign n21144 = n21142 | n21143 ;
  assign n21145 = ( n20990 & n21137 ) | ( n20990 & n21144 ) | ( n21137 & n21144 ) ;
  assign n21146 = ( ~n20990 & n21137 ) | ( ~n20990 & n21144 ) | ( n21137 & n21144 ) ;
  assign n21147 = ( n20990 & ~n21145 ) | ( n20990 & n21146 ) | ( ~n21145 & n21146 ) ;
  assign n21148 = n3501 & ~n15806 ;
  assign n21149 = x29 & n21148 ;
  assign n21150 = n3536 & n15561 ;
  assign n21151 = n4039 | n21150 ;
  assign n21152 = ( ~n15954 & n21150 ) | ( ~n15954 & n21151 ) | ( n21150 & n21151 ) ;
  assign n21153 = n3541 | n21152 ;
  assign n21154 = ( ~n15965 & n21152 ) | ( ~n15965 & n21153 ) | ( n21152 & n21153 ) ;
  assign n21155 = x29 & ~n21154 ;
  assign n21156 = ( ~x29 & n21148 ) | ( ~x29 & n21154 ) | ( n21148 & n21154 ) ;
  assign n21157 = ( ~n21149 & n21155 ) | ( ~n21149 & n21156 ) | ( n21155 & n21156 ) ;
  assign n21158 = ( ~n21113 & n21147 ) | ( ~n21113 & n21157 ) | ( n21147 & n21157 ) ;
  assign n21159 = ( n21113 & n21147 ) | ( n21113 & n21157 ) | ( n21147 & n21157 ) ;
  assign n21160 = ( n21113 & n21158 ) | ( n21113 & ~n21159 ) | ( n21158 & ~n21159 ) ;
  assign n21161 = ( n21003 & ~n21103 ) | ( n21003 & n21160 ) | ( ~n21103 & n21160 ) ;
  assign n21162 = ( n21003 & n21103 ) | ( n21003 & n21160 ) | ( n21103 & n21160 ) ;
  assign n21163 = ( n21103 & n21161 ) | ( n21103 & ~n21162 ) | ( n21161 & ~n21162 ) ;
  assign n21164 = ( n21006 & n21093 ) | ( n21006 & n21163 ) | ( n21093 & n21163 ) ;
  assign n21165 = ( n21006 & ~n21093 ) | ( n21006 & n21163 ) | ( ~n21093 & n21163 ) ;
  assign n21166 = ( n21093 & ~n21164 ) | ( n21093 & n21165 ) | ( ~n21164 & n21165 ) ;
  assign n21167 = ( n21009 & ~n21083 ) | ( n21009 & n21166 ) | ( ~n21083 & n21166 ) ;
  assign n21168 = ( n21009 & n21083 ) | ( n21009 & n21166 ) | ( n21083 & n21166 ) ;
  assign n21169 = ( n21083 & n21167 ) | ( n21083 & ~n21168 ) | ( n21167 & ~n21168 ) ;
  assign n21170 = ( ~n21011 & n21073 ) | ( ~n21011 & n21169 ) | ( n21073 & n21169 ) ;
  assign n21171 = ( n21011 & n21073 ) | ( n21011 & n21169 ) | ( n21073 & n21169 ) ;
  assign n21172 = ( n21011 & n21170 ) | ( n21011 & ~n21171 ) | ( n21170 & ~n21171 ) ;
  assign n21173 = ( ~n21015 & n21063 ) | ( ~n21015 & n21172 ) | ( n21063 & n21172 ) ;
  assign n21174 = ( n21015 & n21063 ) | ( n21015 & n21172 ) | ( n21063 & n21172 ) ;
  assign n21175 = ( n21015 & n21173 ) | ( n21015 & ~n21174 ) | ( n21173 & ~n21174 ) ;
  assign n21176 = ( n21018 & ~n21053 ) | ( n21018 & n21175 ) | ( ~n21053 & n21175 ) ;
  assign n21177 = ( n21018 & n21053 ) | ( n21018 & n21175 ) | ( n21053 & n21175 ) ;
  assign n21178 = ( n21053 & n21176 ) | ( n21053 & ~n21177 ) | ( n21176 & ~n21177 ) ;
  assign n21179 = ( ~n21021 & n21043 ) | ( ~n21021 & n21178 ) | ( n21043 & n21178 ) ;
  assign n21180 = ( n21021 & n21043 ) | ( n21021 & n21178 ) | ( n21043 & n21178 ) ;
  assign n21181 = ( n21021 & n21179 ) | ( n21021 & ~n21180 ) | ( n21179 & ~n21180 ) ;
  assign n21182 = ( n21024 & n21034 ) | ( n21024 & n21181 ) | ( n21034 & n21181 ) ;
  assign n21183 = ( n21024 & ~n21034 ) | ( n21024 & n21181 ) | ( ~n21034 & n21181 ) ;
  assign n21184 = ( n21034 & ~n21182 ) | ( n21034 & n21183 ) | ( ~n21182 & n21183 ) ;
  assign n21185 = n21037 & n21184 ;
  assign n21186 = n21037 | n21184 ;
  assign n21187 = ~n21185 & n21186 ;
  assign n21188 = n7346 & ~n20100 ;
  assign n21189 = x8 & n21188 ;
  assign n21190 = n7341 & n19916 ;
  assign n21191 = n7345 | n21190 ;
  assign n21192 = ( ~n20095 & n21190 ) | ( ~n20095 & n21191 ) | ( n21190 & n21191 ) ;
  assign n21193 = n7644 & n20091 ;
  assign n21194 = n21192 | n21193 ;
  assign n21195 = x8 & ~n21194 ;
  assign n21196 = ( ~x8 & n21188 ) | ( ~x8 & n21194 ) | ( n21188 & n21194 ) ;
  assign n21197 = ( ~n21189 & n21195 ) | ( ~n21189 & n21196 ) | ( n21195 & n21196 ) ;
  assign n21198 = n6796 & ~n19701 ;
  assign n21199 = x11 & n21198 ;
  assign n21200 = n6567 & n19368 ;
  assign n21201 = n6570 | n21200 ;
  assign n21202 = ( n19882 & n21200 ) | ( n19882 & n21201 ) | ( n21200 & n21201 ) ;
  assign n21203 = n6571 | n21202 ;
  assign n21204 = ( ~n19893 & n21202 ) | ( ~n19893 & n21203 ) | ( n21202 & n21203 ) ;
  assign n21205 = x11 & ~n21204 ;
  assign n21206 = ( ~x11 & n21198 ) | ( ~x11 & n21204 ) | ( n21198 & n21204 ) ;
  assign n21207 = ( ~n21199 & n21205 ) | ( ~n21199 & n21206 ) | ( n21205 & n21206 ) ;
  assign n21208 = n6332 & n19248 ;
  assign n21209 = x14 & n21208 ;
  assign n21210 = n5909 & n19177 ;
  assign n21211 = n5914 | n21210 ;
  assign n21212 = ( ~n19315 & n21210 ) | ( ~n19315 & n21211 ) | ( n21210 & n21211 ) ;
  assign n21213 = n5915 | n21212 ;
  assign n21214 = ( ~n19320 & n21212 ) | ( ~n19320 & n21213 ) | ( n21212 & n21213 ) ;
  assign n21215 = x14 & ~n21214 ;
  assign n21216 = ( ~x14 & n21208 ) | ( ~x14 & n21214 ) | ( n21208 & n21214 ) ;
  assign n21217 = ( ~n21209 & n21215 ) | ( ~n21209 & n21216 ) | ( n21215 & n21216 ) ;
  assign n21218 = n5584 & ~n18362 ;
  assign n21219 = x17 & n21218 ;
  assign n21220 = n5413 & ~n18258 ;
  assign n21221 = n5417 | n21220 ;
  assign n21222 = ( n18730 & n21220 ) | ( n18730 & n21221 ) | ( n21220 & n21221 ) ;
  assign n21223 = n5418 | n21222 ;
  assign n21224 = ( n18735 & n21222 ) | ( n18735 & n21223 ) | ( n21222 & n21223 ) ;
  assign n21225 = x17 & ~n21224 ;
  assign n21226 = ( ~x17 & n21218 ) | ( ~x17 & n21224 ) | ( n21218 & n21224 ) ;
  assign n21227 = ( ~n21219 & n21225 ) | ( ~n21219 & n21226 ) | ( n21225 & n21226 ) ;
  assign n21228 = n4879 & ~n17976 ;
  assign n21229 = x20 & n21228 ;
  assign n21230 = n4878 & ~n17963 ;
  assign n21231 = n5232 & n17742 ;
  assign n21232 = n4874 & ~n17635 ;
  assign n21233 = n21231 | n21232 ;
  assign n21234 = n21230 | n21233 ;
  assign n21235 = x20 & ~n21234 ;
  assign n21236 = ( ~x20 & n21228 ) | ( ~x20 & n21234 ) | ( n21228 & n21234 ) ;
  assign n21237 = ( ~n21229 & n21235 ) | ( ~n21229 & n21236 ) | ( n21235 & n21236 ) ;
  assign n21238 = n4637 & ~n17126 ;
  assign n21239 = x23 & n21238 ;
  assign n21240 = n4584 & n16925 ;
  assign n21241 = n4649 | n21240 ;
  assign n21242 = ( n17346 & n21240 ) | ( n17346 & n21241 ) | ( n21240 & n21241 ) ;
  assign n21243 = n4591 | n21242 ;
  assign n21244 = ( ~n17356 & n21242 ) | ( ~n17356 & n21243 ) | ( n21242 & n21243 ) ;
  assign n21245 = x23 & ~n21244 ;
  assign n21246 = ( ~x23 & n21238 ) | ( ~x23 & n21244 ) | ( n21238 & n21244 ) ;
  assign n21247 = ( ~n21239 & n21245 ) | ( ~n21239 & n21246 ) | ( n21245 & n21246 ) ;
  assign n21248 = n4203 & n16735 ;
  assign n21249 = n4215 & n16724 ;
  assign n21250 = n4200 & ~n16531 ;
  assign n21251 = n2083 & ~n16338 ;
  assign n21252 = n21250 | n21251 ;
  assign n21253 = n21249 | n21252 ;
  assign n21254 = n21248 | n21253 ;
  assign n21255 = n4039 & ~n16150 ;
  assign n21256 = n3541 | n21255 ;
  assign n21257 = ( ~n16161 & n21255 ) | ( ~n16161 & n21256 ) | ( n21255 & n21256 ) ;
  assign n21258 = n3501 & ~n15954 ;
  assign n21259 = n21257 | n21258 ;
  assign n21260 = n3536 & ~n15806 ;
  assign n21261 = n21259 | n21260 ;
  assign n21262 = ( x26 & ~x29 ) | ( x26 & n21259 ) | ( ~x29 & n21259 ) ;
  assign n21263 = ( ~x26 & x29 ) | ( ~x26 & n21259 ) | ( x29 & n21259 ) ;
  assign n21264 = ( ~n21261 & n21262 ) | ( ~n21261 & n21263 ) | ( n21262 & n21263 ) ;
  assign n21265 = n3273 & ~n15184 ;
  assign n21266 = n3270 | n21265 ;
  assign n21267 = ( n15561 & n21265 ) | ( n15561 & n21266 ) | ( n21265 & n21266 ) ;
  assign n21268 = n390 | n21267 ;
  assign n21269 = ( n15573 & n21267 ) | ( n15573 & n21268 ) | ( n21267 & n21268 ) ;
  assign n21270 = n3274 & ~n15394 ;
  assign n21271 = n21269 | n21270 ;
  assign n21272 = x2 | n21134 ;
  assign n21273 = ( x2 & ~n20978 ) | ( x2 & n21272 ) | ( ~n20978 & n21272 ) ;
  assign n21274 = ( x2 & n20985 ) | ( x2 & n21273 ) | ( n20985 & n21273 ) ;
  assign n21275 = n329 | n463 ;
  assign n21276 = x23 & x25 ;
  assign n21277 = n98 & n21276 ;
  assign n21278 = n21275 | n21277 ;
  assign n21279 = n1702 | n21278 ;
  assign n21280 = n4756 | n21279 ;
  assign n21281 = n5018 | n21280 ;
  assign n21282 = n184 | n715 ;
  assign n21283 = n587 | n21282 ;
  assign n21284 = n3000 | n21283 ;
  assign n21285 = n2851 | n21284 ;
  assign n21286 = n3732 | n14883 ;
  assign n21287 = n21285 | n21286 ;
  assign n21288 = n21281 | n21287 ;
  assign n21289 = n1245 | n21288 ;
  assign n21290 = n2640 | n21289 ;
  assign n21291 = n1528 | n21290 ;
  assign n21292 = n21274 | n21291 ;
  assign n21293 = n20978 & ~n21134 ;
  assign n21294 = x2 & ~n21293 ;
  assign n21295 = ( x2 & n20985 ) | ( x2 & n21294 ) | ( n20985 & n21294 ) ;
  assign n21296 = ( ~n21274 & n21291 ) | ( ~n21274 & n21295 ) | ( n21291 & n21295 ) ;
  assign n21297 = n21291 | n21295 ;
  assign n21298 = ( n21292 & n21296 ) | ( n21292 & ~n21297 ) | ( n21296 & ~n21297 ) ;
  assign n21299 = ( n21145 & n21271 ) | ( n21145 & n21298 ) | ( n21271 & n21298 ) ;
  assign n21300 = ( ~n21145 & n21271 ) | ( ~n21145 & n21298 ) | ( n21271 & n21298 ) ;
  assign n21301 = ( n21145 & ~n21299 ) | ( n21145 & n21300 ) | ( ~n21299 & n21300 ) ;
  assign n21302 = ( ~n21254 & n21264 ) | ( ~n21254 & n21301 ) | ( n21264 & n21301 ) ;
  assign n21303 = ( n21254 & n21264 ) | ( n21254 & n21301 ) | ( n21264 & n21301 ) ;
  assign n21304 = ( n21254 & n21302 ) | ( n21254 & ~n21303 ) | ( n21302 & ~n21303 ) ;
  assign n21305 = ( n21159 & ~n21247 ) | ( n21159 & n21304 ) | ( ~n21247 & n21304 ) ;
  assign n21306 = ( n21159 & n21247 ) | ( n21159 & n21304 ) | ( n21247 & n21304 ) ;
  assign n21307 = ( n21247 & n21305 ) | ( n21247 & ~n21306 ) | ( n21305 & ~n21306 ) ;
  assign n21308 = ( ~n21162 & n21237 ) | ( ~n21162 & n21307 ) | ( n21237 & n21307 ) ;
  assign n21309 = ( n21162 & n21237 ) | ( n21162 & n21307 ) | ( n21237 & n21307 ) ;
  assign n21310 = ( n21162 & n21308 ) | ( n21162 & ~n21309 ) | ( n21308 & ~n21309 ) ;
  assign n21311 = ( ~n21164 & n21227 ) | ( ~n21164 & n21310 ) | ( n21227 & n21310 ) ;
  assign n21312 = ( n21164 & n21227 ) | ( n21164 & n21310 ) | ( n21227 & n21310 ) ;
  assign n21313 = ( n21164 & n21311 ) | ( n21164 & ~n21312 ) | ( n21311 & ~n21312 ) ;
  assign n21314 = ( ~n21168 & n21217 ) | ( ~n21168 & n21313 ) | ( n21217 & n21313 ) ;
  assign n21315 = ( n21168 & n21217 ) | ( n21168 & n21313 ) | ( n21217 & n21313 ) ;
  assign n21316 = ( n21168 & n21314 ) | ( n21168 & ~n21315 ) | ( n21314 & ~n21315 ) ;
  assign n21317 = ( n21171 & ~n21207 ) | ( n21171 & n21316 ) | ( ~n21207 & n21316 ) ;
  assign n21318 = ( n21171 & n21207 ) | ( n21171 & n21316 ) | ( n21207 & n21316 ) ;
  assign n21319 = ( n21207 & n21317 ) | ( n21207 & ~n21318 ) | ( n21317 & ~n21318 ) ;
  assign n21320 = ( n21174 & ~n21197 ) | ( n21174 & n21319 ) | ( ~n21197 & n21319 ) ;
  assign n21321 = ( n21174 & n21197 ) | ( n21174 & n21319 ) | ( n21197 & n21319 ) ;
  assign n21322 = ( n21197 & n21320 ) | ( n21197 & ~n21321 ) | ( n21320 & ~n21321 ) ;
  assign n21323 = ( x5 & ~n21177 ) | ( x5 & n21322 ) | ( ~n21177 & n21322 ) ;
  assign n21324 = ( x5 & n21177 ) | ( x5 & n21322 ) | ( n21177 & n21322 ) ;
  assign n21325 = ( n21177 & n21323 ) | ( n21177 & ~n21324 ) | ( n21323 & ~n21324 ) ;
  assign n21326 = ( n21180 & ~n21182 ) | ( n21180 & n21325 ) | ( ~n21182 & n21325 ) ;
  assign n21327 = ( n21180 & n21182 ) | ( n21180 & n21325 ) | ( n21182 & n21325 ) ;
  assign n21328 = ( n21182 & n21326 ) | ( n21182 & ~n21327 ) | ( n21326 & ~n21327 ) ;
  assign n21329 = n21185 & n21328 ;
  assign n21330 = n21185 | n21328 ;
  assign n21331 = ~n21329 & n21330 ;
  assign n21332 = n6796 & n19882 ;
  assign n21333 = x11 & n21332 ;
  assign n21334 = n6567 & ~n19701 ;
  assign n21335 = n6570 | n21334 ;
  assign n21336 = ( n19916 & n21334 ) | ( n19916 & n21335 ) | ( n21334 & n21335 ) ;
  assign n21337 = n6571 | n21336 ;
  assign n21338 = ( n19920 & n21336 ) | ( n19920 & n21337 ) | ( n21336 & n21337 ) ;
  assign n21339 = x11 & ~n21338 ;
  assign n21340 = ( ~x11 & n21332 ) | ( ~x11 & n21338 ) | ( n21332 & n21338 ) ;
  assign n21341 = ( ~n21333 & n21339 ) | ( ~n21333 & n21340 ) | ( n21339 & n21340 ) ;
  assign n21342 = n5915 & ~n19374 ;
  assign n21343 = x14 & n21342 ;
  assign n21344 = n5909 & n19248 ;
  assign n21345 = n5914 | n21344 ;
  assign n21346 = ( n19368 & n21344 ) | ( n19368 & n21345 ) | ( n21344 & n21345 ) ;
  assign n21347 = n6332 & ~n19315 ;
  assign n21348 = n21346 | n21347 ;
  assign n21349 = x14 & ~n21348 ;
  assign n21350 = ( ~x14 & n21342 ) | ( ~x14 & n21348 ) | ( n21342 & n21348 ) ;
  assign n21351 = ( ~n21343 & n21349 ) | ( ~n21343 & n21350 ) | ( n21349 & n21350 ) ;
  assign n21352 = n5584 & n18730 ;
  assign n21353 = x17 & n21352 ;
  assign n21354 = n5413 & ~n18362 ;
  assign n21355 = n5417 | n21354 ;
  assign n21356 = ( n19177 & n21354 ) | ( n19177 & n21355 ) | ( n21354 & n21355 ) ;
  assign n21357 = n5418 | n21356 ;
  assign n21358 = ( ~n19182 & n21356 ) | ( ~n19182 & n21357 ) | ( n21356 & n21357 ) ;
  assign n21359 = x17 & ~n21358 ;
  assign n21360 = ( ~x17 & n21352 ) | ( ~x17 & n21358 ) | ( n21352 & n21358 ) ;
  assign n21361 = ( ~n21353 & n21359 ) | ( ~n21353 & n21360 ) | ( n21359 & n21360 ) ;
  assign n21362 = n5232 & ~n17963 ;
  assign n21363 = x20 & n21362 ;
  assign n21364 = n4874 & n17742 ;
  assign n21365 = n4878 | n21364 ;
  assign n21366 = ( ~n18258 & n21364 ) | ( ~n18258 & n21365 ) | ( n21364 & n21365 ) ;
  assign n21367 = n4879 | n21366 ;
  assign n21368 = ( n18268 & n21366 ) | ( n18268 & n21367 ) | ( n21366 & n21367 ) ;
  assign n21369 = x20 & ~n21368 ;
  assign n21370 = ( ~x20 & n21362 ) | ( ~x20 & n21368 ) | ( n21362 & n21368 ) ;
  assign n21371 = ( ~n21363 & n21369 ) | ( ~n21363 & n21370 ) | ( n21369 & n21370 ) ;
  assign n21372 = n4637 & n17346 ;
  assign n21373 = x23 & n21372 ;
  assign n21374 = n4584 & ~n17126 ;
  assign n21375 = n4649 | n21374 ;
  assign n21376 = ( ~n17635 & n21374 ) | ( ~n17635 & n21375 ) | ( n21374 & n21375 ) ;
  assign n21377 = n4591 | n21376 ;
  assign n21378 = ( ~n17646 & n21376 ) | ( ~n17646 & n21377 ) | ( n21376 & n21377 ) ;
  assign n21379 = x23 & ~n21378 ;
  assign n21380 = ( ~x23 & n21372 ) | ( ~x23 & n21378 ) | ( n21372 & n21378 ) ;
  assign n21381 = ( ~n21373 & n21379 ) | ( ~n21373 & n21380 ) | ( n21379 & n21380 ) ;
  assign n21382 = x26 & ~n21254 ;
  assign n21383 = ~x26 & n21254 ;
  assign n21384 = n21382 | n21383 ;
  assign n21385 = x29 & ~n21261 ;
  assign n21386 = ~x29 & n21261 ;
  assign n21387 = n21385 | n21386 ;
  assign n21388 = ( n21301 & n21384 ) | ( n21301 & n21387 ) | ( n21384 & n21387 ) ;
  assign n21389 = n4215 & n16925 ;
  assign n21390 = n4200 & n16724 ;
  assign n21391 = n2083 & ~n16531 ;
  assign n21392 = n21390 | n21391 ;
  assign n21393 = n21389 | n21392 ;
  assign n21394 = x26 & n21393 ;
  assign n21395 = n4203 & ~n16936 ;
  assign n21396 = ( ~x26 & n21393 ) | ( ~x26 & n21395 ) | ( n21393 & n21395 ) ;
  assign n21397 = x26 & ~n21395 ;
  assign n21398 = ( ~n21394 & n21396 ) | ( ~n21394 & n21397 ) | ( n21396 & n21397 ) ;
  assign n21399 = n4039 & ~n16338 ;
  assign n21400 = n3541 | n21399 ;
  assign n21401 = ( ~n16349 & n21399 ) | ( ~n16349 & n21400 ) | ( n21399 & n21400 ) ;
  assign n21402 = n3536 & ~n15954 ;
  assign n21403 = ( ~x29 & n21401 ) | ( ~x29 & n21402 ) | ( n21401 & n21402 ) ;
  assign n21404 = n3501 & ~n16150 ;
  assign n21405 = x29 & ~n21402 ;
  assign n21406 = n21404 | n21405 ;
  assign n21407 = ( n21401 & n21404 ) | ( n21401 & n21405 ) | ( n21404 & n21405 ) ;
  assign n21408 = ( n21403 & n21406 ) | ( n21403 & ~n21407 ) | ( n21406 & ~n21407 ) ;
  assign n21409 = n3273 & ~n15394 ;
  assign n21410 = n3270 | n21409 ;
  assign n21411 = ( ~n15806 & n21409 ) | ( ~n15806 & n21410 ) | ( n21409 & n21410 ) ;
  assign n21412 = n390 | n21411 ;
  assign n21413 = ( n15817 & n21411 ) | ( n15817 & n21412 ) | ( n21411 & n21412 ) ;
  assign n21414 = n3274 & n15561 ;
  assign n21415 = n21413 | n21414 ;
  assign n21416 = n1292 | n4348 ;
  assign n21417 = n1780 | n2897 ;
  assign n21418 = n21416 | n21417 ;
  assign n21419 = n469 | n536 ;
  assign n21420 = n357 | n700 ;
  assign n21421 = n222 | n21420 ;
  assign n21422 = n4903 | n21421 ;
  assign n21423 = n21419 | n21422 ;
  assign n21424 = n21418 | n21423 ;
  assign n21425 = n17077 | n21424 ;
  assign n21426 = n18472 | n21425 ;
  assign n21427 = n4013 | n21426 ;
  assign n21428 = n2363 | n21427 ;
  assign n21429 = ( x2 & ~x5 ) | ( x2 & n21428 ) | ( ~x5 & n21428 ) ;
  assign n21430 = ( x2 & x5 ) | ( x2 & ~n21428 ) | ( x5 & ~n21428 ) ;
  assign n21431 = ( ~x2 & n21429 ) | ( ~x2 & n21430 ) | ( n21429 & n21430 ) ;
  assign n21432 = n21274 & n21297 ;
  assign n21433 = ( n21415 & n21431 ) | ( n21415 & n21432 ) | ( n21431 & n21432 ) ;
  assign n21434 = ( ~n21415 & n21431 ) | ( ~n21415 & n21432 ) | ( n21431 & n21432 ) ;
  assign n21435 = ( n21415 & ~n21433 ) | ( n21415 & n21434 ) | ( ~n21433 & n21434 ) ;
  assign n21436 = ( n21299 & n21408 ) | ( n21299 & n21435 ) | ( n21408 & n21435 ) ;
  assign n21437 = ( ~n21299 & n21408 ) | ( ~n21299 & n21435 ) | ( n21408 & n21435 ) ;
  assign n21438 = ( n21299 & ~n21436 ) | ( n21299 & n21437 ) | ( ~n21436 & n21437 ) ;
  assign n21439 = ( ~n21388 & n21398 ) | ( ~n21388 & n21438 ) | ( n21398 & n21438 ) ;
  assign n21440 = ( n21388 & n21398 ) | ( n21388 & n21438 ) | ( n21398 & n21438 ) ;
  assign n21441 = ( n21388 & n21439 ) | ( n21388 & ~n21440 ) | ( n21439 & ~n21440 ) ;
  assign n21442 = ( ~n21306 & n21381 ) | ( ~n21306 & n21441 ) | ( n21381 & n21441 ) ;
  assign n21443 = ( n21306 & n21381 ) | ( n21306 & n21441 ) | ( n21381 & n21441 ) ;
  assign n21444 = ( n21306 & n21442 ) | ( n21306 & ~n21443 ) | ( n21442 & ~n21443 ) ;
  assign n21445 = ( n21309 & ~n21371 ) | ( n21309 & n21444 ) | ( ~n21371 & n21444 ) ;
  assign n21446 = ( n21309 & n21371 ) | ( n21309 & n21444 ) | ( n21371 & n21444 ) ;
  assign n21447 = ( n21371 & n21445 ) | ( n21371 & ~n21446 ) | ( n21445 & ~n21446 ) ;
  assign n21448 = ( ~n21312 & n21361 ) | ( ~n21312 & n21447 ) | ( n21361 & n21447 ) ;
  assign n21449 = ( n21312 & n21361 ) | ( n21312 & n21447 ) | ( n21361 & n21447 ) ;
  assign n21450 = ( n21312 & n21448 ) | ( n21312 & ~n21449 ) | ( n21448 & ~n21449 ) ;
  assign n21451 = ( n21315 & ~n21351 ) | ( n21315 & n21450 ) | ( ~n21351 & n21450 ) ;
  assign n21452 = ( n21315 & n21351 ) | ( n21315 & n21450 ) | ( n21351 & n21450 ) ;
  assign n21453 = ( n21351 & n21451 ) | ( n21351 & ~n21452 ) | ( n21451 & ~n21452 ) ;
  assign n21454 = ( ~n21318 & n21341 ) | ( ~n21318 & n21453 ) | ( n21341 & n21453 ) ;
  assign n21455 = ( n21318 & n21341 ) | ( n21318 & n21453 ) | ( n21341 & n21453 ) ;
  assign n21456 = ( n21318 & n21454 ) | ( n21318 & ~n21455 ) | ( n21454 & ~n21455 ) ;
  assign n21457 = n7644 & ~n20095 ;
  assign n21458 = n7341 & n20091 ;
  assign n21459 = n21457 | n21458 ;
  assign n21460 = x8 & n21459 ;
  assign n21461 = n7346 & ~n20097 ;
  assign n21462 = ( ~x8 & n21459 ) | ( ~x8 & n21461 ) | ( n21459 & n21461 ) ;
  assign n21463 = x8 & ~n21461 ;
  assign n21464 = ( ~n21460 & n21462 ) | ( ~n21460 & n21463 ) | ( n21462 & n21463 ) ;
  assign n21465 = ( ~n21321 & n21456 ) | ( ~n21321 & n21464 ) | ( n21456 & n21464 ) ;
  assign n21466 = ( n21321 & n21456 ) | ( n21321 & n21464 ) | ( n21456 & n21464 ) ;
  assign n21467 = ( n21321 & n21465 ) | ( n21321 & ~n21466 ) | ( n21465 & ~n21466 ) ;
  assign n21468 = ( n21324 & n21327 ) | ( n21324 & n21467 ) | ( n21327 & n21467 ) ;
  assign n21469 = ( n21324 & ~n21327 ) | ( n21324 & n21467 ) | ( ~n21327 & n21467 ) ;
  assign n21470 = ( n21327 & ~n21468 ) | ( n21327 & n21469 ) | ( ~n21468 & n21469 ) ;
  assign n21471 = n21329 & ~n21470 ;
  assign n21472 = n21329 & n21470 ;
  assign n21473 = ( n21470 & n21471 ) | ( n21470 & ~n21472 ) | ( n21471 & ~n21472 ) ;
  assign n21474 = n6796 & n19916 ;
  assign n21475 = x11 & n21474 ;
  assign n21476 = n6567 & n19882 ;
  assign n21477 = n6570 | n21476 ;
  assign n21478 = ( n20091 & n21476 ) | ( n20091 & n21477 ) | ( n21476 & n21477 ) ;
  assign n21479 = n6571 | n21478 ;
  assign n21480 = ( n20101 & n21478 ) | ( n20101 & n21479 ) | ( n21478 & n21479 ) ;
  assign n21481 = x11 & ~n21480 ;
  assign n21482 = ( ~x11 & n21474 ) | ( ~x11 & n21480 ) | ( n21474 & n21480 ) ;
  assign n21483 = ( ~n21475 & n21481 ) | ( ~n21475 & n21482 ) | ( n21481 & n21482 ) ;
  assign n21484 = n5914 & ~n19701 ;
  assign n21485 = n5915 | n21484 ;
  assign n21486 = ( ~n19706 & n21484 ) | ( ~n19706 & n21485 ) | ( n21484 & n21485 ) ;
  assign n21487 = n6332 & n19368 ;
  assign n21488 = n21486 | n21487 ;
  assign n21489 = n5908 & ~n19315 ;
  assign n21490 = n5909 & ~n19315 ;
  assign n21491 = x14 & ~n21490 ;
  assign n21492 = ( ~n21488 & n21489 ) | ( ~n21488 & n21491 ) | ( n21489 & n21491 ) ;
  assign n21493 = n21488 | n21491 ;
  assign n21494 = ( ~x14 & n21492 ) | ( ~x14 & n21493 ) | ( n21492 & n21493 ) ;
  assign n21495 = n5584 & n19177 ;
  assign n21496 = x17 & n21495 ;
  assign n21497 = n5413 & n18730 ;
  assign n21498 = n5417 | n21497 ;
  assign n21499 = ( n19248 & n21497 ) | ( n19248 & n21498 ) | ( n21497 & n21498 ) ;
  assign n21500 = n5418 | n21499 ;
  assign n21501 = ( n19253 & n21499 ) | ( n19253 & n21500 ) | ( n21499 & n21500 ) ;
  assign n21502 = x17 & ~n21501 ;
  assign n21503 = ( ~x17 & n21495 ) | ( ~x17 & n21501 ) | ( n21495 & n21501 ) ;
  assign n21504 = ( ~n21496 & n21502 ) | ( ~n21496 & n21503 ) | ( n21502 & n21503 ) ;
  assign n21505 = n5232 & ~n18258 ;
  assign n21506 = x20 & n21505 ;
  assign n21507 = n4874 & ~n17963 ;
  assign n21508 = n4878 | n21507 ;
  assign n21509 = ( ~n18362 & n21507 ) | ( ~n18362 & n21508 ) | ( n21507 & n21508 ) ;
  assign n21510 = n4879 | n21509 ;
  assign n21511 = ( ~n18373 & n21509 ) | ( ~n18373 & n21510 ) | ( n21509 & n21510 ) ;
  assign n21512 = x20 & ~n21511 ;
  assign n21513 = ( ~x20 & n21505 ) | ( ~x20 & n21511 ) | ( n21505 & n21511 ) ;
  assign n21514 = ( ~n21506 & n21512 ) | ( ~n21506 & n21513 ) | ( n21512 & n21513 ) ;
  assign n21515 = n4649 & n17742 ;
  assign n21516 = x23 & n21515 ;
  assign n21517 = n4637 & ~n17635 ;
  assign n21518 = n4584 & n17346 ;
  assign n21519 = n21517 | n21518 ;
  assign n21520 = n4591 | n21519 ;
  assign n21521 = ( ~n17749 & n21519 ) | ( ~n17749 & n21520 ) | ( n21519 & n21520 ) ;
  assign n21522 = x23 & ~n21521 ;
  assign n21523 = ( ~x23 & n21515 ) | ( ~x23 & n21521 ) | ( n21515 & n21521 ) ;
  assign n21524 = ( ~n21516 & n21522 ) | ( ~n21516 & n21523 ) | ( n21522 & n21523 ) ;
  assign n21525 = n4215 & ~n17126 ;
  assign n21526 = n4200 & n16925 ;
  assign n21527 = n2083 & n16724 ;
  assign n21528 = n21526 | n21527 ;
  assign n21529 = n21525 | n21528 ;
  assign n21530 = x26 & n21529 ;
  assign n21531 = n4203 & ~n17139 ;
  assign n21532 = ( ~x26 & n21529 ) | ( ~x26 & n21531 ) | ( n21529 & n21531 ) ;
  assign n21533 = x26 & ~n21531 ;
  assign n21534 = ( ~n21530 & n21532 ) | ( ~n21530 & n21533 ) | ( n21532 & n21533 ) ;
  assign n21535 = n3541 & ~n16542 ;
  assign n21536 = x29 & n21535 ;
  assign n21537 = n3536 & ~n16150 ;
  assign n21538 = n4039 | n21537 ;
  assign n21539 = ( ~n16531 & n21537 ) | ( ~n16531 & n21538 ) | ( n21537 & n21538 ) ;
  assign n21540 = n3501 & ~n16338 ;
  assign n21541 = n21539 | n21540 ;
  assign n21542 = x29 & ~n21541 ;
  assign n21543 = ( ~x29 & n21535 ) | ( ~x29 & n21541 ) | ( n21535 & n21541 ) ;
  assign n21544 = ( ~n21536 & n21542 ) | ( ~n21536 & n21543 ) | ( n21542 & n21543 ) ;
  assign n21545 = n4286 | n5988 ;
  assign n21546 = n13414 | n21545 ;
  assign n21547 = n1329 | n21546 ;
  assign n21548 = n129 | n198 ;
  assign n21549 = n97 | n21548 ;
  assign n21550 = n1007 | n21549 ;
  assign n21551 = n3025 | n3072 ;
  assign n21552 = n21550 | n21551 ;
  assign n21553 = n1102 | n3905 ;
  assign n21554 = n221 | n794 ;
  assign n21555 = n1113 | n21554 ;
  assign n21556 = n21553 | n21555 ;
  assign n21557 = n21552 | n21556 ;
  assign n21558 = n21547 | n21557 ;
  assign n21559 = n2013 | n21558 ;
  assign n21560 = n1281 | n21559 ;
  assign n21561 = n982 | n1130 ;
  assign n21562 = n1149 | n1835 ;
  assign n21563 = n21561 | n21562 ;
  assign n21564 = n485 | n689 ;
  assign n21565 = n5635 | n21564 ;
  assign n21566 = n403 | n1126 ;
  assign n21567 = n1926 | n2836 ;
  assign n21568 = n21566 | n21567 ;
  assign n21569 = n21565 | n21568 ;
  assign n21570 = n6011 | n21569 ;
  assign n21571 = n21563 | n21570 ;
  assign n21572 = n21560 | n21571 ;
  assign n21573 = n3273 & n15561 ;
  assign n21574 = n3270 | n21573 ;
  assign n21575 = ( ~n15954 & n21573 ) | ( ~n15954 & n21574 ) | ( n21573 & n21574 ) ;
  assign n21576 = n390 | n21575 ;
  assign n21577 = ( ~n15965 & n21575 ) | ( ~n15965 & n21576 ) | ( n21575 & n21576 ) ;
  assign n21578 = n3274 & ~n15806 ;
  assign n21579 = n21577 | n21578 ;
  assign n21580 = ( n21430 & n21572 ) | ( n21430 & n21579 ) | ( n21572 & n21579 ) ;
  assign n21581 = ( n21430 & ~n21572 ) | ( n21430 & n21579 ) | ( ~n21572 & n21579 ) ;
  assign n21582 = ( n21572 & ~n21580 ) | ( n21572 & n21581 ) | ( ~n21580 & n21581 ) ;
  assign n21583 = ( ~n21433 & n21544 ) | ( ~n21433 & n21582 ) | ( n21544 & n21582 ) ;
  assign n21584 = ( n21433 & n21544 ) | ( n21433 & n21582 ) | ( n21544 & n21582 ) ;
  assign n21585 = ( n21433 & n21583 ) | ( n21433 & ~n21584 ) | ( n21583 & ~n21584 ) ;
  assign n21586 = ( n21436 & ~n21534 ) | ( n21436 & n21585 ) | ( ~n21534 & n21585 ) ;
  assign n21587 = ( n21436 & n21534 ) | ( n21436 & n21585 ) | ( n21534 & n21585 ) ;
  assign n21588 = ( n21534 & n21586 ) | ( n21534 & ~n21587 ) | ( n21586 & ~n21587 ) ;
  assign n21589 = ( n21440 & n21524 ) | ( n21440 & n21588 ) | ( n21524 & n21588 ) ;
  assign n21590 = ( n21440 & ~n21524 ) | ( n21440 & n21588 ) | ( ~n21524 & n21588 ) ;
  assign n21591 = ( n21524 & ~n21589 ) | ( n21524 & n21590 ) | ( ~n21589 & n21590 ) ;
  assign n21592 = ( n21443 & ~n21514 ) | ( n21443 & n21591 ) | ( ~n21514 & n21591 ) ;
  assign n21593 = ( n21443 & n21514 ) | ( n21443 & n21591 ) | ( n21514 & n21591 ) ;
  assign n21594 = ( n21514 & n21592 ) | ( n21514 & ~n21593 ) | ( n21592 & ~n21593 ) ;
  assign n21595 = ( n21446 & ~n21504 ) | ( n21446 & n21594 ) | ( ~n21504 & n21594 ) ;
  assign n21596 = ( n21446 & n21504 ) | ( n21446 & n21594 ) | ( n21504 & n21594 ) ;
  assign n21597 = ( n21504 & n21595 ) | ( n21504 & ~n21596 ) | ( n21595 & ~n21596 ) ;
  assign n21598 = ( n21449 & ~n21494 ) | ( n21449 & n21597 ) | ( ~n21494 & n21597 ) ;
  assign n21599 = ( n21449 & n21494 ) | ( n21449 & n21597 ) | ( n21494 & n21597 ) ;
  assign n21600 = ( n21494 & n21598 ) | ( n21494 & ~n21599 ) | ( n21598 & ~n21599 ) ;
  assign n21601 = ( n21452 & n21483 ) | ( n21452 & n21600 ) | ( n21483 & n21600 ) ;
  assign n21602 = ( n21452 & ~n21483 ) | ( n21452 & n21600 ) | ( ~n21483 & n21600 ) ;
  assign n21603 = ( n21483 & ~n21601 ) | ( n21483 & n21602 ) | ( ~n21601 & n21602 ) ;
  assign n21604 = n7336 & ~n20095 ;
  assign n21605 = n7340 | n20095 ;
  assign n21606 = ( x8 & n21604 ) | ( x8 & n21605 ) | ( n21604 & n21605 ) ;
  assign n21607 = ( n21455 & ~n21603 ) | ( n21455 & n21606 ) | ( ~n21603 & n21606 ) ;
  assign n21608 = ( n21455 & n21603 ) | ( n21455 & n21606 ) | ( n21603 & n21606 ) ;
  assign n21609 = ( n21603 & n21607 ) | ( n21603 & ~n21608 ) | ( n21607 & ~n21608 ) ;
  assign n21610 = ( n21466 & ~n21468 ) | ( n21466 & n21609 ) | ( ~n21468 & n21609 ) ;
  assign n21611 = ( n21466 & n21468 ) | ( n21466 & n21609 ) | ( n21468 & n21609 ) ;
  assign n21612 = ( n21468 & n21610 ) | ( n21468 & ~n21611 ) | ( n21610 & ~n21611 ) ;
  assign n21613 = n21472 & ~n21612 ;
  assign n21614 = n21472 & n21612 ;
  assign n21615 = ( n21612 & n21613 ) | ( n21612 & ~n21614 ) | ( n21613 & ~n21614 ) ;
  assign n21616 = n6567 & n19916 ;
  assign n21617 = n6570 | n21616 ;
  assign n21618 = ( ~n20095 & n21616 ) | ( ~n20095 & n21617 ) | ( n21616 & n21617 ) ;
  assign n21619 = n6796 & n20091 ;
  assign n21620 = n21618 | n21619 ;
  assign n21621 = x11 & n21620 ;
  assign n21622 = n6571 & ~n20100 ;
  assign n21623 = ( ~x11 & n21620 ) | ( ~x11 & n21622 ) | ( n21620 & n21622 ) ;
  assign n21624 = x11 & ~n21622 ;
  assign n21625 = ( ~n21621 & n21623 ) | ( ~n21621 & n21624 ) | ( n21623 & n21624 ) ;
  assign n21626 = n6332 & ~n19701 ;
  assign n21627 = x14 & n21626 ;
  assign n21628 = n5909 & n19368 ;
  assign n21629 = n5914 | n21628 ;
  assign n21630 = ( n19882 & n21628 ) | ( n19882 & n21629 ) | ( n21628 & n21629 ) ;
  assign n21631 = n5915 | n21630 ;
  assign n21632 = ( ~n19893 & n21630 ) | ( ~n19893 & n21631 ) | ( n21630 & n21631 ) ;
  assign n21633 = x14 & ~n21632 ;
  assign n21634 = ( ~x14 & n21626 ) | ( ~x14 & n21632 ) | ( n21626 & n21632 ) ;
  assign n21635 = ( ~n21627 & n21633 ) | ( ~n21627 & n21634 ) | ( n21633 & n21634 ) ;
  assign n21636 = n5584 & n19248 ;
  assign n21637 = x17 & n21636 ;
  assign n21638 = n5413 & n19177 ;
  assign n21639 = n5417 | n21638 ;
  assign n21640 = ( ~n19315 & n21638 ) | ( ~n19315 & n21639 ) | ( n21638 & n21639 ) ;
  assign n21641 = n5418 | n21640 ;
  assign n21642 = ( ~n19320 & n21640 ) | ( ~n19320 & n21641 ) | ( n21640 & n21641 ) ;
  assign n21643 = x17 & ~n21642 ;
  assign n21644 = ( ~x17 & n21636 ) | ( ~x17 & n21642 ) | ( n21636 & n21642 ) ;
  assign n21645 = ( ~n21637 & n21643 ) | ( ~n21637 & n21644 ) | ( n21643 & n21644 ) ;
  assign n21646 = n5232 & ~n18362 ;
  assign n21647 = x20 & n21646 ;
  assign n21648 = n4874 & ~n18258 ;
  assign n21649 = n4878 | n21648 ;
  assign n21650 = ( n18730 & n21648 ) | ( n18730 & n21649 ) | ( n21648 & n21649 ) ;
  assign n21651 = n4879 | n21650 ;
  assign n21652 = ( n18735 & n21650 ) | ( n18735 & n21651 ) | ( n21650 & n21651 ) ;
  assign n21653 = x20 & ~n21652 ;
  assign n21654 = ( ~x20 & n21646 ) | ( ~x20 & n21652 ) | ( n21646 & n21652 ) ;
  assign n21655 = ( ~n21647 & n21653 ) | ( ~n21647 & n21654 ) | ( n21653 & n21654 ) ;
  assign n21656 = n4591 & ~n17976 ;
  assign n21657 = x23 & n21656 ;
  assign n21658 = n4649 & ~n17963 ;
  assign n21659 = n4637 & n17742 ;
  assign n21660 = n4584 & ~n17635 ;
  assign n21661 = n21659 | n21660 ;
  assign n21662 = n21658 | n21661 ;
  assign n21663 = x23 & ~n21662 ;
  assign n21664 = ( ~x23 & n21656 ) | ( ~x23 & n21662 ) | ( n21656 & n21662 ) ;
  assign n21665 = ( ~n21657 & n21663 ) | ( ~n21657 & n21664 ) | ( n21663 & n21664 ) ;
  assign n21666 = n4215 & n17346 ;
  assign n21667 = n4200 & ~n17126 ;
  assign n21668 = n2083 & n16925 ;
  assign n21669 = n21667 | n21668 ;
  assign n21670 = n21666 | n21669 ;
  assign n21671 = x26 & n21670 ;
  assign n21672 = n4203 & ~n17356 ;
  assign n21673 = ( ~x26 & n21670 ) | ( ~x26 & n21672 ) | ( n21670 & n21672 ) ;
  assign n21674 = x26 & ~n21672 ;
  assign n21675 = ( ~n21671 & n21673 ) | ( ~n21671 & n21674 ) | ( n21673 & n21674 ) ;
  assign n21676 = n4039 & n16724 ;
  assign n21677 = n3501 & ~n16531 ;
  assign n21678 = n3536 & ~n16338 ;
  assign n21679 = n21677 | n21678 ;
  assign n21680 = n21676 | n21679 ;
  assign n21681 = x29 & n21680 ;
  assign n21682 = n3541 & n16735 ;
  assign n21683 = ( ~x29 & n21680 ) | ( ~x29 & n21682 ) | ( n21680 & n21682 ) ;
  assign n21684 = x29 & ~n21682 ;
  assign n21685 = ( ~n21681 & n21683 ) | ( ~n21681 & n21684 ) | ( n21683 & n21684 ) ;
  assign n21686 = n329 | n616 ;
  assign n21687 = n2629 | n21686 ;
  assign n21688 = n5140 | n21687 ;
  assign n21689 = n3223 | n6118 ;
  assign n21690 = n21688 | n21689 ;
  assign n21691 = n17682 | n21690 ;
  assign n21692 = n4018 | n21691 ;
  assign n21693 = n3808 | n21692 ;
  assign n21694 = n471 | n679 ;
  assign n21695 = n226 | n21694 ;
  assign n21696 = n5974 | n21695 ;
  assign n21697 = n745 | n1542 ;
  assign n21698 = n21696 | n21697 ;
  assign n21699 = n1556 | n21698 ;
  assign n21700 = n325 | n4382 ;
  assign n21701 = n2850 | n2866 ;
  assign n21702 = n21700 | n21701 ;
  assign n21703 = n2844 & ~n21702 ;
  assign n21704 = ~n21699 & n21703 ;
  assign n21705 = n185 | n465 ;
  assign n21706 = n308 | n21705 ;
  assign n21707 = n661 | n750 ;
  assign n21708 = n21706 | n21707 ;
  assign n21709 = n318 | n912 ;
  assign n21710 = n592 | n21709 ;
  assign n21711 = n21708 | n21710 ;
  assign n21712 = n21704 & ~n21711 ;
  assign n21713 = ~n21693 & n21712 ;
  assign n21714 = ~n16687 & n21713 ;
  assign n21715 = ( n21430 & n21579 ) | ( n21430 & ~n21714 ) | ( n21579 & ~n21714 ) ;
  assign n21716 = ( n21430 & n21572 ) | ( n21430 & ~n21715 ) | ( n21572 & ~n21715 ) ;
  assign n21717 = ( n21430 & ~n21580 ) | ( n21430 & n21714 ) | ( ~n21580 & n21714 ) ;
  assign n21718 = ( n21572 & ~n21716 ) | ( n21572 & n21717 ) | ( ~n21716 & n21717 ) ;
  assign n21719 = n390 & ~n16161 ;
  assign n21720 = n3270 & ~n16150 ;
  assign n21721 = n3274 & ~n15954 ;
  assign n21722 = n3273 & ~n15806 ;
  assign n21723 = n21721 | n21722 ;
  assign n21724 = n21720 | n21723 ;
  assign n21725 = n21719 | n21724 ;
  assign n21726 = ( n21584 & n21718 ) | ( n21584 & n21725 ) | ( n21718 & n21725 ) ;
  assign n21727 = ( n21584 & ~n21718 ) | ( n21584 & n21725 ) | ( ~n21718 & n21725 ) ;
  assign n21728 = ( n21718 & ~n21726 ) | ( n21718 & n21727 ) | ( ~n21726 & n21727 ) ;
  assign n21729 = ( n21675 & n21685 ) | ( n21675 & ~n21728 ) | ( n21685 & ~n21728 ) ;
  assign n21730 = ( n21675 & ~n21685 ) | ( n21675 & n21728 ) | ( ~n21685 & n21728 ) ;
  assign n21731 = ( ~n21675 & n21729 ) | ( ~n21675 & n21730 ) | ( n21729 & n21730 ) ;
  assign n21732 = ( ~n21587 & n21665 ) | ( ~n21587 & n21731 ) | ( n21665 & n21731 ) ;
  assign n21733 = ( n21587 & n21665 ) | ( n21587 & ~n21731 ) | ( n21665 & ~n21731 ) ;
  assign n21734 = ( ~n21665 & n21732 ) | ( ~n21665 & n21733 ) | ( n21732 & n21733 ) ;
  assign n21735 = ( ~n21589 & n21655 ) | ( ~n21589 & n21734 ) | ( n21655 & n21734 ) ;
  assign n21736 = ( n21589 & n21655 ) | ( n21589 & ~n21734 ) | ( n21655 & ~n21734 ) ;
  assign n21737 = ( ~n21655 & n21735 ) | ( ~n21655 & n21736 ) | ( n21735 & n21736 ) ;
  assign n21738 = ( ~n21593 & n21645 ) | ( ~n21593 & n21737 ) | ( n21645 & n21737 ) ;
  assign n21739 = ( n21593 & n21645 ) | ( n21593 & ~n21737 ) | ( n21645 & ~n21737 ) ;
  assign n21740 = ( ~n21645 & n21738 ) | ( ~n21645 & n21739 ) | ( n21738 & n21739 ) ;
  assign n21741 = ( ~n21596 & n21635 ) | ( ~n21596 & n21740 ) | ( n21635 & n21740 ) ;
  assign n21742 = ( n21596 & n21635 ) | ( n21596 & ~n21740 ) | ( n21635 & ~n21740 ) ;
  assign n21743 = ( ~n21635 & n21741 ) | ( ~n21635 & n21742 ) | ( n21741 & n21742 ) ;
  assign n21744 = ( n21599 & n21625 ) | ( n21599 & ~n21743 ) | ( n21625 & ~n21743 ) ;
  assign n21745 = ( ~n21599 & n21625 ) | ( ~n21599 & n21743 ) | ( n21625 & n21743 ) ;
  assign n21746 = ( ~n21625 & n21744 ) | ( ~n21625 & n21745 ) | ( n21744 & n21745 ) ;
  assign n21747 = ( ~x8 & n21601 ) | ( ~x8 & n21746 ) | ( n21601 & n21746 ) ;
  assign n21748 = ( x8 & n21601 ) | ( x8 & ~n21746 ) | ( n21601 & ~n21746 ) ;
  assign n21749 = ( ~n21601 & n21747 ) | ( ~n21601 & n21748 ) | ( n21747 & n21748 ) ;
  assign n21750 = ( ~n21608 & n21611 ) | ( ~n21608 & n21749 ) | ( n21611 & n21749 ) ;
  assign n21751 = ( n21608 & n21611 ) | ( n21608 & ~n21749 ) | ( n21611 & ~n21749 ) ;
  assign n21752 = ( ~n21611 & n21750 ) | ( ~n21611 & n21751 ) | ( n21750 & n21751 ) ;
  assign n21753 = n21614 & ~n21752 ;
  assign n21754 = ~n21614 & n21752 ;
  assign n21755 = n21753 | n21754 ;
  assign n21756 = n6796 & ~n20095 ;
  assign n21757 = n6567 & n20091 ;
  assign n21758 = n21756 | n21757 ;
  assign n21759 = x11 & n21758 ;
  assign n21760 = n6571 & ~n20097 ;
  assign n21761 = ( ~x11 & n21758 ) | ( ~x11 & n21760 ) | ( n21758 & n21760 ) ;
  assign n21762 = x11 & ~n21760 ;
  assign n21763 = ( ~n21759 & n21761 ) | ( ~n21759 & n21762 ) | ( n21761 & n21762 ) ;
  assign n21764 = n6332 & n19882 ;
  assign n21765 = x14 & n21764 ;
  assign n21766 = n5909 & ~n19701 ;
  assign n21767 = n5914 | n21766 ;
  assign n21768 = ( n19916 & n21766 ) | ( n19916 & n21767 ) | ( n21766 & n21767 ) ;
  assign n21769 = n5915 | n21768 ;
  assign n21770 = ( n19920 & n21768 ) | ( n19920 & n21769 ) | ( n21768 & n21769 ) ;
  assign n21771 = x14 & ~n21770 ;
  assign n21772 = ( ~x14 & n21764 ) | ( ~x14 & n21770 ) | ( n21764 & n21770 ) ;
  assign n21773 = ( ~n21765 & n21771 ) | ( ~n21765 & n21772 ) | ( n21771 & n21772 ) ;
  assign n21774 = n5418 & ~n19374 ;
  assign n21775 = x17 & n21774 ;
  assign n21776 = n5413 & n19248 ;
  assign n21777 = n5417 | n21776 ;
  assign n21778 = ( n19368 & n21776 ) | ( n19368 & n21777 ) | ( n21776 & n21777 ) ;
  assign n21779 = n5584 & ~n19315 ;
  assign n21780 = n21778 | n21779 ;
  assign n21781 = x17 & ~n21780 ;
  assign n21782 = ( ~x17 & n21774 ) | ( ~x17 & n21780 ) | ( n21774 & n21780 ) ;
  assign n21783 = ( ~n21775 & n21781 ) | ( ~n21775 & n21782 ) | ( n21781 & n21782 ) ;
  assign n21784 = n4879 & ~n19182 ;
  assign n21785 = x20 & n21784 ;
  assign n21786 = n4874 & ~n18362 ;
  assign n21787 = n4878 | n21786 ;
  assign n21788 = ( n19177 & n21786 ) | ( n19177 & n21787 ) | ( n21786 & n21787 ) ;
  assign n21789 = n5232 & n18730 ;
  assign n21790 = n21788 | n21789 ;
  assign n21791 = x20 & ~n21790 ;
  assign n21792 = ( ~x20 & n21784 ) | ( ~x20 & n21790 ) | ( n21784 & n21790 ) ;
  assign n21793 = ( ~n21785 & n21791 ) | ( ~n21785 & n21792 ) | ( n21791 & n21792 ) ;
  assign n21794 = n4637 & ~n17963 ;
  assign n21795 = x23 & n21794 ;
  assign n21796 = n4584 & n17742 ;
  assign n21797 = n4649 | n21796 ;
  assign n21798 = ( ~n18258 & n21796 ) | ( ~n18258 & n21797 ) | ( n21796 & n21797 ) ;
  assign n21799 = n4591 | n21798 ;
  assign n21800 = ( n18268 & n21798 ) | ( n18268 & n21799 ) | ( n21798 & n21799 ) ;
  assign n21801 = x23 & ~n21800 ;
  assign n21802 = ( ~x23 & n21794 ) | ( ~x23 & n21800 ) | ( n21794 & n21800 ) ;
  assign n21803 = ( ~n21795 & n21801 ) | ( ~n21795 & n21802 ) | ( n21801 & n21802 ) ;
  assign n21804 = n3273 & ~n15954 ;
  assign n21805 = n3270 | n21804 ;
  assign n21806 = ( ~n16338 & n21804 ) | ( ~n16338 & n21805 ) | ( n21804 & n21805 ) ;
  assign n21807 = n390 | n21806 ;
  assign n21808 = ( ~n16349 & n21806 ) | ( ~n16349 & n21807 ) | ( n21806 & n21807 ) ;
  assign n21809 = n3274 & ~n16150 ;
  assign n21810 = n21808 | n21809 ;
  assign n21811 = n306 | n600 ;
  assign n21812 = n572 | n21811 ;
  assign n21813 = n957 | n2206 ;
  assign n21814 = n21812 | n21813 ;
  assign n21815 = n4945 | n21814 ;
  assign n21816 = n17284 | n17296 ;
  assign n21817 = n21815 | n21816 ;
  assign n21818 = n1134 | n1635 ;
  assign n21819 = n1991 | n21818 ;
  assign n21820 = n21817 | n21819 ;
  assign n21821 = n2498 | n21820 ;
  assign n21822 = n1079 | n21821 ;
  assign n21823 = n3048 & ~n21822 ;
  assign n21824 = ( x8 & n21572 ) | ( x8 & ~n21823 ) | ( n21572 & ~n21823 ) ;
  assign n21825 = ( x8 & ~n21572 ) | ( x8 & n21823 ) | ( ~n21572 & n21823 ) ;
  assign n21826 = ( ~x8 & n21824 ) | ( ~x8 & n21825 ) | ( n21824 & n21825 ) ;
  assign n21827 = ( n21716 & n21810 ) | ( n21716 & ~n21826 ) | ( n21810 & ~n21826 ) ;
  assign n21828 = ( ~n21716 & n21810 ) | ( ~n21716 & n21826 ) | ( n21810 & n21826 ) ;
  assign n21829 = ( ~n21810 & n21827 ) | ( ~n21810 & n21828 ) | ( n21827 & n21828 ) ;
  assign n21830 = n3541 & ~n16936 ;
  assign n21831 = x29 & n21830 ;
  assign n21832 = n3536 & ~n16531 ;
  assign n21833 = n4039 | n21832 ;
  assign n21834 = ( n16925 & n21832 ) | ( n16925 & n21833 ) | ( n21832 & n21833 ) ;
  assign n21835 = n3501 & n16724 ;
  assign n21836 = n21834 | n21835 ;
  assign n21837 = x29 & ~n21836 ;
  assign n21838 = ( ~x29 & n21830 ) | ( ~x29 & n21836 ) | ( n21830 & n21836 ) ;
  assign n21839 = ( ~n21831 & n21837 ) | ( ~n21831 & n21838 ) | ( n21837 & n21838 ) ;
  assign n21840 = ( n21727 & ~n21829 ) | ( n21727 & n21839 ) | ( ~n21829 & n21839 ) ;
  assign n21841 = ( n21727 & n21829 ) | ( n21727 & ~n21839 ) | ( n21829 & ~n21839 ) ;
  assign n21842 = ( ~n21727 & n21840 ) | ( ~n21727 & n21841 ) | ( n21840 & n21841 ) ;
  assign n21843 = n4215 & ~n17635 ;
  assign n21844 = n4200 & n17346 ;
  assign n21845 = n2083 & ~n17126 ;
  assign n21846 = n21844 | n21845 ;
  assign n21847 = n21843 | n21846 ;
  assign n21848 = x26 & n21847 ;
  assign n21849 = n4203 & ~n17646 ;
  assign n21850 = ( ~x26 & n21847 ) | ( ~x26 & n21849 ) | ( n21847 & n21849 ) ;
  assign n21851 = x26 & ~n21849 ;
  assign n21852 = ( ~n21848 & n21850 ) | ( ~n21848 & n21851 ) | ( n21850 & n21851 ) ;
  assign n21853 = ( n21729 & n21842 ) | ( n21729 & ~n21852 ) | ( n21842 & ~n21852 ) ;
  assign n21854 = ( n21729 & ~n21842 ) | ( n21729 & n21852 ) | ( ~n21842 & n21852 ) ;
  assign n21855 = ( ~n21729 & n21853 ) | ( ~n21729 & n21854 ) | ( n21853 & n21854 ) ;
  assign n21856 = ( n21733 & n21803 ) | ( n21733 & ~n21855 ) | ( n21803 & ~n21855 ) ;
  assign n21857 = ( n21733 & ~n21803 ) | ( n21733 & n21855 ) | ( ~n21803 & n21855 ) ;
  assign n21858 = ( ~n21733 & n21856 ) | ( ~n21733 & n21857 ) | ( n21856 & n21857 ) ;
  assign n21859 = ( n21736 & n21793 ) | ( n21736 & ~n21858 ) | ( n21793 & ~n21858 ) ;
  assign n21860 = ( n21736 & ~n21793 ) | ( n21736 & n21858 ) | ( ~n21793 & n21858 ) ;
  assign n21861 = ( ~n21736 & n21859 ) | ( ~n21736 & n21860 ) | ( n21859 & n21860 ) ;
  assign n21862 = ( n21739 & n21783 ) | ( n21739 & ~n21861 ) | ( n21783 & ~n21861 ) ;
  assign n21863 = ( ~n21739 & n21783 ) | ( ~n21739 & n21861 ) | ( n21783 & n21861 ) ;
  assign n21864 = ( ~n21783 & n21862 ) | ( ~n21783 & n21863 ) | ( n21862 & n21863 ) ;
  assign n21865 = ( n21742 & n21773 ) | ( n21742 & ~n21864 ) | ( n21773 & ~n21864 ) ;
  assign n21866 = ( ~n21742 & n21773 ) | ( ~n21742 & n21864 ) | ( n21773 & n21864 ) ;
  assign n21867 = ( ~n21773 & n21865 ) | ( ~n21773 & n21866 ) | ( n21865 & n21866 ) ;
  assign n21868 = ( n21744 & ~n21763 ) | ( n21744 & n21867 ) | ( ~n21763 & n21867 ) ;
  assign n21869 = ( n21744 & n21763 ) | ( n21744 & ~n21867 ) | ( n21763 & ~n21867 ) ;
  assign n21870 = ( ~n21744 & n21868 ) | ( ~n21744 & n21869 ) | ( n21868 & n21869 ) ;
  assign n21871 = ( n21748 & n21751 ) | ( n21748 & ~n21870 ) | ( n21751 & ~n21870 ) ;
  assign n21872 = ( ~n21748 & n21751 ) | ( ~n21748 & n21870 ) | ( n21751 & n21870 ) ;
  assign n21873 = ( ~n21751 & n21871 ) | ( ~n21751 & n21872 ) | ( n21871 & n21872 ) ;
  assign n21874 = n21753 & ~n21873 ;
  assign n21875 = ~n21753 & n21873 ;
  assign n21876 = n21874 | n21875 ;
  assign n21877 = n5584 & n19368 ;
  assign n21878 = x17 & n21877 ;
  assign n21879 = n5413 & ~n19315 ;
  assign n21880 = n5417 | n21879 ;
  assign n21881 = ( ~n19701 & n21879 ) | ( ~n19701 & n21880 ) | ( n21879 & n21880 ) ;
  assign n21882 = n5418 | n21881 ;
  assign n21883 = ( ~n19706 & n21881 ) | ( ~n19706 & n21882 ) | ( n21881 & n21882 ) ;
  assign n21884 = x17 & ~n21883 ;
  assign n21885 = ( ~x17 & n21877 ) | ( ~x17 & n21883 ) | ( n21877 & n21883 ) ;
  assign n21886 = ( ~n21878 & n21884 ) | ( ~n21878 & n21885 ) | ( n21884 & n21885 ) ;
  assign n21887 = n5232 & n19177 ;
  assign n21888 = x20 & n21887 ;
  assign n21889 = n4874 & n18730 ;
  assign n21890 = n4878 | n21889 ;
  assign n21891 = ( n19248 & n21889 ) | ( n19248 & n21890 ) | ( n21889 & n21890 ) ;
  assign n21892 = n4879 | n21891 ;
  assign n21893 = ( n19253 & n21891 ) | ( n19253 & n21892 ) | ( n21891 & n21892 ) ;
  assign n21894 = x20 & ~n21893 ;
  assign n21895 = ( ~x20 & n21887 ) | ( ~x20 & n21893 ) | ( n21887 & n21893 ) ;
  assign n21896 = ( ~n21888 & n21894 ) | ( ~n21888 & n21895 ) | ( n21894 & n21895 ) ;
  assign n21897 = n4637 & ~n18258 ;
  assign n21898 = x23 & n21897 ;
  assign n21899 = n4584 & ~n17963 ;
  assign n21900 = n4649 | n21899 ;
  assign n21901 = ( ~n18362 & n21899 ) | ( ~n18362 & n21900 ) | ( n21899 & n21900 ) ;
  assign n21902 = n4591 | n21901 ;
  assign n21903 = ( ~n18373 & n21901 ) | ( ~n18373 & n21902 ) | ( n21901 & n21902 ) ;
  assign n21904 = x23 & ~n21903 ;
  assign n21905 = ( ~x23 & n21897 ) | ( ~x23 & n21903 ) | ( n21897 & n21903 ) ;
  assign n21906 = ( ~n21898 & n21904 ) | ( ~n21898 & n21905 ) | ( n21904 & n21905 ) ;
  assign n21907 = n4215 & n17742 ;
  assign n21908 = x26 & n21907 ;
  assign n21909 = n4200 & ~n17635 ;
  assign n21910 = n2083 & n17346 ;
  assign n21911 = n21909 | n21910 ;
  assign n21912 = n4203 | n21911 ;
  assign n21913 = ( ~n17749 & n21911 ) | ( ~n17749 & n21912 ) | ( n21911 & n21912 ) ;
  assign n21914 = x26 & ~n21913 ;
  assign n21915 = ( ~x26 & n21907 ) | ( ~x26 & n21913 ) | ( n21907 & n21913 ) ;
  assign n21916 = ( ~n21908 & n21914 ) | ( ~n21908 & n21915 ) | ( n21914 & n21915 ) ;
  assign n21917 = n3501 & n16925 ;
  assign n21918 = x29 & n21917 ;
  assign n21919 = n3536 & n16724 ;
  assign n21920 = n4039 | n21919 ;
  assign n21921 = ( ~n17126 & n21919 ) | ( ~n17126 & n21920 ) | ( n21919 & n21920 ) ;
  assign n21922 = n3541 | n21921 ;
  assign n21923 = ( ~n17139 & n21921 ) | ( ~n17139 & n21922 ) | ( n21921 & n21922 ) ;
  assign n21924 = x29 & ~n21923 ;
  assign n21925 = ( ~x29 & n21917 ) | ( ~x29 & n21923 ) | ( n21917 & n21923 ) ;
  assign n21926 = ( ~n21918 & n21924 ) | ( ~n21918 & n21925 ) | ( n21924 & n21925 ) ;
  assign n21927 = n298 | n1606 ;
  assign n21928 = n1935 | n21927 ;
  assign n21929 = n285 | n308 ;
  assign n21930 = n2964 | n21929 ;
  assign n21931 = n21928 | n21930 ;
  assign n21932 = n16491 | n21931 ;
  assign n21933 = n80 | n147 ;
  assign n21934 = n21932 | n21933 ;
  assign n21935 = n922 | n1678 ;
  assign n21936 = n2097 | n2979 ;
  assign n21937 = n21935 | n21936 ;
  assign n21938 = n4777 | n21937 ;
  assign n21939 = n21934 | n21938 ;
  assign n21940 = n857 | n21939 ;
  assign n21941 = n2230 & ~n21940 ;
  assign n21942 = n3273 & ~n16150 ;
  assign n21943 = n3270 | n21942 ;
  assign n21944 = ( ~n16531 & n21942 ) | ( ~n16531 & n21943 ) | ( n21942 & n21943 ) ;
  assign n21945 = n390 | n21944 ;
  assign n21946 = ( ~n16542 & n21944 ) | ( ~n16542 & n21945 ) | ( n21944 & n21945 ) ;
  assign n21947 = n3274 & ~n16338 ;
  assign n21948 = n21946 | n21947 ;
  assign n21949 = ( n21825 & n21941 ) | ( n21825 & ~n21948 ) | ( n21941 & ~n21948 ) ;
  assign n21950 = ( ~n21825 & n21941 ) | ( ~n21825 & n21948 ) | ( n21941 & n21948 ) ;
  assign n21951 = ( ~n21941 & n21949 ) | ( ~n21941 & n21950 ) | ( n21949 & n21950 ) ;
  assign n21952 = ( ~n21828 & n21926 ) | ( ~n21828 & n21951 ) | ( n21926 & n21951 ) ;
  assign n21953 = ( n21828 & n21926 ) | ( n21828 & ~n21951 ) | ( n21926 & ~n21951 ) ;
  assign n21954 = ( ~n21926 & n21952 ) | ( ~n21926 & n21953 ) | ( n21952 & n21953 ) ;
  assign n21955 = ( n21840 & n21916 ) | ( n21840 & ~n21954 ) | ( n21916 & ~n21954 ) ;
  assign n21956 = ( ~n21840 & n21916 ) | ( ~n21840 & n21954 ) | ( n21916 & n21954 ) ;
  assign n21957 = ( ~n21916 & n21955 ) | ( ~n21916 & n21956 ) | ( n21955 & n21956 ) ;
  assign n21958 = ( n21854 & n21906 ) | ( n21854 & ~n21957 ) | ( n21906 & ~n21957 ) ;
  assign n21959 = ( ~n21854 & n21906 ) | ( ~n21854 & n21957 ) | ( n21906 & n21957 ) ;
  assign n21960 = ( ~n21906 & n21958 ) | ( ~n21906 & n21959 ) | ( n21958 & n21959 ) ;
  assign n21961 = ( n21856 & n21896 ) | ( n21856 & ~n21960 ) | ( n21896 & ~n21960 ) ;
  assign n21962 = ( ~n21856 & n21896 ) | ( ~n21856 & n21960 ) | ( n21896 & n21960 ) ;
  assign n21963 = ( ~n21896 & n21961 ) | ( ~n21896 & n21962 ) | ( n21961 & n21962 ) ;
  assign n21964 = ( n21859 & n21886 ) | ( n21859 & ~n21963 ) | ( n21886 & ~n21963 ) ;
  assign n21965 = ( ~n21859 & n21886 ) | ( ~n21859 & n21963 ) | ( n21886 & n21963 ) ;
  assign n21966 = ( ~n21886 & n21964 ) | ( ~n21886 & n21965 ) | ( n21964 & n21965 ) ;
  assign n21967 = n5914 & n20091 ;
  assign n21968 = n5915 | n21967 ;
  assign n21969 = ( n20101 & n21967 ) | ( n20101 & n21968 ) | ( n21967 & n21968 ) ;
  assign n21970 = n6332 & n19916 ;
  assign n21971 = n21969 | n21970 ;
  assign n21972 = n5908 & n19882 ;
  assign n21973 = n5909 & n19882 ;
  assign n21974 = x14 & ~n21973 ;
  assign n21975 = ( ~n21971 & n21972 ) | ( ~n21971 & n21974 ) | ( n21972 & n21974 ) ;
  assign n21976 = n21971 | n21974 ;
  assign n21977 = ( ~x14 & n21975 ) | ( ~x14 & n21976 ) | ( n21975 & n21976 ) ;
  assign n21978 = ( n21862 & n21966 ) | ( n21862 & n21977 ) | ( n21966 & n21977 ) ;
  assign n21979 = ( n21862 & ~n21966 ) | ( n21862 & n21977 ) | ( ~n21966 & n21977 ) ;
  assign n21980 = ( n21966 & ~n21978 ) | ( n21966 & n21979 ) | ( ~n21978 & n21979 ) ;
  assign n21981 = n6565 & ~n20095 ;
  assign n21982 = n6563 | n20095 ;
  assign n21983 = ( x11 & n21981 ) | ( x11 & n21982 ) | ( n21981 & n21982 ) ;
  assign n21984 = ( n21865 & ~n21980 ) | ( n21865 & n21983 ) | ( ~n21980 & n21983 ) ;
  assign n21985 = ( n21865 & n21980 ) | ( n21865 & n21983 ) | ( n21980 & n21983 ) ;
  assign n21986 = ( n21980 & n21984 ) | ( n21980 & ~n21985 ) | ( n21984 & ~n21985 ) ;
  assign n21987 = ( n21869 & n21871 ) | ( n21869 & ~n21986 ) | ( n21871 & ~n21986 ) ;
  assign n21988 = ( ~n21869 & n21871 ) | ( ~n21869 & n21986 ) | ( n21871 & n21986 ) ;
  assign n21989 = ( ~n21871 & n21987 ) | ( ~n21871 & n21988 ) | ( n21987 & n21988 ) ;
  assign n21990 = n21874 & ~n21989 ;
  assign n21991 = ~n21874 & n21989 ;
  assign n21992 = n21990 | n21991 ;
  assign n21993 = n5909 & n19916 ;
  assign n21994 = n5914 | n21993 ;
  assign n21995 = ( ~n20095 & n21993 ) | ( ~n20095 & n21994 ) | ( n21993 & n21994 ) ;
  assign n21996 = n6332 & n20091 ;
  assign n21997 = n21995 | n21996 ;
  assign n21998 = x14 & n21997 ;
  assign n21999 = n5915 & ~n20100 ;
  assign n22000 = ( ~x14 & n21997 ) | ( ~x14 & n21999 ) | ( n21997 & n21999 ) ;
  assign n22001 = x14 & ~n21999 ;
  assign n22002 = ( ~n21998 & n22000 ) | ( ~n21998 & n22001 ) | ( n22000 & n22001 ) ;
  assign n22003 = n5584 & ~n19701 ;
  assign n22004 = x17 & n22003 ;
  assign n22005 = n5413 & n19368 ;
  assign n22006 = n5417 | n22005 ;
  assign n22007 = ( n19882 & n22005 ) | ( n19882 & n22006 ) | ( n22005 & n22006 ) ;
  assign n22008 = n5418 | n22007 ;
  assign n22009 = ( ~n19893 & n22007 ) | ( ~n19893 & n22008 ) | ( n22007 & n22008 ) ;
  assign n22010 = x17 & ~n22009 ;
  assign n22011 = ( ~x17 & n22003 ) | ( ~x17 & n22009 ) | ( n22003 & n22009 ) ;
  assign n22012 = ( ~n22004 & n22010 ) | ( ~n22004 & n22011 ) | ( n22010 & n22011 ) ;
  assign n22013 = n5232 & n19248 ;
  assign n22014 = x20 & n22013 ;
  assign n22015 = n4874 & n19177 ;
  assign n22016 = n4878 | n22015 ;
  assign n22017 = ( ~n19315 & n22015 ) | ( ~n19315 & n22016 ) | ( n22015 & n22016 ) ;
  assign n22018 = n4879 | n22017 ;
  assign n22019 = ( ~n19320 & n22017 ) | ( ~n19320 & n22018 ) | ( n22017 & n22018 ) ;
  assign n22020 = x20 & ~n22019 ;
  assign n22021 = ( ~x20 & n22013 ) | ( ~x20 & n22019 ) | ( n22013 & n22019 ) ;
  assign n22022 = ( ~n22014 & n22020 ) | ( ~n22014 & n22021 ) | ( n22020 & n22021 ) ;
  assign n22023 = n4649 & n18730 ;
  assign n22024 = n4591 | n22023 ;
  assign n22025 = ( n18735 & n22023 ) | ( n18735 & n22024 ) | ( n22023 & n22024 ) ;
  assign n22026 = n4637 & ~n18362 ;
  assign n22027 = n22025 | n22026 ;
  assign n22028 = n4583 & ~n18258 ;
  assign n22029 = n4584 & ~n18258 ;
  assign n22030 = x23 & ~n22029 ;
  assign n22031 = ( ~n22027 & n22028 ) | ( ~n22027 & n22030 ) | ( n22028 & n22030 ) ;
  assign n22032 = n22027 | n22030 ;
  assign n22033 = ( ~x23 & n22031 ) | ( ~x23 & n22032 ) | ( n22031 & n22032 ) ;
  assign n22034 = n4215 & ~n17963 ;
  assign n22035 = n4200 & n17742 ;
  assign n22036 = n2083 & ~n17635 ;
  assign n22037 = n22035 | n22036 ;
  assign n22038 = n22034 | n22037 ;
  assign n22039 = x26 & n22038 ;
  assign n22040 = n4203 & ~n17976 ;
  assign n22041 = ( ~x26 & n22038 ) | ( ~x26 & n22040 ) | ( n22038 & n22040 ) ;
  assign n22042 = x26 & ~n22040 ;
  assign n22043 = ( ~n22039 & n22041 ) | ( ~n22039 & n22042 ) | ( n22041 & n22042 ) ;
  assign n22044 = n3501 & ~n17126 ;
  assign n22045 = x29 & n22044 ;
  assign n22046 = n3536 & n16925 ;
  assign n22047 = n4039 | n22046 ;
  assign n22048 = ( n17346 & n22046 ) | ( n17346 & n22047 ) | ( n22046 & n22047 ) ;
  assign n22049 = n3541 | n22048 ;
  assign n22050 = ( ~n17356 & n22048 ) | ( ~n17356 & n22049 ) | ( n22048 & n22049 ) ;
  assign n22051 = x29 & ~n22050 ;
  assign n22052 = ( ~x29 & n22044 ) | ( ~x29 & n22050 ) | ( n22044 & n22050 ) ;
  assign n22053 = ( ~n22045 & n22051 ) | ( ~n22045 & n22052 ) | ( n22051 & n22052 ) ;
  assign n22054 = n3273 & ~n16338 ;
  assign n22055 = n3270 | n22054 ;
  assign n22056 = ( n16724 & n22054 ) | ( n16724 & n22055 ) | ( n22054 & n22055 ) ;
  assign n22057 = n390 | n22056 ;
  assign n22058 = ( n16735 & n22056 ) | ( n16735 & n22057 ) | ( n22056 & n22057 ) ;
  assign n22059 = n3274 & ~n16531 ;
  assign n22060 = n22058 | n22059 ;
  assign n22061 = n917 | n1601 ;
  assign n22062 = n1518 | n22061 ;
  assign n22063 = n13914 | n22062 ;
  assign n22064 = n271 | n3154 ;
  assign n22065 = n891 | n22064 ;
  assign n22066 = n22063 | n22065 ;
  assign n22067 = n1876 | n1939 ;
  assign n22068 = n304 | n22067 ;
  assign n22069 = n987 | n1360 ;
  assign n22070 = n2995 | n22069 ;
  assign n22071 = n22068 | n22070 ;
  assign n22072 = n17309 | n22071 ;
  assign n22073 = n22066 | n22072 ;
  assign n22074 = n5126 | n22073 ;
  assign n22075 = n21571 | n22074 ;
  assign n22076 = ( n21941 & n21950 ) | ( n21941 & n22075 ) | ( n21950 & n22075 ) ;
  assign n22077 = ( ~n21941 & n21950 ) | ( ~n21941 & n22075 ) | ( n21950 & n22075 ) ;
  assign n22078 = ( n21941 & ~n22076 ) | ( n21941 & n22077 ) | ( ~n22076 & n22077 ) ;
  assign n22079 = ( ~n22053 & n22060 ) | ( ~n22053 & n22078 ) | ( n22060 & n22078 ) ;
  assign n22080 = ( n22053 & n22060 ) | ( n22053 & n22078 ) | ( n22060 & n22078 ) ;
  assign n22081 = ( n22053 & n22079 ) | ( n22053 & ~n22080 ) | ( n22079 & ~n22080 ) ;
  assign n22082 = ( ~n21953 & n22043 ) | ( ~n21953 & n22081 ) | ( n22043 & n22081 ) ;
  assign n22083 = ( n21953 & n22043 ) | ( n21953 & n22081 ) | ( n22043 & n22081 ) ;
  assign n22084 = ( n21953 & n22082 ) | ( n21953 & ~n22083 ) | ( n22082 & ~n22083 ) ;
  assign n22085 = ( n21955 & n22033 ) | ( n21955 & n22084 ) | ( n22033 & n22084 ) ;
  assign n22086 = ( n21955 & ~n22033 ) | ( n21955 & n22084 ) | ( ~n22033 & n22084 ) ;
  assign n22087 = ( n22033 & ~n22085 ) | ( n22033 & n22086 ) | ( ~n22085 & n22086 ) ;
  assign n22088 = ( ~n21958 & n22022 ) | ( ~n21958 & n22087 ) | ( n22022 & n22087 ) ;
  assign n22089 = ( n21958 & n22022 ) | ( n21958 & n22087 ) | ( n22022 & n22087 ) ;
  assign n22090 = ( n21958 & n22088 ) | ( n21958 & ~n22089 ) | ( n22088 & ~n22089 ) ;
  assign n22091 = ( n21961 & n22012 ) | ( n21961 & n22090 ) | ( n22012 & n22090 ) ;
  assign n22092 = ( n21961 & ~n22012 ) | ( n21961 & n22090 ) | ( ~n22012 & n22090 ) ;
  assign n22093 = ( n22012 & ~n22091 ) | ( n22012 & n22092 ) | ( ~n22091 & n22092 ) ;
  assign n22094 = ( n21964 & ~n22002 ) | ( n21964 & n22093 ) | ( ~n22002 & n22093 ) ;
  assign n22095 = ( n21964 & n22002 ) | ( n21964 & n22093 ) | ( n22002 & n22093 ) ;
  assign n22096 = ( n22002 & n22094 ) | ( n22002 & ~n22095 ) | ( n22094 & ~n22095 ) ;
  assign n22097 = ( ~x11 & n21979 ) | ( ~x11 & n22096 ) | ( n21979 & n22096 ) ;
  assign n22098 = ( x11 & n21979 ) | ( x11 & n22096 ) | ( n21979 & n22096 ) ;
  assign n22099 = ( x11 & n22097 ) | ( x11 & ~n22098 ) | ( n22097 & ~n22098 ) ;
  assign n22100 = ( n21984 & ~n21987 ) | ( n21984 & n22099 ) | ( ~n21987 & n22099 ) ;
  assign n22101 = ( n21984 & n21987 ) | ( n21984 & n22099 ) | ( n21987 & n22099 ) ;
  assign n22102 = ( n21987 & n22100 ) | ( n21987 & ~n22101 ) | ( n22100 & ~n22101 ) ;
  assign n22103 = n21990 & ~n22102 ;
  assign n22104 = n21990 & n22102 ;
  assign n22105 = ( n22102 & n22103 ) | ( n22102 & ~n22104 ) | ( n22103 & ~n22104 ) ;
  assign n22106 = n6332 & ~n20095 ;
  assign n22107 = n5909 & n20091 ;
  assign n22108 = n22106 | n22107 ;
  assign n22109 = x14 & n22108 ;
  assign n22110 = n5915 & ~n20097 ;
  assign n22111 = ( ~x14 & n22108 ) | ( ~x14 & n22110 ) | ( n22108 & n22110 ) ;
  assign n22112 = x14 & ~n22110 ;
  assign n22113 = ( ~n22109 & n22111 ) | ( ~n22109 & n22112 ) | ( n22111 & n22112 ) ;
  assign n22114 = n5418 & n19920 ;
  assign n22115 = x17 & n22114 ;
  assign n22116 = n5413 & ~n19701 ;
  assign n22117 = n5417 | n22116 ;
  assign n22118 = ( n19916 & n22116 ) | ( n19916 & n22117 ) | ( n22116 & n22117 ) ;
  assign n22119 = n5584 & n19882 ;
  assign n22120 = n22118 | n22119 ;
  assign n22121 = x17 & ~n22120 ;
  assign n22122 = ( ~x17 & n22114 ) | ( ~x17 & n22120 ) | ( n22114 & n22120 ) ;
  assign n22123 = ( ~n22115 & n22121 ) | ( ~n22115 & n22122 ) | ( n22121 & n22122 ) ;
  assign n22124 = n4879 & ~n19374 ;
  assign n22125 = x20 & n22124 ;
  assign n22126 = n4874 & n19248 ;
  assign n22127 = n4878 | n22126 ;
  assign n22128 = ( n19368 & n22126 ) | ( n19368 & n22127 ) | ( n22126 & n22127 ) ;
  assign n22129 = n5232 & ~n19315 ;
  assign n22130 = n22128 | n22129 ;
  assign n22131 = x20 & ~n22130 ;
  assign n22132 = ( ~x20 & n22124 ) | ( ~x20 & n22130 ) | ( n22124 & n22130 ) ;
  assign n22133 = ( ~n22125 & n22131 ) | ( ~n22125 & n22132 ) | ( n22131 & n22132 ) ;
  assign n22134 = n4637 & n18730 ;
  assign n22135 = x23 & n22134 ;
  assign n22136 = n4584 & ~n18362 ;
  assign n22137 = n4649 | n22136 ;
  assign n22138 = ( n19177 & n22136 ) | ( n19177 & n22137 ) | ( n22136 & n22137 ) ;
  assign n22139 = n4591 | n22138 ;
  assign n22140 = ( ~n19182 & n22138 ) | ( ~n19182 & n22139 ) | ( n22138 & n22139 ) ;
  assign n22141 = x23 & ~n22140 ;
  assign n22142 = ( ~x23 & n22134 ) | ( ~x23 & n22140 ) | ( n22134 & n22140 ) ;
  assign n22143 = ( ~n22135 & n22141 ) | ( ~n22135 & n22142 ) | ( n22141 & n22142 ) ;
  assign n22144 = n4215 & ~n18258 ;
  assign n22145 = n4200 & ~n17963 ;
  assign n22146 = n2083 & n17742 ;
  assign n22147 = n22145 | n22146 ;
  assign n22148 = n22144 | n22147 ;
  assign n22149 = x26 & n22148 ;
  assign n22150 = n4203 & n18268 ;
  assign n22151 = ( ~x26 & n22148 ) | ( ~x26 & n22150 ) | ( n22148 & n22150 ) ;
  assign n22152 = x26 & ~n22150 ;
  assign n22153 = ( ~n22149 & n22151 ) | ( ~n22149 & n22152 ) | ( n22151 & n22152 ) ;
  assign n22154 = n3501 & n17346 ;
  assign n22155 = x29 & n22154 ;
  assign n22156 = n3536 & ~n17126 ;
  assign n22157 = n4039 | n22156 ;
  assign n22158 = ( ~n17635 & n22156 ) | ( ~n17635 & n22157 ) | ( n22156 & n22157 ) ;
  assign n22159 = n3541 | n22158 ;
  assign n22160 = ( ~n17646 & n22158 ) | ( ~n17646 & n22159 ) | ( n22158 & n22159 ) ;
  assign n22161 = x29 & ~n22160 ;
  assign n22162 = ( ~x29 & n22154 ) | ( ~x29 & n22160 ) | ( n22154 & n22160 ) ;
  assign n22163 = ( ~n22155 & n22161 ) | ( ~n22155 & n22162 ) | ( n22161 & n22162 ) ;
  assign n22164 = n3273 & ~n16531 ;
  assign n22165 = n3270 | n22164 ;
  assign n22166 = ( n16925 & n22164 ) | ( n16925 & n22165 ) | ( n22164 & n22165 ) ;
  assign n22167 = n390 | n22166 ;
  assign n22168 = ( ~n16936 & n22166 ) | ( ~n16936 & n22167 ) | ( n22166 & n22167 ) ;
  assign n22169 = n3274 & n16724 ;
  assign n22170 = n22168 | n22169 ;
  assign n22171 = n269 | n287 ;
  assign n22172 = n257 | n22171 ;
  assign n22173 = n123 | n22172 ;
  assign n22174 = n1364 | n1843 ;
  assign n22175 = n22173 | n22174 ;
  assign n22176 = n1138 | n4889 ;
  assign n22177 = n22175 | n22176 ;
  assign n22178 = n956 | n3448 ;
  assign n22179 = n2629 | n22178 ;
  assign n22180 = n22177 | n22179 ;
  assign n22181 = n2616 | n4931 ;
  assign n22182 = n1973 | n22181 ;
  assign n22183 = n22180 | n22182 ;
  assign n22184 = n2039 & ~n22183 ;
  assign n22185 = ~n898 & n22184 ;
  assign n22186 = ( ~x11 & n21941 ) | ( ~x11 & n22185 ) | ( n21941 & n22185 ) ;
  assign n22187 = ( x11 & n21941 ) | ( x11 & n22185 ) | ( n21941 & n22185 ) ;
  assign n22188 = ( x11 & n22186 ) | ( x11 & ~n22187 ) | ( n22186 & ~n22187 ) ;
  assign n22189 = ( n22076 & n22170 ) | ( n22076 & ~n22188 ) | ( n22170 & ~n22188 ) ;
  assign n22190 = ( n22076 & ~n22170 ) | ( n22076 & n22188 ) | ( ~n22170 & n22188 ) ;
  assign n22191 = ( ~n22076 & n22189 ) | ( ~n22076 & n22190 ) | ( n22189 & n22190 ) ;
  assign n22192 = ( n22080 & n22163 ) | ( n22080 & ~n22191 ) | ( n22163 & ~n22191 ) ;
  assign n22193 = ( n22080 & ~n22163 ) | ( n22080 & n22191 ) | ( ~n22163 & n22191 ) ;
  assign n22194 = ( ~n22080 & n22192 ) | ( ~n22080 & n22193 ) | ( n22192 & n22193 ) ;
  assign n22195 = ( n22083 & n22153 ) | ( n22083 & ~n22194 ) | ( n22153 & ~n22194 ) ;
  assign n22196 = ( ~n22083 & n22153 ) | ( ~n22083 & n22194 ) | ( n22153 & n22194 ) ;
  assign n22197 = ( ~n22153 & n22195 ) | ( ~n22153 & n22196 ) | ( n22195 & n22196 ) ;
  assign n22198 = ( n22085 & n22143 ) | ( n22085 & ~n22197 ) | ( n22143 & ~n22197 ) ;
  assign n22199 = ( n22085 & ~n22143 ) | ( n22085 & n22197 ) | ( ~n22143 & n22197 ) ;
  assign n22200 = ( ~n22085 & n22198 ) | ( ~n22085 & n22199 ) | ( n22198 & n22199 ) ;
  assign n22201 = ( ~n22089 & n22133 ) | ( ~n22089 & n22200 ) | ( n22133 & n22200 ) ;
  assign n22202 = ( n22089 & n22133 ) | ( n22089 & ~n22200 ) | ( n22133 & ~n22200 ) ;
  assign n22203 = ( ~n22133 & n22201 ) | ( ~n22133 & n22202 ) | ( n22201 & n22202 ) ;
  assign n22204 = ( n22091 & ~n22123 ) | ( n22091 & n22203 ) | ( ~n22123 & n22203 ) ;
  assign n22205 = ( n22091 & n22123 ) | ( n22091 & ~n22203 ) | ( n22123 & ~n22203 ) ;
  assign n22206 = ( ~n22091 & n22204 ) | ( ~n22091 & n22205 ) | ( n22204 & n22205 ) ;
  assign n22207 = ( n22095 & n22113 ) | ( n22095 & ~n22206 ) | ( n22113 & ~n22206 ) ;
  assign n22208 = ( n22095 & ~n22113 ) | ( n22095 & n22206 ) | ( ~n22113 & n22206 ) ;
  assign n22209 = ( ~n22095 & n22207 ) | ( ~n22095 & n22208 ) | ( n22207 & n22208 ) ;
  assign n22210 = ( ~n22098 & n22101 ) | ( ~n22098 & n22209 ) | ( n22101 & n22209 ) ;
  assign n22211 = ( n22098 & n22101 ) | ( n22098 & ~n22209 ) | ( n22101 & ~n22209 ) ;
  assign n22212 = ( ~n22101 & n22210 ) | ( ~n22101 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22213 = n22104 & ~n22212 ;
  assign n22214 = ~n22104 & n22212 ;
  assign n22215 = n22213 | n22214 ;
  assign n22216 = n5584 & n19916 ;
  assign n22217 = x17 & n22216 ;
  assign n22218 = n5413 & n19882 ;
  assign n22219 = n5417 | n22218 ;
  assign n22220 = ( n20091 & n22218 ) | ( n20091 & n22219 ) | ( n22218 & n22219 ) ;
  assign n22221 = n5418 | n22220 ;
  assign n22222 = ( n20101 & n22220 ) | ( n20101 & n22221 ) | ( n22220 & n22221 ) ;
  assign n22223 = x17 & ~n22222 ;
  assign n22224 = ( ~x17 & n22216 ) | ( ~x17 & n22222 ) | ( n22216 & n22222 ) ;
  assign n22225 = ( ~n22217 & n22223 ) | ( ~n22217 & n22224 ) | ( n22223 & n22224 ) ;
  assign n22226 = n4874 & ~n19315 ;
  assign n22227 = n4878 | n22226 ;
  assign n22228 = ( ~n19701 & n22226 ) | ( ~n19701 & n22227 ) | ( n22226 & n22227 ) ;
  assign n22229 = n5232 & n19368 ;
  assign n22230 = n22228 | n22229 ;
  assign n22231 = x20 & n22230 ;
  assign n22232 = n4879 & ~n19706 ;
  assign n22233 = x20 & ~n22232 ;
  assign n22234 = ( ~x20 & n22230 ) | ( ~x20 & n22232 ) | ( n22230 & n22232 ) ;
  assign n22235 = ( ~n22231 & n22233 ) | ( ~n22231 & n22234 ) | ( n22233 & n22234 ) ;
  assign n22236 = n4637 & n19177 ;
  assign n22237 = x23 & n22236 ;
  assign n22238 = n4584 & n18730 ;
  assign n22239 = n4649 | n22238 ;
  assign n22240 = ( n19248 & n22238 ) | ( n19248 & n22239 ) | ( n22238 & n22239 ) ;
  assign n22241 = n4591 | n22240 ;
  assign n22242 = ( n19253 & n22240 ) | ( n19253 & n22241 ) | ( n22240 & n22241 ) ;
  assign n22243 = x23 & ~n22242 ;
  assign n22244 = ( ~x23 & n22236 ) | ( ~x23 & n22242 ) | ( n22236 & n22242 ) ;
  assign n22245 = ( ~n22237 & n22243 ) | ( ~n22237 & n22244 ) | ( n22243 & n22244 ) ;
  assign n22246 = n4215 & ~n18362 ;
  assign n22247 = n4200 & ~n18258 ;
  assign n22248 = n2083 & ~n17963 ;
  assign n22249 = n22247 | n22248 ;
  assign n22250 = n22246 | n22249 ;
  assign n22251 = x26 & n22250 ;
  assign n22252 = n4203 & ~n18373 ;
  assign n22253 = ( ~x26 & n22250 ) | ( ~x26 & n22252 ) | ( n22250 & n22252 ) ;
  assign n22254 = x26 & ~n22252 ;
  assign n22255 = ( ~n22251 & n22253 ) | ( ~n22251 & n22254 ) | ( n22253 & n22254 ) ;
  assign n22256 = n3541 & ~n17749 ;
  assign n22257 = x29 & n22256 ;
  assign n22258 = n4039 & n17742 ;
  assign n22259 = n3501 & ~n17635 ;
  assign n22260 = n3536 & n17346 ;
  assign n22261 = n22259 | n22260 ;
  assign n22262 = n22258 | n22261 ;
  assign n22263 = x29 & ~n22262 ;
  assign n22264 = ( ~x29 & n22256 ) | ( ~x29 & n22262 ) | ( n22256 & n22262 ) ;
  assign n22265 = ( ~n22257 & n22263 ) | ( ~n22257 & n22264 ) | ( n22263 & n22264 ) ;
  assign n22266 = n2760 | n4366 ;
  assign n22267 = n2175 | n2576 ;
  assign n22268 = n22266 | n22267 ;
  assign n22269 = n18231 | n22268 ;
  assign n22270 = n20805 | n22269 ;
  assign n22271 = n20481 | n22270 ;
  assign n22272 = n773 | n957 ;
  assign n22273 = n1102 | n2079 ;
  assign n22274 = n3551 | n22273 ;
  assign n22275 = n22272 | n22274 ;
  assign n22276 = n22271 | n22275 ;
  assign n22277 = n13923 | n18343 ;
  assign n22278 = n22276 | n22277 ;
  assign n22279 = n3273 & n16724 ;
  assign n22280 = n3270 | n22279 ;
  assign n22281 = ( ~n17126 & n22279 ) | ( ~n17126 & n22280 ) | ( n22279 & n22280 ) ;
  assign n22282 = n390 | n22281 ;
  assign n22283 = ( ~n17139 & n22281 ) | ( ~n17139 & n22282 ) | ( n22281 & n22282 ) ;
  assign n22284 = n3274 & n16925 ;
  assign n22285 = n22283 | n22284 ;
  assign n22286 = ( ~n22187 & n22278 ) | ( ~n22187 & n22285 ) | ( n22278 & n22285 ) ;
  assign n22287 = ( n22187 & n22278 ) | ( n22187 & ~n22285 ) | ( n22278 & ~n22285 ) ;
  assign n22288 = ( ~n22278 & n22286 ) | ( ~n22278 & n22287 ) | ( n22286 & n22287 ) ;
  assign n22289 = ( n22189 & ~n22265 ) | ( n22189 & n22288 ) | ( ~n22265 & n22288 ) ;
  assign n22290 = ( n22189 & n22265 ) | ( n22189 & n22288 ) | ( n22265 & n22288 ) ;
  assign n22291 = ( n22265 & n22289 ) | ( n22265 & ~n22290 ) | ( n22289 & ~n22290 ) ;
  assign n22292 = ( ~n22192 & n22255 ) | ( ~n22192 & n22291 ) | ( n22255 & n22291 ) ;
  assign n22293 = ( n22192 & n22255 ) | ( n22192 & n22291 ) | ( n22255 & n22291 ) ;
  assign n22294 = ( n22192 & n22292 ) | ( n22192 & ~n22293 ) | ( n22292 & ~n22293 ) ;
  assign n22295 = ( ~n22195 & n22245 ) | ( ~n22195 & n22294 ) | ( n22245 & n22294 ) ;
  assign n22296 = ( n22195 & n22245 ) | ( n22195 & n22294 ) | ( n22245 & n22294 ) ;
  assign n22297 = ( n22195 & n22295 ) | ( n22195 & ~n22296 ) | ( n22295 & ~n22296 ) ;
  assign n22298 = ( ~n22198 & n22235 ) | ( ~n22198 & n22297 ) | ( n22235 & n22297 ) ;
  assign n22299 = ( n22198 & n22235 ) | ( n22198 & n22297 ) | ( n22235 & n22297 ) ;
  assign n22300 = ( n22198 & n22298 ) | ( n22198 & ~n22299 ) | ( n22298 & ~n22299 ) ;
  assign n22301 = ( ~n22202 & n22225 ) | ( ~n22202 & n22300 ) | ( n22225 & n22300 ) ;
  assign n22302 = ( n22202 & n22225 ) | ( n22202 & n22300 ) | ( n22225 & n22300 ) ;
  assign n22303 = ( n22202 & n22301 ) | ( n22202 & ~n22302 ) | ( n22301 & ~n22302 ) ;
  assign n22304 = n5904 & ~n20095 ;
  assign n22305 = n5908 | n20095 ;
  assign n22306 = ( x14 & n22304 ) | ( x14 & n22305 ) | ( n22304 & n22305 ) ;
  assign n22307 = ( ~n22205 & n22303 ) | ( ~n22205 & n22306 ) | ( n22303 & n22306 ) ;
  assign n22308 = ( n22205 & n22303 ) | ( n22205 & n22306 ) | ( n22303 & n22306 ) ;
  assign n22309 = ( n22205 & n22307 ) | ( n22205 & ~n22308 ) | ( n22307 & ~n22308 ) ;
  assign n22310 = ( ~n22207 & n22211 ) | ( ~n22207 & n22309 ) | ( n22211 & n22309 ) ;
  assign n22311 = ( n22207 & n22211 ) | ( n22207 & n22309 ) | ( n22211 & n22309 ) ;
  assign n22312 = ( n22207 & n22310 ) | ( n22207 & ~n22311 ) | ( n22310 & ~n22311 ) ;
  assign n22313 = n22213 & ~n22312 ;
  assign n22314 = n22213 & n22312 ;
  assign n22315 = ( n22312 & n22313 ) | ( n22312 & ~n22314 ) | ( n22313 & ~n22314 ) ;
  assign n22316 = n5413 & n19916 ;
  assign n22317 = n5417 | n22316 ;
  assign n22318 = ( ~n20095 & n22316 ) | ( ~n20095 & n22317 ) | ( n22316 & n22317 ) ;
  assign n22319 = n5584 & n20091 ;
  assign n22320 = n22318 | n22319 ;
  assign n22321 = x17 & n22320 ;
  assign n22322 = n5418 & ~n20100 ;
  assign n22323 = ( ~x17 & n22320 ) | ( ~x17 & n22322 ) | ( n22320 & n22322 ) ;
  assign n22324 = x17 & ~n22322 ;
  assign n22325 = ( ~n22321 & n22323 ) | ( ~n22321 & n22324 ) | ( n22323 & n22324 ) ;
  assign n22326 = n5232 & ~n19701 ;
  assign n22327 = x20 & n22326 ;
  assign n22328 = n4874 & n19368 ;
  assign n22329 = n4878 | n22328 ;
  assign n22330 = ( n19882 & n22328 ) | ( n19882 & n22329 ) | ( n22328 & n22329 ) ;
  assign n22331 = n4879 | n22330 ;
  assign n22332 = ( ~n19893 & n22330 ) | ( ~n19893 & n22331 ) | ( n22330 & n22331 ) ;
  assign n22333 = x20 & ~n22332 ;
  assign n22334 = ( ~x20 & n22326 ) | ( ~x20 & n22332 ) | ( n22326 & n22332 ) ;
  assign n22335 = ( ~n22327 & n22333 ) | ( ~n22327 & n22334 ) | ( n22333 & n22334 ) ;
  assign n22336 = n4637 & n19248 ;
  assign n22337 = x23 & n22336 ;
  assign n22338 = n4584 & n19177 ;
  assign n22339 = n4649 | n22338 ;
  assign n22340 = ( ~n19315 & n22338 ) | ( ~n19315 & n22339 ) | ( n22338 & n22339 ) ;
  assign n22341 = n4591 | n22340 ;
  assign n22342 = ( ~n19320 & n22340 ) | ( ~n19320 & n22341 ) | ( n22340 & n22341 ) ;
  assign n22343 = x23 & ~n22342 ;
  assign n22344 = ( ~x23 & n22336 ) | ( ~x23 & n22342 ) | ( n22336 & n22342 ) ;
  assign n22345 = ( ~n22337 & n22343 ) | ( ~n22337 & n22344 ) | ( n22343 & n22344 ) ;
  assign n22346 = n4215 & n18730 ;
  assign n22347 = n4200 & ~n18362 ;
  assign n22348 = n2083 & ~n18258 ;
  assign n22349 = n22347 | n22348 ;
  assign n22350 = n22346 | n22349 ;
  assign n22351 = x26 & n22350 ;
  assign n22352 = n4203 & n18735 ;
  assign n22353 = ( ~x26 & n22350 ) | ( ~x26 & n22352 ) | ( n22350 & n22352 ) ;
  assign n22354 = x26 & ~n22352 ;
  assign n22355 = ( ~n22351 & n22353 ) | ( ~n22351 & n22354 ) | ( n22353 & n22354 ) ;
  assign n22356 = n3541 & ~n17976 ;
  assign n22357 = x29 & n22356 ;
  assign n22358 = n3536 & ~n17635 ;
  assign n22359 = n4039 | n22358 ;
  assign n22360 = ( ~n17963 & n22358 ) | ( ~n17963 & n22359 ) | ( n22358 & n22359 ) ;
  assign n22361 = n3501 & n17742 ;
  assign n22362 = n22360 | n22361 ;
  assign n22363 = x29 & ~n22362 ;
  assign n22364 = ( ~x29 & n22356 ) | ( ~x29 & n22362 ) | ( n22356 & n22362 ) ;
  assign n22365 = ( ~n22357 & n22363 ) | ( ~n22357 & n22364 ) | ( n22363 & n22364 ) ;
  assign n22366 = n3273 & n16925 ;
  assign n22367 = n3270 | n22366 ;
  assign n22368 = ( n17346 & n22366 ) | ( n17346 & n22367 ) | ( n22366 & n22367 ) ;
  assign n22369 = n390 | n22368 ;
  assign n22370 = ( ~n17356 & n22368 ) | ( ~n17356 & n22369 ) | ( n22368 & n22369 ) ;
  assign n22371 = n3274 & ~n17126 ;
  assign n22372 = n22370 | n22371 ;
  assign n22373 = n642 | n10137 ;
  assign n22374 = n383 | n2610 ;
  assign n22375 = n22373 | n22374 ;
  assign n22376 = n1339 | n2492 ;
  assign n22377 = n16297 | n22376 ;
  assign n22378 = n2438 | n3325 ;
  assign n22379 = n471 | n3082 ;
  assign n22380 = n22378 | n22379 ;
  assign n22381 = n22377 | n22380 ;
  assign n22382 = n5026 & ~n22381 ;
  assign n22383 = ~n22375 & n22382 ;
  assign n22384 = n2942 | n3903 ;
  assign n22385 = n22383 & ~n22384 ;
  assign n22386 = ( n22278 & ~n22372 ) | ( n22278 & n22385 ) | ( ~n22372 & n22385 ) ;
  assign n22387 = ( n22278 & n22372 ) | ( n22278 & ~n22385 ) | ( n22372 & ~n22385 ) ;
  assign n22388 = ( ~n22278 & n22386 ) | ( ~n22278 & n22387 ) | ( n22386 & n22387 ) ;
  assign n22389 = ( ~n22287 & n22290 ) | ( ~n22287 & n22388 ) | ( n22290 & n22388 ) ;
  assign n22390 = ( n22287 & n22290 ) | ( n22287 & ~n22388 ) | ( n22290 & ~n22388 ) ;
  assign n22391 = ( ~n22290 & n22389 ) | ( ~n22290 & n22390 ) | ( n22389 & n22390 ) ;
  assign n22392 = ( n22355 & ~n22365 ) | ( n22355 & n22391 ) | ( ~n22365 & n22391 ) ;
  assign n22393 = ( n22355 & n22365 ) | ( n22355 & ~n22391 ) | ( n22365 & ~n22391 ) ;
  assign n22394 = ( ~n22355 & n22392 ) | ( ~n22355 & n22393 ) | ( n22392 & n22393 ) ;
  assign n22395 = ( n22293 & n22345 ) | ( n22293 & ~n22394 ) | ( n22345 & ~n22394 ) ;
  assign n22396 = ( ~n22293 & n22345 ) | ( ~n22293 & n22394 ) | ( n22345 & n22394 ) ;
  assign n22397 = ( ~n22345 & n22395 ) | ( ~n22345 & n22396 ) | ( n22395 & n22396 ) ;
  assign n22398 = ( n22296 & n22335 ) | ( n22296 & ~n22397 ) | ( n22335 & ~n22397 ) ;
  assign n22399 = ( ~n22296 & n22335 ) | ( ~n22296 & n22397 ) | ( n22335 & n22397 ) ;
  assign n22400 = ( ~n22335 & n22398 ) | ( ~n22335 & n22399 ) | ( n22398 & n22399 ) ;
  assign n22401 = ( n22299 & n22325 ) | ( n22299 & ~n22400 ) | ( n22325 & ~n22400 ) ;
  assign n22402 = ( ~n22299 & n22325 ) | ( ~n22299 & n22400 ) | ( n22325 & n22400 ) ;
  assign n22403 = ( ~n22325 & n22401 ) | ( ~n22325 & n22402 ) | ( n22401 & n22402 ) ;
  assign n22404 = ( ~x14 & n22302 ) | ( ~x14 & n22403 ) | ( n22302 & n22403 ) ;
  assign n22405 = ( x14 & n22302 ) | ( x14 & ~n22403 ) | ( n22302 & ~n22403 ) ;
  assign n22406 = ( ~n22302 & n22404 ) | ( ~n22302 & n22405 ) | ( n22404 & n22405 ) ;
  assign n22407 = ( n22308 & n22311 ) | ( n22308 & ~n22406 ) | ( n22311 & ~n22406 ) ;
  assign n22408 = ( ~n22308 & n22311 ) | ( ~n22308 & n22406 ) | ( n22311 & n22406 ) ;
  assign n22409 = ( ~n22311 & n22407 ) | ( ~n22311 & n22408 ) | ( n22407 & n22408 ) ;
  assign n22410 = n22314 & ~n22409 ;
  assign n22411 = ~n22314 & n22409 ;
  assign n22412 = n22410 | n22411 ;
  assign n22413 = n5232 & n19882 ;
  assign n22414 = x20 & n22413 ;
  assign n22415 = n4874 & ~n19701 ;
  assign n22416 = n4878 | n22415 ;
  assign n22417 = ( n19916 & n22415 ) | ( n19916 & n22416 ) | ( n22415 & n22416 ) ;
  assign n22418 = n4879 | n22417 ;
  assign n22419 = ( n19920 & n22417 ) | ( n19920 & n22418 ) | ( n22417 & n22418 ) ;
  assign n22420 = x20 & ~n22419 ;
  assign n22421 = ( ~x20 & n22413 ) | ( ~x20 & n22419 ) | ( n22413 & n22419 ) ;
  assign n22422 = ( ~n22414 & n22420 ) | ( ~n22414 & n22421 ) | ( n22420 & n22421 ) ;
  assign n22423 = n4591 & ~n19374 ;
  assign n22424 = x23 & n22423 ;
  assign n22425 = n4584 & n19248 ;
  assign n22426 = n4649 | n22425 ;
  assign n22427 = ( n19368 & n22425 ) | ( n19368 & n22426 ) | ( n22425 & n22426 ) ;
  assign n22428 = n4637 & ~n19315 ;
  assign n22429 = n22427 | n22428 ;
  assign n22430 = x23 & ~n22429 ;
  assign n22431 = ( ~x23 & n22423 ) | ( ~x23 & n22429 ) | ( n22423 & n22429 ) ;
  assign n22432 = ( ~n22424 & n22430 ) | ( ~n22424 & n22431 ) | ( n22430 & n22431 ) ;
  assign n22433 = n4215 & n19177 ;
  assign n22434 = n4200 & n18730 ;
  assign n22435 = n2083 & ~n18362 ;
  assign n22436 = n22434 | n22435 ;
  assign n22437 = n22433 | n22436 ;
  assign n22438 = x26 & n22437 ;
  assign n22439 = n4203 & ~n19182 ;
  assign n22440 = ( ~x26 & n22437 ) | ( ~x26 & n22439 ) | ( n22437 & n22439 ) ;
  assign n22441 = x26 & ~n22439 ;
  assign n22442 = ( ~n22438 & n22440 ) | ( ~n22438 & n22441 ) | ( n22440 & n22441 ) ;
  assign n22443 = n3501 & ~n17963 ;
  assign n22444 = x29 & n22443 ;
  assign n22445 = n3536 & n17742 ;
  assign n22446 = n4039 | n22445 ;
  assign n22447 = ( ~n18258 & n22445 ) | ( ~n18258 & n22446 ) | ( n22445 & n22446 ) ;
  assign n22448 = n3541 | n22447 ;
  assign n22449 = ( n18268 & n22447 ) | ( n18268 & n22448 ) | ( n22447 & n22448 ) ;
  assign n22450 = x29 & ~n22449 ;
  assign n22451 = ( ~x29 & n22443 ) | ( ~x29 & n22449 ) | ( n22443 & n22449 ) ;
  assign n22452 = ( ~n22444 & n22450 ) | ( ~n22444 & n22451 ) | ( n22450 & n22451 ) ;
  assign n22453 = n3273 & ~n17126 ;
  assign n22454 = n3270 | n22453 ;
  assign n22455 = ( ~n17635 & n22453 ) | ( ~n17635 & n22454 ) | ( n22453 & n22454 ) ;
  assign n22456 = n390 | n22455 ;
  assign n22457 = ( ~n17646 & n22455 ) | ( ~n17646 & n22456 ) | ( n22455 & n22456 ) ;
  assign n22458 = n3274 & n17346 ;
  assign n22459 = n22457 | n22458 ;
  assign n22460 = n996 | n3304 ;
  assign n22461 = n1745 | n2922 ;
  assign n22462 = n3995 | n22461 ;
  assign n22463 = n22460 | n22462 ;
  assign n22464 = n2719 | n2947 ;
  assign n22465 = n22463 | n22464 ;
  assign n22466 = n1648 | n12843 ;
  assign n22467 = n22465 | n22466 ;
  assign n22468 = n6030 & ~n22467 ;
  assign n22469 = ~n1883 & n22468 ;
  assign n22470 = ~n16900 & n22469 ;
  assign n22471 = ( x14 & n22278 ) | ( x14 & ~n22470 ) | ( n22278 & ~n22470 ) ;
  assign n22472 = ( x14 & ~n22278 ) | ( x14 & n22470 ) | ( ~n22278 & n22470 ) ;
  assign n22473 = ( ~x14 & n22471 ) | ( ~x14 & n22472 ) | ( n22471 & n22472 ) ;
  assign n22474 = ( ~n22386 & n22459 ) | ( ~n22386 & n22473 ) | ( n22459 & n22473 ) ;
  assign n22475 = ( n22386 & n22459 ) | ( n22386 & n22473 ) | ( n22459 & n22473 ) ;
  assign n22476 = ( n22386 & n22474 ) | ( n22386 & ~n22475 ) | ( n22474 & ~n22475 ) ;
  assign n22477 = ( n22389 & n22452 ) | ( n22389 & ~n22476 ) | ( n22452 & ~n22476 ) ;
  assign n22478 = ( ~n22389 & n22452 ) | ( ~n22389 & n22476 ) | ( n22452 & n22476 ) ;
  assign n22479 = ( ~n22452 & n22477 ) | ( ~n22452 & n22478 ) | ( n22477 & n22478 ) ;
  assign n22480 = ( n22393 & n22442 ) | ( n22393 & ~n22479 ) | ( n22442 & ~n22479 ) ;
  assign n22481 = ( n22393 & ~n22442 ) | ( n22393 & n22479 ) | ( ~n22442 & n22479 ) ;
  assign n22482 = ( ~n22393 & n22480 ) | ( ~n22393 & n22481 ) | ( n22480 & n22481 ) ;
  assign n22483 = ( n22395 & n22432 ) | ( n22395 & ~n22482 ) | ( n22432 & ~n22482 ) ;
  assign n22484 = ( ~n22395 & n22432 ) | ( ~n22395 & n22482 ) | ( n22432 & n22482 ) ;
  assign n22485 = ( ~n22432 & n22483 ) | ( ~n22432 & n22484 ) | ( n22483 & n22484 ) ;
  assign n22486 = ( n22398 & n22422 ) | ( n22398 & ~n22485 ) | ( n22422 & ~n22485 ) ;
  assign n22487 = ( n22398 & ~n22422 ) | ( n22398 & n22485 ) | ( ~n22422 & n22485 ) ;
  assign n22488 = ( ~n22398 & n22486 ) | ( ~n22398 & n22487 ) | ( n22486 & n22487 ) ;
  assign n22489 = n5584 & ~n20095 ;
  assign n22490 = n5413 & n20091 ;
  assign n22491 = n22489 | n22490 ;
  assign n22492 = x17 & n22491 ;
  assign n22493 = n5418 & ~n20097 ;
  assign n22494 = ( ~x17 & n22491 ) | ( ~x17 & n22493 ) | ( n22491 & n22493 ) ;
  assign n22495 = x17 & ~n22493 ;
  assign n22496 = ( ~n22492 & n22494 ) | ( ~n22492 & n22495 ) | ( n22494 & n22495 ) ;
  assign n22497 = ( n22401 & n22488 ) | ( n22401 & n22496 ) | ( n22488 & n22496 ) ;
  assign n22498 = ( n22401 & ~n22488 ) | ( n22401 & n22496 ) | ( ~n22488 & n22496 ) ;
  assign n22499 = ( n22488 & ~n22497 ) | ( n22488 & n22498 ) | ( ~n22497 & n22498 ) ;
  assign n22500 = ( n22405 & n22407 ) | ( n22405 & ~n22499 ) | ( n22407 & ~n22499 ) ;
  assign n22501 = ( ~n22405 & n22407 ) | ( ~n22405 & n22499 ) | ( n22407 & n22499 ) ;
  assign n22502 = ( ~n22407 & n22500 ) | ( ~n22407 & n22501 ) | ( n22500 & n22501 ) ;
  assign n22503 = n22410 & ~n22502 ;
  assign n22504 = ~n22410 & n22502 ;
  assign n22505 = n22503 | n22504 ;
  assign n22506 = n5232 & n19916 ;
  assign n22507 = x20 & n22506 ;
  assign n22508 = n4874 & n19882 ;
  assign n22509 = n4878 | n22508 ;
  assign n22510 = ( n20091 & n22508 ) | ( n20091 & n22509 ) | ( n22508 & n22509 ) ;
  assign n22511 = n4879 | n22510 ;
  assign n22512 = ( n20101 & n22510 ) | ( n20101 & n22511 ) | ( n22510 & n22511 ) ;
  assign n22513 = x20 & ~n22512 ;
  assign n22514 = ( ~x20 & n22506 ) | ( ~x20 & n22512 ) | ( n22506 & n22512 ) ;
  assign n22515 = ( ~n22507 & n22513 ) | ( ~n22507 & n22514 ) | ( n22513 & n22514 ) ;
  assign n22516 = n4649 & ~n19701 ;
  assign n22517 = n4591 | n22516 ;
  assign n22518 = ( ~n19706 & n22516 ) | ( ~n19706 & n22517 ) | ( n22516 & n22517 ) ;
  assign n22519 = n4637 & n19368 ;
  assign n22520 = n22518 | n22519 ;
  assign n22521 = n4583 & ~n19315 ;
  assign n22522 = n4584 & ~n19315 ;
  assign n22523 = x23 & ~n22522 ;
  assign n22524 = ( ~n22520 & n22521 ) | ( ~n22520 & n22523 ) | ( n22521 & n22523 ) ;
  assign n22525 = n22520 | n22523 ;
  assign n22526 = ( ~x23 & n22524 ) | ( ~x23 & n22525 ) | ( n22524 & n22525 ) ;
  assign n22527 = n4215 & n19248 ;
  assign n22528 = n4200 & n19177 ;
  assign n22529 = n2083 & n18730 ;
  assign n22530 = n22528 | n22529 ;
  assign n22531 = n22527 | n22530 ;
  assign n22532 = x26 & n22531 ;
  assign n22533 = n4203 & n19253 ;
  assign n22534 = ( ~x26 & n22531 ) | ( ~x26 & n22533 ) | ( n22531 & n22533 ) ;
  assign n22535 = x26 & ~n22533 ;
  assign n22536 = ( ~n22532 & n22534 ) | ( ~n22532 & n22535 ) | ( n22534 & n22535 ) ;
  assign n22537 = n3541 & ~n18373 ;
  assign n22538 = x29 & n22537 ;
  assign n22539 = n3536 & ~n17963 ;
  assign n22540 = n4039 | n22539 ;
  assign n22541 = ( ~n18362 & n22539 ) | ( ~n18362 & n22540 ) | ( n22539 & n22540 ) ;
  assign n22542 = n3501 & ~n18258 ;
  assign n22543 = n22541 | n22542 ;
  assign n22544 = x29 & ~n22543 ;
  assign n22545 = ( ~x29 & n22537 ) | ( ~x29 & n22543 ) | ( n22537 & n22543 ) ;
  assign n22546 = ( ~n22538 & n22544 ) | ( ~n22538 & n22545 ) | ( n22544 & n22545 ) ;
  assign n22547 = n3274 & ~n17635 ;
  assign n22548 = n3273 & n17346 ;
  assign n22549 = n22547 | n22548 ;
  assign n22550 = n390 | n22549 ;
  assign n22551 = ( ~n17749 & n22549 ) | ( ~n17749 & n22550 ) | ( n22549 & n22550 ) ;
  assign n22552 = n3270 & n17742 ;
  assign n22553 = n22551 | n22552 ;
  assign n22554 = n5443 | n15514 ;
  assign n22555 = n290 | n2011 ;
  assign n22556 = n82 | n1649 ;
  assign n22557 = n12679 | n22556 ;
  assign n22558 = n22555 | n22557 ;
  assign n22559 = n22554 | n22558 ;
  assign n22560 = n3048 & ~n22559 ;
  assign n22561 = n1793 | n2321 ;
  assign n22562 = n683 | n2754 ;
  assign n22563 = n22561 | n22562 ;
  assign n22564 = n19447 | n22563 ;
  assign n22565 = n646 | n22564 ;
  assign n22566 = n4933 | n22565 ;
  assign n22567 = n22560 & ~n22566 ;
  assign n22568 = ( ~n22472 & n22553 ) | ( ~n22472 & n22567 ) | ( n22553 & n22567 ) ;
  assign n22569 = ( n22472 & n22553 ) | ( n22472 & ~n22567 ) | ( n22553 & ~n22567 ) ;
  assign n22570 = ( ~n22553 & n22568 ) | ( ~n22553 & n22569 ) | ( n22568 & n22569 ) ;
  assign n22571 = ( n22474 & n22546 ) | ( n22474 & ~n22570 ) | ( n22546 & ~n22570 ) ;
  assign n22572 = ( ~n22474 & n22546 ) | ( ~n22474 & n22570 ) | ( n22546 & n22570 ) ;
  assign n22573 = ( ~n22546 & n22571 ) | ( ~n22546 & n22572 ) | ( n22571 & n22572 ) ;
  assign n22574 = ( n22477 & n22536 ) | ( n22477 & ~n22573 ) | ( n22536 & ~n22573 ) ;
  assign n22575 = ( ~n22477 & n22536 ) | ( ~n22477 & n22573 ) | ( n22536 & n22573 ) ;
  assign n22576 = ( ~n22536 & n22574 ) | ( ~n22536 & n22575 ) | ( n22574 & n22575 ) ;
  assign n22577 = ( n22480 & n22526 ) | ( n22480 & ~n22576 ) | ( n22526 & ~n22576 ) ;
  assign n22578 = ( ~n22480 & n22526 ) | ( ~n22480 & n22576 ) | ( n22526 & n22576 ) ;
  assign n22579 = ( ~n22526 & n22577 ) | ( ~n22526 & n22578 ) | ( n22577 & n22578 ) ;
  assign n22580 = ( n22483 & n22515 ) | ( n22483 & ~n22579 ) | ( n22515 & ~n22579 ) ;
  assign n22581 = ( ~n22483 & n22515 ) | ( ~n22483 & n22579 ) | ( n22515 & n22579 ) ;
  assign n22582 = ( ~n22515 & n22580 ) | ( ~n22515 & n22581 ) | ( n22580 & n22581 ) ;
  assign n22583 = n5408 & ~n20095 ;
  assign n22584 = n5412 | n20095 ;
  assign n22585 = ( x17 & n22583 ) | ( x17 & n22584 ) | ( n22583 & n22584 ) ;
  assign n22586 = ( n22486 & n22582 ) | ( n22486 & n22585 ) | ( n22582 & n22585 ) ;
  assign n22587 = ( n22486 & ~n22582 ) | ( n22486 & n22585 ) | ( ~n22582 & n22585 ) ;
  assign n22588 = ( n22582 & ~n22586 ) | ( n22582 & n22587 ) | ( ~n22586 & n22587 ) ;
  assign n22589 = ( n22498 & n22500 ) | ( n22498 & ~n22588 ) | ( n22500 & ~n22588 ) ;
  assign n22590 = ( ~n22498 & n22500 ) | ( ~n22498 & n22588 ) | ( n22500 & n22588 ) ;
  assign n22591 = ( ~n22500 & n22589 ) | ( ~n22500 & n22590 ) | ( n22589 & n22590 ) ;
  assign n22592 = n22503 & ~n22591 ;
  assign n22593 = ~n22503 & n22591 ;
  assign n22594 = n22592 | n22593 ;
  assign n22595 = n4879 & ~n20100 ;
  assign n22596 = x20 & n22595 ;
  assign n22597 = n4874 & n19916 ;
  assign n22598 = n4878 | n22597 ;
  assign n22599 = ( ~n20095 & n22597 ) | ( ~n20095 & n22598 ) | ( n22597 & n22598 ) ;
  assign n22600 = n5232 & n20091 ;
  assign n22601 = n22599 | n22600 ;
  assign n22602 = x20 & ~n22601 ;
  assign n22603 = ( ~x20 & n22595 ) | ( ~x20 & n22601 ) | ( n22595 & n22601 ) ;
  assign n22604 = ( ~n22596 & n22602 ) | ( ~n22596 & n22603 ) | ( n22602 & n22603 ) ;
  assign n22605 = n4637 & ~n19701 ;
  assign n22606 = x23 & n22605 ;
  assign n22607 = n4584 & n19368 ;
  assign n22608 = n4649 | n22607 ;
  assign n22609 = ( n19882 & n22607 ) | ( n19882 & n22608 ) | ( n22607 & n22608 ) ;
  assign n22610 = n4591 | n22609 ;
  assign n22611 = ( ~n19893 & n22609 ) | ( ~n19893 & n22610 ) | ( n22609 & n22610 ) ;
  assign n22612 = x23 & ~n22611 ;
  assign n22613 = ( ~x23 & n22605 ) | ( ~x23 & n22611 ) | ( n22605 & n22611 ) ;
  assign n22614 = ( ~n22606 & n22612 ) | ( ~n22606 & n22613 ) | ( n22612 & n22613 ) ;
  assign n22615 = n4215 & ~n19315 ;
  assign n22616 = n4200 & n19248 ;
  assign n22617 = n2083 & n19177 ;
  assign n22618 = n22616 | n22617 ;
  assign n22619 = n22615 | n22618 ;
  assign n22620 = x26 & n22619 ;
  assign n22621 = n4203 & ~n19320 ;
  assign n22622 = ( ~x26 & n22619 ) | ( ~x26 & n22621 ) | ( n22619 & n22621 ) ;
  assign n22623 = x26 & ~n22621 ;
  assign n22624 = ( ~n22620 & n22622 ) | ( ~n22620 & n22623 ) | ( n22622 & n22623 ) ;
  assign n22625 = n3501 & ~n18362 ;
  assign n22626 = x29 & n22625 ;
  assign n22627 = n3536 & ~n18258 ;
  assign n22628 = n4039 | n22627 ;
  assign n22629 = ( n18730 & n22627 ) | ( n18730 & n22628 ) | ( n22627 & n22628 ) ;
  assign n22630 = n3541 | n22629 ;
  assign n22631 = ( n18735 & n22629 ) | ( n18735 & n22630 ) | ( n22629 & n22630 ) ;
  assign n22632 = x29 & ~n22631 ;
  assign n22633 = ( ~x29 & n22625 ) | ( ~x29 & n22631 ) | ( n22625 & n22631 ) ;
  assign n22634 = ( ~n22626 & n22632 ) | ( ~n22626 & n22633 ) | ( n22632 & n22633 ) ;
  assign n22635 = n2019 | n2470 ;
  assign n22636 = n4008 | n22635 ;
  assign n22637 = n647 | n1102 ;
  assign n22638 = n1177 | n22637 ;
  assign n22639 = n22636 | n22638 ;
  assign n22640 = n438 | n2916 ;
  assign n22641 = n22639 | n22640 ;
  assign n22642 = n2895 | n4284 ;
  assign n22643 = n13194 | n14656 ;
  assign n22644 = n22642 | n22643 ;
  assign n22645 = n22641 | n22644 ;
  assign n22646 = n3371 | n22645 ;
  assign n22647 = n1790 | n5056 ;
  assign n22648 = n22646 | n22647 ;
  assign n22649 = ( n22567 & n22568 ) | ( n22567 & ~n22648 ) | ( n22568 & ~n22648 ) ;
  assign n22650 = ( n22472 & ~n22569 ) | ( n22472 & n22648 ) | ( ~n22569 & n22648 ) ;
  assign n22651 = ( ~n22567 & n22649 ) | ( ~n22567 & n22650 ) | ( n22649 & n22650 ) ;
  assign n22652 = n3270 & ~n17963 ;
  assign n22653 = n3274 & n17742 ;
  assign n22654 = n3273 & ~n17635 ;
  assign n22655 = n22653 | n22654 ;
  assign n22656 = n22652 | n22655 ;
  assign n22657 = n390 & ~n17976 ;
  assign n22658 = n22656 | n22657 ;
  assign n22659 = ( ~n22634 & n22651 ) | ( ~n22634 & n22658 ) | ( n22651 & n22658 ) ;
  assign n22660 = ( n22634 & n22651 ) | ( n22634 & n22658 ) | ( n22651 & n22658 ) ;
  assign n22661 = ( n22634 & n22659 ) | ( n22634 & ~n22660 ) | ( n22659 & ~n22660 ) ;
  assign n22662 = ( ~n22571 & n22624 ) | ( ~n22571 & n22661 ) | ( n22624 & n22661 ) ;
  assign n22663 = ( n22571 & n22624 ) | ( n22571 & n22661 ) | ( n22624 & n22661 ) ;
  assign n22664 = ( n22571 & n22662 ) | ( n22571 & ~n22663 ) | ( n22662 & ~n22663 ) ;
  assign n22665 = ( n22574 & ~n22614 ) | ( n22574 & n22664 ) | ( ~n22614 & n22664 ) ;
  assign n22666 = ( n22574 & n22614 ) | ( n22574 & n22664 ) | ( n22614 & n22664 ) ;
  assign n22667 = ( n22614 & n22665 ) | ( n22614 & ~n22666 ) | ( n22665 & ~n22666 ) ;
  assign n22668 = ( n22577 & ~n22604 ) | ( n22577 & n22667 ) | ( ~n22604 & n22667 ) ;
  assign n22669 = ( n22577 & n22604 ) | ( n22577 & n22667 ) | ( n22604 & n22667 ) ;
  assign n22670 = ( n22604 & n22668 ) | ( n22604 & ~n22669 ) | ( n22668 & ~n22669 ) ;
  assign n22671 = ( ~x17 & n22580 ) | ( ~x17 & n22670 ) | ( n22580 & n22670 ) ;
  assign n22672 = ( x17 & n22580 ) | ( x17 & n22670 ) | ( n22580 & n22670 ) ;
  assign n22673 = ( x17 & n22671 ) | ( x17 & ~n22672 ) | ( n22671 & ~n22672 ) ;
  assign n22674 = ( n22587 & ~n22589 ) | ( n22587 & n22673 ) | ( ~n22589 & n22673 ) ;
  assign n22675 = ( n22587 & n22589 ) | ( n22587 & n22673 ) | ( n22589 & n22673 ) ;
  assign n22676 = ( n22589 & n22674 ) | ( n22589 & ~n22675 ) | ( n22674 & ~n22675 ) ;
  assign n22677 = n22592 & ~n22676 ;
  assign n22678 = n22592 & n22676 ;
  assign n22679 = ( n22676 & n22677 ) | ( n22676 & ~n22678 ) | ( n22677 & ~n22678 ) ;
  assign n22680 = n4637 & n19882 ;
  assign n22681 = x23 & n22680 ;
  assign n22682 = n4584 & ~n19701 ;
  assign n22683 = n4649 | n22682 ;
  assign n22684 = ( n19916 & n22682 ) | ( n19916 & n22683 ) | ( n22682 & n22683 ) ;
  assign n22685 = n4591 | n22684 ;
  assign n22686 = ( n19920 & n22684 ) | ( n19920 & n22685 ) | ( n22684 & n22685 ) ;
  assign n22687 = x23 & ~n22686 ;
  assign n22688 = ( ~x23 & n22680 ) | ( ~x23 & n22686 ) | ( n22680 & n22686 ) ;
  assign n22689 = ( ~n22681 & n22687 ) | ( ~n22681 & n22688 ) | ( n22687 & n22688 ) ;
  assign n22690 = n4215 & n19368 ;
  assign n22691 = n4200 & ~n19315 ;
  assign n22692 = n2083 & n19248 ;
  assign n22693 = n22691 | n22692 ;
  assign n22694 = n22690 | n22693 ;
  assign n22695 = x26 & n22694 ;
  assign n22696 = n4203 & ~n19374 ;
  assign n22697 = ( ~x26 & n22694 ) | ( ~x26 & n22696 ) | ( n22694 & n22696 ) ;
  assign n22698 = x26 & ~n22696 ;
  assign n22699 = ( ~n22695 & n22697 ) | ( ~n22695 & n22698 ) | ( n22697 & n22698 ) ;
  assign n22700 = n3541 & ~n19182 ;
  assign n22701 = x29 & n22700 ;
  assign n22702 = n3536 & ~n18362 ;
  assign n22703 = n4039 | n22702 ;
  assign n22704 = ( n19177 & n22702 ) | ( n19177 & n22703 ) | ( n22702 & n22703 ) ;
  assign n22705 = n3501 & n18730 ;
  assign n22706 = n22704 | n22705 ;
  assign n22707 = x29 & ~n22706 ;
  assign n22708 = ( ~x29 & n22700 ) | ( ~x29 & n22706 ) | ( n22700 & n22706 ) ;
  assign n22709 = ( ~n22701 & n22707 ) | ( ~n22701 & n22708 ) | ( n22707 & n22708 ) ;
  assign n22710 = n3273 & n17742 ;
  assign n22711 = n3270 | n22710 ;
  assign n22712 = ( ~n18258 & n22710 ) | ( ~n18258 & n22711 ) | ( n22710 & n22711 ) ;
  assign n22713 = n390 | n22712 ;
  assign n22714 = ( n18268 & n22712 ) | ( n18268 & n22713 ) | ( n22712 & n22713 ) ;
  assign n22715 = n3274 & ~n17963 ;
  assign n22716 = n22714 | n22715 ;
  assign n22717 = n1199 | n1571 ;
  assign n22718 = n1738 | n22717 ;
  assign n22719 = n4135 | n22718 ;
  assign n22720 = n21566 | n22719 ;
  assign n22721 = n3018 | n19457 ;
  assign n22722 = n22720 | n22721 ;
  assign n22723 = n1596 | n17913 ;
  assign n22724 = n22722 | n22723 ;
  assign n22725 = n1274 | n22724 ;
  assign n22726 = n4115 | n4821 ;
  assign n22727 = n22725 | n22726 ;
  assign n22728 = ( x17 & n22648 ) | ( x17 & n22727 ) | ( n22648 & n22727 ) ;
  assign n22729 = ( ~x17 & n22648 ) | ( ~x17 & n22727 ) | ( n22648 & n22727 ) ;
  assign n22730 = ( x17 & ~n22728 ) | ( x17 & n22729 ) | ( ~n22728 & n22729 ) ;
  assign n22731 = ( n22650 & ~n22716 ) | ( n22650 & n22730 ) | ( ~n22716 & n22730 ) ;
  assign n22732 = ( n22650 & n22716 ) | ( n22650 & n22730 ) | ( n22716 & n22730 ) ;
  assign n22733 = ( n22716 & n22731 ) | ( n22716 & ~n22732 ) | ( n22731 & ~n22732 ) ;
  assign n22734 = ( ~n22660 & n22709 ) | ( ~n22660 & n22733 ) | ( n22709 & n22733 ) ;
  assign n22735 = ( n22660 & n22709 ) | ( n22660 & n22733 ) | ( n22709 & n22733 ) ;
  assign n22736 = ( n22660 & n22734 ) | ( n22660 & ~n22735 ) | ( n22734 & ~n22735 ) ;
  assign n22737 = ( n22663 & ~n22699 ) | ( n22663 & n22736 ) | ( ~n22699 & n22736 ) ;
  assign n22738 = ( n22663 & n22699 ) | ( n22663 & n22736 ) | ( n22699 & n22736 ) ;
  assign n22739 = ( n22699 & n22737 ) | ( n22699 & ~n22738 ) | ( n22737 & ~n22738 ) ;
  assign n22740 = ( n22666 & n22689 ) | ( n22666 & n22739 ) | ( n22689 & n22739 ) ;
  assign n22741 = ( n22666 & ~n22689 ) | ( n22666 & n22739 ) | ( ~n22689 & n22739 ) ;
  assign n22742 = ( n22689 & ~n22740 ) | ( n22689 & n22741 ) | ( ~n22740 & n22741 ) ;
  assign n22743 = n5232 & ~n20095 ;
  assign n22744 = n4874 & n20091 ;
  assign n22745 = n22743 | n22744 ;
  assign n22746 = x20 & n22745 ;
  assign n22747 = n4879 & ~n20097 ;
  assign n22748 = ( ~x20 & n22745 ) | ( ~x20 & n22747 ) | ( n22745 & n22747 ) ;
  assign n22749 = x20 & ~n22747 ;
  assign n22750 = ( ~n22746 & n22748 ) | ( ~n22746 & n22749 ) | ( n22748 & n22749 ) ;
  assign n22751 = ( ~n22669 & n22742 ) | ( ~n22669 & n22750 ) | ( n22742 & n22750 ) ;
  assign n22752 = ( n22669 & n22742 ) | ( n22669 & n22750 ) | ( n22742 & n22750 ) ;
  assign n22753 = ( n22669 & n22751 ) | ( n22669 & ~n22752 ) | ( n22751 & ~n22752 ) ;
  assign n22754 = ( n22672 & n22675 ) | ( n22672 & n22753 ) | ( n22675 & n22753 ) ;
  assign n22755 = ( n22672 & ~n22675 ) | ( n22672 & n22753 ) | ( ~n22675 & n22753 ) ;
  assign n22756 = ( n22675 & ~n22754 ) | ( n22675 & n22755 ) | ( ~n22754 & n22755 ) ;
  assign n22757 = n22678 & ~n22756 ;
  assign n22758 = n22678 & n22756 ;
  assign n22759 = ( n22756 & n22757 ) | ( n22756 & ~n22758 ) | ( n22757 & ~n22758 ) ;
  assign n22760 = n4215 & ~n19701 ;
  assign n22761 = n4200 & n19368 ;
  assign n22762 = n2083 & ~n19315 ;
  assign n22763 = n22761 | n22762 ;
  assign n22764 = n22760 | n22763 ;
  assign n22765 = x26 & n22764 ;
  assign n22766 = n4203 & ~n19706 ;
  assign n22767 = ( ~x26 & n22764 ) | ( ~x26 & n22766 ) | ( n22764 & n22766 ) ;
  assign n22768 = x26 & ~n22766 ;
  assign n22769 = ( ~n22765 & n22767 ) | ( ~n22765 & n22768 ) | ( n22767 & n22768 ) ;
  assign n22770 = n3501 & n19177 ;
  assign n22771 = x29 & n22770 ;
  assign n22772 = n3536 & n18730 ;
  assign n22773 = n4039 | n22772 ;
  assign n22774 = ( n19248 & n22772 ) | ( n19248 & n22773 ) | ( n22772 & n22773 ) ;
  assign n22775 = n3541 | n22774 ;
  assign n22776 = ( n19253 & n22774 ) | ( n19253 & n22775 ) | ( n22774 & n22775 ) ;
  assign n22777 = x29 & ~n22776 ;
  assign n22778 = ( ~x29 & n22770 ) | ( ~x29 & n22776 ) | ( n22770 & n22776 ) ;
  assign n22779 = ( ~n22771 & n22777 ) | ( ~n22771 & n22778 ) | ( n22777 & n22778 ) ;
  assign n22780 = n164 | n1041 ;
  assign n22781 = n413 | n22780 ;
  assign n22782 = n1380 | n22781 ;
  assign n22783 = n4771 | n22782 ;
  assign n22784 = n888 | n22783 ;
  assign n22785 = n2952 | n22784 ;
  assign n22786 = n1253 | n4253 ;
  assign n22787 = n1159 | n22786 ;
  assign n22788 = n3051 | n22787 ;
  assign n22789 = n18698 | n22788 ;
  assign n22790 = n22785 | n22789 ;
  assign n22791 = n6188 | n22790 ;
  assign n22792 = n21704 & ~n22791 ;
  assign n22793 = n3273 & ~n17963 ;
  assign n22794 = n3270 | n22793 ;
  assign n22795 = ( ~n18362 & n22793 ) | ( ~n18362 & n22794 ) | ( n22793 & n22794 ) ;
  assign n22796 = n390 | n22795 ;
  assign n22797 = ( ~n18373 & n22795 ) | ( ~n18373 & n22796 ) | ( n22795 & n22796 ) ;
  assign n22798 = n3274 & ~n18258 ;
  assign n22799 = n22797 | n22798 ;
  assign n22800 = ( n22729 & ~n22792 ) | ( n22729 & n22799 ) | ( ~n22792 & n22799 ) ;
  assign n22801 = ( n22729 & n22792 ) | ( n22729 & n22799 ) | ( n22792 & n22799 ) ;
  assign n22802 = ( n22792 & n22800 ) | ( n22792 & ~n22801 ) | ( n22800 & ~n22801 ) ;
  assign n22803 = ( ~n22731 & n22779 ) | ( ~n22731 & n22802 ) | ( n22779 & n22802 ) ;
  assign n22804 = ( n22731 & n22779 ) | ( n22731 & ~n22802 ) | ( n22779 & ~n22802 ) ;
  assign n22805 = ( ~n22779 & n22803 ) | ( ~n22779 & n22804 ) | ( n22803 & n22804 ) ;
  assign n22806 = ( n22735 & n22769 ) | ( n22735 & ~n22805 ) | ( n22769 & ~n22805 ) ;
  assign n22807 = ( ~n22735 & n22769 ) | ( ~n22735 & n22805 ) | ( n22769 & n22805 ) ;
  assign n22808 = ( ~n22769 & n22806 ) | ( ~n22769 & n22807 ) | ( n22806 & n22807 ) ;
  assign n22809 = n4649 & n20091 ;
  assign n22810 = n4591 | n22809 ;
  assign n22811 = ( n20101 & n22809 ) | ( n20101 & n22810 ) | ( n22809 & n22810 ) ;
  assign n22812 = n4637 & n19916 ;
  assign n22813 = n22811 | n22812 ;
  assign n22814 = n4583 & n19882 ;
  assign n22815 = n4584 & n19882 ;
  assign n22816 = x23 & ~n22815 ;
  assign n22817 = ( ~n22813 & n22814 ) | ( ~n22813 & n22816 ) | ( n22814 & n22816 ) ;
  assign n22818 = n22813 | n22816 ;
  assign n22819 = ( ~x23 & n22817 ) | ( ~x23 & n22818 ) | ( n22817 & n22818 ) ;
  assign n22820 = ( n22738 & n22808 ) | ( n22738 & n22819 ) | ( n22808 & n22819 ) ;
  assign n22821 = ( n22738 & ~n22808 ) | ( n22738 & n22819 ) | ( ~n22808 & n22819 ) ;
  assign n22822 = ( n22808 & ~n22820 ) | ( n22808 & n22821 ) | ( ~n22820 & n22821 ) ;
  assign n22823 = n4869 | n20095 ;
  assign n22824 = n4873 | n20095 ;
  assign n22825 = ( x20 & n22823 ) | ( x20 & ~n22824 ) | ( n22823 & ~n22824 ) ;
  assign n22826 = ( n22740 & n22822 ) | ( n22740 & n22825 ) | ( n22822 & n22825 ) ;
  assign n22827 = ( n22740 & ~n22822 ) | ( n22740 & n22825 ) | ( ~n22822 & n22825 ) ;
  assign n22828 = ( n22822 & ~n22826 ) | ( n22822 & n22827 ) | ( ~n22826 & n22827 ) ;
  assign n22829 = ( n22752 & n22754 ) | ( n22752 & ~n22828 ) | ( n22754 & ~n22828 ) ;
  assign n22830 = ( ~n22752 & n22754 ) | ( ~n22752 & n22828 ) | ( n22754 & n22828 ) ;
  assign n22831 = ( ~n22754 & n22829 ) | ( ~n22754 & n22830 ) | ( n22829 & n22830 ) ;
  assign n22832 = n22758 & ~n22831 ;
  assign n22833 = ~n22758 & n22831 ;
  assign n22834 = n22832 | n22833 ;
  assign n22835 = n4584 & n19916 ;
  assign n22836 = n4649 | n22835 ;
  assign n22837 = ( ~n20095 & n22835 ) | ( ~n20095 & n22836 ) | ( n22835 & n22836 ) ;
  assign n22838 = n4637 & n20091 ;
  assign n22839 = n22837 | n22838 ;
  assign n22840 = x23 & n22839 ;
  assign n22841 = n4591 & ~n20100 ;
  assign n22842 = ( ~x23 & n22839 ) | ( ~x23 & n22841 ) | ( n22839 & n22841 ) ;
  assign n22843 = x23 & ~n22841 ;
  assign n22844 = ( ~n22840 & n22842 ) | ( ~n22840 & n22843 ) | ( n22842 & n22843 ) ;
  assign n22845 = n4203 & ~n19893 ;
  assign n22846 = x26 & n22845 ;
  assign n22847 = n4215 & n19882 ;
  assign n22848 = n4200 & ~n19701 ;
  assign n22849 = n2083 & n19368 ;
  assign n22850 = n22848 | n22849 ;
  assign n22851 = n22847 | n22850 ;
  assign n22852 = x26 & ~n22851 ;
  assign n22853 = ( ~x26 & n22845 ) | ( ~x26 & n22851 ) | ( n22845 & n22851 ) ;
  assign n22854 = ( ~n22846 & n22852 ) | ( ~n22846 & n22853 ) | ( n22852 & n22853 ) ;
  assign n22855 = n3273 & ~n18258 ;
  assign n22856 = n3270 | n22855 ;
  assign n22857 = ( n18730 & n22855 ) | ( n18730 & n22856 ) | ( n22855 & n22856 ) ;
  assign n22858 = n390 | n22857 ;
  assign n22859 = ( n18735 & n22857 ) | ( n18735 & n22858 ) | ( n22857 & n22858 ) ;
  assign n22860 = n3274 & ~n18362 ;
  assign n22861 = n22859 | n22860 ;
  assign n22862 = n162 | n918 ;
  assign n22863 = n17929 | n22862 ;
  assign n22864 = n4105 | n22863 ;
  assign n22865 = n677 | n2534 ;
  assign n22866 = n21131 | n22865 ;
  assign n22867 = n22864 | n22866 ;
  assign n22868 = n6126 | n22867 ;
  assign n22869 = n1281 | n22868 ;
  assign n22870 = n244 | n14296 ;
  assign n22871 = n13194 | n22870 ;
  assign n22872 = n4474 & ~n22871 ;
  assign n22873 = ~n22869 & n22872 ;
  assign n22874 = ( n22792 & n22861 ) | ( n22792 & ~n22873 ) | ( n22861 & ~n22873 ) ;
  assign n22875 = ( n22792 & ~n22861 ) | ( n22792 & n22873 ) | ( ~n22861 & n22873 ) ;
  assign n22876 = ( ~n22792 & n22874 ) | ( ~n22792 & n22875 ) | ( n22874 & n22875 ) ;
  assign n22877 = ( ~n22801 & n22803 ) | ( ~n22801 & n22876 ) | ( n22803 & n22876 ) ;
  assign n22878 = ( n22801 & n22803 ) | ( n22801 & ~n22876 ) | ( n22803 & ~n22876 ) ;
  assign n22879 = ( ~n22803 & n22877 ) | ( ~n22803 & n22878 ) | ( n22877 & n22878 ) ;
  assign n22880 = n3501 & n19248 ;
  assign n22881 = x29 & n22880 ;
  assign n22882 = n3536 & n19177 ;
  assign n22883 = n4039 | n22882 ;
  assign n22884 = ( ~n19315 & n22882 ) | ( ~n19315 & n22883 ) | ( n22882 & n22883 ) ;
  assign n22885 = n3541 | n22884 ;
  assign n22886 = ( ~n19320 & n22884 ) | ( ~n19320 & n22885 ) | ( n22884 & n22885 ) ;
  assign n22887 = x29 & ~n22886 ;
  assign n22888 = ( ~x29 & n22880 ) | ( ~x29 & n22886 ) | ( n22880 & n22886 ) ;
  assign n22889 = ( ~n22881 & n22887 ) | ( ~n22881 & n22888 ) | ( n22887 & n22888 ) ;
  assign n22890 = ( n22854 & ~n22879 ) | ( n22854 & n22889 ) | ( ~n22879 & n22889 ) ;
  assign n22891 = ( n22854 & n22879 ) | ( n22854 & ~n22889 ) | ( n22879 & ~n22889 ) ;
  assign n22892 = ( ~n22854 & n22890 ) | ( ~n22854 & n22891 ) | ( n22890 & n22891 ) ;
  assign n22893 = ( n22806 & n22844 ) | ( n22806 & ~n22892 ) | ( n22844 & ~n22892 ) ;
  assign n22894 = ( ~n22806 & n22844 ) | ( ~n22806 & n22892 ) | ( n22844 & n22892 ) ;
  assign n22895 = ( ~n22844 & n22893 ) | ( ~n22844 & n22894 ) | ( n22893 & n22894 ) ;
  assign n22896 = ( x20 & ~n22821 ) | ( x20 & n22895 ) | ( ~n22821 & n22895 ) ;
  assign n22897 = ( x20 & n22821 ) | ( x20 & ~n22895 ) | ( n22821 & ~n22895 ) ;
  assign n22898 = ( ~x20 & n22896 ) | ( ~x20 & n22897 ) | ( n22896 & n22897 ) ;
  assign n22899 = ( ~n22827 & n22829 ) | ( ~n22827 & n22898 ) | ( n22829 & n22898 ) ;
  assign n22900 = ( n22827 & n22829 ) | ( n22827 & ~n22898 ) | ( n22829 & ~n22898 ) ;
  assign n22901 = ( ~n22829 & n22899 ) | ( ~n22829 & n22900 ) | ( n22899 & n22900 ) ;
  assign n22902 = n22832 & ~n22901 ;
  assign n22903 = ~n22832 & n22901 ;
  assign n22904 = n22902 | n22903 ;
  assign n22905 = n4215 & n19916 ;
  assign n22906 = n4200 & n19882 ;
  assign n22907 = n2083 & ~n19701 ;
  assign n22908 = n22906 | n22907 ;
  assign n22909 = n22905 | n22908 ;
  assign n22910 = x26 & n22909 ;
  assign n22911 = n4203 & n19920 ;
  assign n22912 = ( ~x26 & n22909 ) | ( ~x26 & n22911 ) | ( n22909 & n22911 ) ;
  assign n22913 = x26 & ~n22911 ;
  assign n22914 = ( ~n22910 & n22912 ) | ( ~n22910 & n22913 ) | ( n22912 & n22913 ) ;
  assign n22915 = n3541 & ~n19374 ;
  assign n22916 = x29 & n22915 ;
  assign n22917 = n3536 & n19248 ;
  assign n22918 = n4039 | n22917 ;
  assign n22919 = ( n19368 & n22917 ) | ( n19368 & n22918 ) | ( n22917 & n22918 ) ;
  assign n22920 = n3501 & ~n19315 ;
  assign n22921 = n22919 | n22920 ;
  assign n22922 = x29 & ~n22921 ;
  assign n22923 = ( ~x29 & n22915 ) | ( ~x29 & n22921 ) | ( n22915 & n22921 ) ;
  assign n22924 = ( ~n22916 & n22922 ) | ( ~n22916 & n22923 ) | ( n22922 & n22923 ) ;
  assign n22925 = n1289 | n2916 ;
  assign n22926 = n5078 | n22925 ;
  assign n22927 = n1401 | n2246 ;
  assign n22928 = n842 | n1711 ;
  assign n22929 = n22927 | n22928 ;
  assign n22930 = n13210 & ~n22929 ;
  assign n22931 = ~n22926 & n22930 ;
  assign n22932 = n335 | n1086 ;
  assign n22933 = n350 | n412 ;
  assign n22934 = n22932 | n22933 ;
  assign n22935 = n693 | n22934 ;
  assign n22936 = n22931 & ~n22935 ;
  assign n22937 = n1686 | n14847 ;
  assign n22938 = n22936 & ~n22937 ;
  assign n22939 = ~n4415 & n22938 ;
  assign n22940 = ( ~x20 & n22792 ) | ( ~x20 & n22939 ) | ( n22792 & n22939 ) ;
  assign n22941 = ( x20 & n22792 ) | ( x20 & n22939 ) | ( n22792 & n22939 ) ;
  assign n22942 = ( x20 & n22940 ) | ( x20 & ~n22941 ) | ( n22940 & ~n22941 ) ;
  assign n22943 = n3273 & ~n18362 ;
  assign n22944 = n3270 | n22943 ;
  assign n22945 = ( n19177 & n22943 ) | ( n19177 & n22944 ) | ( n22943 & n22944 ) ;
  assign n22946 = n390 | n22945 ;
  assign n22947 = ( ~n19182 & n22945 ) | ( ~n19182 & n22946 ) | ( n22945 & n22946 ) ;
  assign n22948 = n3274 & n18730 ;
  assign n22949 = n22947 | n22948 ;
  assign n22950 = ( n22874 & ~n22942 ) | ( n22874 & n22949 ) | ( ~n22942 & n22949 ) ;
  assign n22951 = ( n22874 & n22942 ) | ( n22874 & ~n22949 ) | ( n22942 & ~n22949 ) ;
  assign n22952 = ( ~n22874 & n22950 ) | ( ~n22874 & n22951 ) | ( n22950 & n22951 ) ;
  assign n22953 = ( n22878 & n22924 ) | ( n22878 & ~n22952 ) | ( n22924 & ~n22952 ) ;
  assign n22954 = ( ~n22878 & n22924 ) | ( ~n22878 & n22952 ) | ( n22924 & n22952 ) ;
  assign n22955 = ( ~n22924 & n22953 ) | ( ~n22924 & n22954 ) | ( n22953 & n22954 ) ;
  assign n22956 = ( n22890 & n22914 ) | ( n22890 & ~n22955 ) | ( n22914 & ~n22955 ) ;
  assign n22957 = ( n22890 & ~n22914 ) | ( n22890 & n22955 ) | ( ~n22914 & n22955 ) ;
  assign n22958 = ( ~n22890 & n22956 ) | ( ~n22890 & n22957 ) | ( n22956 & n22957 ) ;
  assign n22959 = n4637 & ~n20095 ;
  assign n22960 = n4584 & n20091 ;
  assign n22961 = n22959 | n22960 ;
  assign n22962 = x23 & n22961 ;
  assign n22963 = n4591 & ~n20097 ;
  assign n22964 = ( ~x23 & n22961 ) | ( ~x23 & n22963 ) | ( n22961 & n22963 ) ;
  assign n22965 = x23 & ~n22963 ;
  assign n22966 = ( ~n22962 & n22964 ) | ( ~n22962 & n22965 ) | ( n22964 & n22965 ) ;
  assign n22967 = ( n22893 & n22958 ) | ( n22893 & n22966 ) | ( n22958 & n22966 ) ;
  assign n22968 = ( n22893 & ~n22958 ) | ( n22893 & n22966 ) | ( ~n22958 & n22966 ) ;
  assign n22969 = ( n22958 & ~n22967 ) | ( n22958 & n22968 ) | ( ~n22967 & n22968 ) ;
  assign n22970 = ( ~n22897 & n22900 ) | ( ~n22897 & n22969 ) | ( n22900 & n22969 ) ;
  assign n22971 = ( n22897 & n22900 ) | ( n22897 & ~n22969 ) | ( n22900 & ~n22969 ) ;
  assign n22972 = ( ~n22900 & n22970 ) | ( ~n22900 & n22971 ) | ( n22970 & n22971 ) ;
  assign n22973 = n22902 & ~n22972 ;
  assign n22974 = ~n22902 & n22972 ;
  assign n22975 = n22973 | n22974 ;
  assign n22976 = n4579 & ~n20095 ;
  assign n22977 = n4583 | n20095 ;
  assign n22978 = ( x23 & n22976 ) | ( x23 & n22977 ) | ( n22976 & n22977 ) ;
  assign n22979 = n2083 & n19882 ;
  assign n22980 = x26 & n22979 ;
  assign n22981 = n4215 & n20091 ;
  assign n22982 = n4200 & n19916 ;
  assign n22983 = n22981 | n22982 ;
  assign n22984 = n4203 | n22983 ;
  assign n22985 = ( n20101 & n22983 ) | ( n20101 & n22984 ) | ( n22983 & n22984 ) ;
  assign n22986 = x26 & ~n22985 ;
  assign n22987 = ( ~x26 & n22979 ) | ( ~x26 & n22985 ) | ( n22979 & n22985 ) ;
  assign n22988 = ( ~n22980 & n22986 ) | ( ~n22980 & n22987 ) | ( n22986 & n22987 ) ;
  assign n22989 = n3536 & ~n19315 ;
  assign n22990 = n4039 | n22989 ;
  assign n22991 = ( ~n19701 & n22989 ) | ( ~n19701 & n22990 ) | ( n22989 & n22990 ) ;
  assign n22992 = n3501 & n19368 ;
  assign n22993 = n22991 | n22992 ;
  assign n22994 = x29 & n22993 ;
  assign n22995 = n3541 & ~n19706 ;
  assign n22996 = x29 & ~n22995 ;
  assign n22997 = ( ~x29 & n22993 ) | ( ~x29 & n22995 ) | ( n22993 & n22995 ) ;
  assign n22998 = ( ~n22994 & n22996 ) | ( ~n22994 & n22997 ) | ( n22996 & n22997 ) ;
  assign n22999 = n3273 & n18730 ;
  assign n23000 = n3270 | n22999 ;
  assign n23001 = ( n19248 & n22999 ) | ( n19248 & n23000 ) | ( n22999 & n23000 ) ;
  assign n23002 = n390 | n23001 ;
  assign n23003 = ( n19253 & n23001 ) | ( n19253 & n23002 ) | ( n23001 & n23002 ) ;
  assign n23004 = n3274 & n19177 ;
  assign n23005 = n23003 | n23004 ;
  assign n23006 = n314 | n2269 ;
  assign n23007 = n4781 | n23006 ;
  assign n23008 = n2122 | n23007 ;
  assign n23009 = n4012 | n23008 ;
  assign n23010 = n928 | n1843 ;
  assign n23011 = n2156 | n23010 ;
  assign n23012 = n279 | n915 ;
  assign n23013 = n5031 | n23012 ;
  assign n23014 = n23011 | n23013 ;
  assign n23015 = n23009 | n23014 ;
  assign n23016 = n12681 | n15507 ;
  assign n23017 = n2200 | n23016 ;
  assign n23018 = n23015 | n23017 ;
  assign n23019 = n4115 | n23018 ;
  assign n23020 = ( n22941 & n23005 ) | ( n22941 & n23019 ) | ( n23005 & n23019 ) ;
  assign n23021 = ( n22941 & ~n23005 ) | ( n22941 & n23019 ) | ( ~n23005 & n23019 ) ;
  assign n23022 = ( n23005 & ~n23020 ) | ( n23005 & n23021 ) | ( ~n23020 & n23021 ) ;
  assign n23023 = ( n22950 & n22998 ) | ( n22950 & n23022 ) | ( n22998 & n23022 ) ;
  assign n23024 = ( n22950 & ~n22998 ) | ( n22950 & n23022 ) | ( ~n22998 & n23022 ) ;
  assign n23025 = ( n22998 & ~n23023 ) | ( n22998 & n23024 ) | ( ~n23023 & n23024 ) ;
  assign n23026 = ( n22953 & ~n22988 ) | ( n22953 & n23025 ) | ( ~n22988 & n23025 ) ;
  assign n23027 = ( n22953 & n22988 ) | ( n22953 & n23025 ) | ( n22988 & n23025 ) ;
  assign n23028 = ( n22988 & n23026 ) | ( n22988 & ~n23027 ) | ( n23026 & ~n23027 ) ;
  assign n23029 = ( ~n22956 & n22978 ) | ( ~n22956 & n23028 ) | ( n22978 & n23028 ) ;
  assign n23030 = ( n22956 & n22978 ) | ( n22956 & n23028 ) | ( n22978 & n23028 ) ;
  assign n23031 = ( n22956 & n23029 ) | ( n22956 & ~n23030 ) | ( n23029 & ~n23030 ) ;
  assign n23032 = ( n22968 & ~n22971 ) | ( n22968 & n23031 ) | ( ~n22971 & n23031 ) ;
  assign n23033 = ( n22968 & n22971 ) | ( n22968 & n23031 ) | ( n22971 & n23031 ) ;
  assign n23034 = ( n22971 & n23032 ) | ( n22971 & ~n23033 ) | ( n23032 & ~n23033 ) ;
  assign n23035 = n22973 & ~n23034 ;
  assign n23036 = n22973 & n23034 ;
  assign n23037 = ( n23034 & n23035 ) | ( n23034 & ~n23036 ) | ( n23035 & ~n23036 ) ;
  assign n23038 = n2083 & n19916 ;
  assign n23039 = x26 & n23038 ;
  assign n23040 = n4215 & ~n20095 ;
  assign n23041 = n4200 & n20091 ;
  assign n23042 = n23040 | n23041 ;
  assign n23043 = n4203 & ~n20100 ;
  assign n23044 = n23042 | n23043 ;
  assign n23045 = x26 & ~n23044 ;
  assign n23046 = ( ~x26 & n23038 ) | ( ~x26 & n23044 ) | ( n23038 & n23044 ) ;
  assign n23047 = ( ~n23039 & n23045 ) | ( ~n23039 & n23046 ) | ( n23045 & n23046 ) ;
  assign n23048 = n3501 & ~n19701 ;
  assign n23049 = x29 & n23048 ;
  assign n23050 = n3536 & n19368 ;
  assign n23051 = n4039 | n23050 ;
  assign n23052 = ( n19882 & n23050 ) | ( n19882 & n23051 ) | ( n23050 & n23051 ) ;
  assign n23053 = n3541 | n23052 ;
  assign n23054 = ( ~n19893 & n23052 ) | ( ~n19893 & n23053 ) | ( n23052 & n23053 ) ;
  assign n23055 = x29 & ~n23054 ;
  assign n23056 = ( ~x29 & n23048 ) | ( ~x29 & n23054 ) | ( n23048 & n23054 ) ;
  assign n23057 = ( ~n23049 & n23055 ) | ( ~n23049 & n23056 ) | ( n23055 & n23056 ) ;
  assign n23058 = n3484 | n18695 ;
  assign n23059 = n1843 | n13590 ;
  assign n23060 = n23058 | n23059 ;
  assign n23061 = n21711 | n23060 ;
  assign n23062 = n330 | n342 ;
  assign n23063 = n1184 | n23062 ;
  assign n23064 = n290 | n939 ;
  assign n23065 = n23063 | n23064 ;
  assign n23066 = n917 | n3327 ;
  assign n23067 = n23065 | n23066 ;
  assign n23068 = n19288 | n23067 ;
  assign n23069 = n23061 | n23068 ;
  assign n23070 = n18497 & ~n23069 ;
  assign n23071 = ~n3629 & n23070 ;
  assign n23072 = ( n23019 & n23021 ) | ( n23019 & ~n23071 ) | ( n23021 & ~n23071 ) ;
  assign n23073 = ( ~n22941 & n23020 ) | ( ~n22941 & n23071 ) | ( n23020 & n23071 ) ;
  assign n23074 = ( ~n23019 & n23072 ) | ( ~n23019 & n23073 ) | ( n23072 & n23073 ) ;
  assign n23075 = n3273 & n19177 ;
  assign n23076 = n3270 | n23075 ;
  assign n23077 = ( ~n19315 & n23075 ) | ( ~n19315 & n23076 ) | ( n23075 & n23076 ) ;
  assign n23078 = n390 | n23077 ;
  assign n23079 = ( ~n19320 & n23077 ) | ( ~n19320 & n23078 ) | ( n23077 & n23078 ) ;
  assign n23080 = n3274 & n19248 ;
  assign n23081 = n23079 | n23080 ;
  assign n23082 = ( n23023 & n23074 ) | ( n23023 & n23081 ) | ( n23074 & n23081 ) ;
  assign n23083 = ( n23023 & ~n23074 ) | ( n23023 & n23081 ) | ( ~n23074 & n23081 ) ;
  assign n23084 = ( n23074 & ~n23082 ) | ( n23074 & n23083 ) | ( ~n23082 & n23083 ) ;
  assign n23085 = ( n23047 & ~n23057 ) | ( n23047 & n23084 ) | ( ~n23057 & n23084 ) ;
  assign n23086 = ( n23047 & n23057 ) | ( n23047 & ~n23084 ) | ( n23057 & ~n23084 ) ;
  assign n23087 = ( ~n23047 & n23085 ) | ( ~n23047 & n23086 ) | ( n23085 & n23086 ) ;
  assign n23088 = ( ~x23 & n23027 ) | ( ~x23 & n23087 ) | ( n23027 & n23087 ) ;
  assign n23089 = ( x23 & n23027 ) | ( x23 & ~n23087 ) | ( n23027 & ~n23087 ) ;
  assign n23090 = ( ~n23027 & n23088 ) | ( ~n23027 & n23089 ) | ( n23088 & n23089 ) ;
  assign n23091 = ( n23030 & n23033 ) | ( n23030 & ~n23090 ) | ( n23033 & ~n23090 ) ;
  assign n23092 = ( ~n23030 & n23033 ) | ( ~n23030 & n23090 ) | ( n23033 & n23090 ) ;
  assign n23093 = ( ~n23033 & n23091 ) | ( ~n23033 & n23092 ) | ( n23091 & n23092 ) ;
  assign n23094 = n23036 & ~n23093 ;
  assign n23095 = ~n23036 & n23093 ;
  assign n23096 = n23094 | n23095 ;
  assign n23097 = n4200 & ~n20095 ;
  assign n23098 = n2083 & n20091 ;
  assign n23099 = n23097 | n23098 ;
  assign n23100 = x26 & n23099 ;
  assign n23101 = n4203 & ~n20097 ;
  assign n23102 = ( ~x26 & n23099 ) | ( ~x26 & n23101 ) | ( n23099 & n23101 ) ;
  assign n23103 = x26 & ~n23101 ;
  assign n23104 = ( ~n23100 & n23102 ) | ( ~n23100 & n23103 ) | ( n23102 & n23103 ) ;
  assign n23105 = n3541 & n19920 ;
  assign n23106 = x29 & n23105 ;
  assign n23107 = n3536 & ~n19701 ;
  assign n23108 = n4039 | n23107 ;
  assign n23109 = ( n19916 & n23107 ) | ( n19916 & n23108 ) | ( n23107 & n23108 ) ;
  assign n23110 = n3501 & n19882 ;
  assign n23111 = n23109 | n23110 ;
  assign n23112 = x29 & ~n23111 ;
  assign n23113 = ( ~x29 & n23105 ) | ( ~x29 & n23111 ) | ( n23105 & n23111 ) ;
  assign n23114 = ( ~n23106 & n23112 ) | ( ~n23106 & n23113 ) | ( n23112 & n23113 ) ;
  assign n23115 = n3273 & n19248 ;
  assign n23116 = n3270 | n23115 ;
  assign n23117 = ( n19368 & n23115 ) | ( n19368 & n23116 ) | ( n23115 & n23116 ) ;
  assign n23118 = n390 | n23117 ;
  assign n23119 = ( ~n19374 & n23117 ) | ( ~n19374 & n23118 ) | ( n23117 & n23118 ) ;
  assign n23120 = n3274 & ~n19315 ;
  assign n23121 = n23119 | n23120 ;
  assign n23122 = n44 | n794 ;
  assign n23123 = n131 | n712 ;
  assign n23124 = n23122 | n23123 ;
  assign n23125 = n237 | n1107 ;
  assign n23126 = n23124 | n23125 ;
  assign n23127 = n4789 | n23126 ;
  assign n23128 = n13617 | n23127 ;
  assign n23129 = n1724 | n2084 ;
  assign n23130 = n4916 | n23129 ;
  assign n23131 = n23128 | n23130 ;
  assign n23132 = n3567 & ~n23131 ;
  assign n23133 = ~n10204 & n23132 ;
  assign n23134 = ( ~x23 & n23071 ) | ( ~x23 & n23133 ) | ( n23071 & n23133 ) ;
  assign n23135 = ( x23 & n23071 ) | ( x23 & n23133 ) | ( n23071 & n23133 ) ;
  assign n23136 = ( x23 & n23134 ) | ( x23 & ~n23135 ) | ( n23134 & ~n23135 ) ;
  assign n23137 = ( ~n23073 & n23121 ) | ( ~n23073 & n23136 ) | ( n23121 & n23136 ) ;
  assign n23138 = ( n23073 & n23121 ) | ( n23073 & ~n23136 ) | ( n23121 & ~n23136 ) ;
  assign n23139 = ( ~n23121 & n23137 ) | ( ~n23121 & n23138 ) | ( n23137 & n23138 ) ;
  assign n23140 = ( n23083 & n23114 ) | ( n23083 & ~n23139 ) | ( n23114 & ~n23139 ) ;
  assign n23141 = ( n23083 & ~n23114 ) | ( n23083 & n23139 ) | ( ~n23114 & n23139 ) ;
  assign n23142 = ( ~n23083 & n23140 ) | ( ~n23083 & n23141 ) | ( n23140 & n23141 ) ;
  assign n23143 = ( n23086 & n23104 ) | ( n23086 & ~n23142 ) | ( n23104 & ~n23142 ) ;
  assign n23144 = ( n23086 & ~n23104 ) | ( n23086 & n23142 ) | ( ~n23104 & n23142 ) ;
  assign n23145 = ( ~n23086 & n23143 ) | ( ~n23086 & n23144 ) | ( n23143 & n23144 ) ;
  assign n23146 = n23089 & ~n23145 ;
  assign n23147 = ~n23089 & n23145 ;
  assign n23148 = n23146 | n23147 ;
  assign n23149 = ( n23091 & ~n23094 ) | ( n23091 & n23148 ) | ( ~n23094 & n23148 ) ;
  assign n23150 = ( n23091 & n23094 ) | ( n23091 & ~n23148 ) | ( n23094 & ~n23148 ) ;
  assign n23151 = ( ~n23091 & n23149 ) | ( ~n23091 & n23150 ) | ( n23149 & n23150 ) ;
  assign n23152 = n23091 | n23146 ;
  assign n23153 = ( n23094 & ~n23147 ) | ( n23094 & n23152 ) | ( ~n23147 & n23152 ) ;
  assign n23154 = n23091 & n23146 ;
  assign n23155 = n23094 & n23154 ;
  assign n23156 = n23153 & ~n23155 ;
  assign n23157 = n3536 & n19882 ;
  assign n23158 = x29 & n23157 ;
  assign n23159 = n4039 & n20091 ;
  assign n23160 = n3541 | n23159 ;
  assign n23161 = ( n20101 & n23159 ) | ( n20101 & n23160 ) | ( n23159 & n23160 ) ;
  assign n23162 = n3501 & n19916 ;
  assign n23163 = n23161 | n23162 ;
  assign n23164 = x29 & ~n23163 ;
  assign n23165 = ( ~x29 & n23157 ) | ( ~x29 & n23163 ) | ( n23157 & n23163 ) ;
  assign n23166 = ( ~n23158 & n23164 ) | ( ~n23158 & n23165 ) | ( n23164 & n23165 ) ;
  assign n23167 = n91 | n15764 ;
  assign n23168 = n6085 | n23167 ;
  assign n23169 = n3470 | n23168 ;
  assign n23170 = n3557 | n4101 ;
  assign n23171 = n150 | n264 ;
  assign n23172 = n3116 | n23171 ;
  assign n23173 = n572 | n23172 ;
  assign n23174 = n23170 | n23173 ;
  assign n23175 = n329 | n674 ;
  assign n23176 = n351 | n23175 ;
  assign n23177 = n844 | n12844 ;
  assign n23178 = n23176 | n23177 ;
  assign n23179 = n3413 | n23178 ;
  assign n23180 = n23174 | n23179 ;
  assign n23181 = n23169 | n23180 ;
  assign n23182 = n13628 | n23181 ;
  assign n23183 = n3273 & ~n19315 ;
  assign n23184 = n3270 | n23183 ;
  assign n23185 = ( ~n19701 & n23183 ) | ( ~n19701 & n23184 ) | ( n23183 & n23184 ) ;
  assign n23186 = n390 | n23185 ;
  assign n23187 = ( ~n19706 & n23185 ) | ( ~n19706 & n23186 ) | ( n23185 & n23186 ) ;
  assign n23188 = n3274 & n19368 ;
  assign n23189 = n23187 | n23188 ;
  assign n23190 = ( ~n23135 & n23182 ) | ( ~n23135 & n23189 ) | ( n23182 & n23189 ) ;
  assign n23191 = ( n23135 & n23182 ) | ( n23135 & ~n23189 ) | ( n23182 & ~n23189 ) ;
  assign n23192 = ( ~n23182 & n23190 ) | ( ~n23182 & n23191 ) | ( n23190 & n23191 ) ;
  assign n23193 = ( n23138 & n23166 ) | ( n23138 & n23192 ) | ( n23166 & n23192 ) ;
  assign n23194 = ( n23138 & ~n23166 ) | ( n23138 & n23192 ) | ( ~n23166 & n23192 ) ;
  assign n23195 = ( n23166 & ~n23193 ) | ( n23166 & n23194 ) | ( ~n23193 & n23194 ) ;
  assign n23196 = x26 & n13475 ;
  assign n23197 = n19266 | n23196 ;
  assign n23198 = ( n23140 & ~n23195 ) | ( n23140 & n23197 ) | ( ~n23195 & n23197 ) ;
  assign n23199 = ( n23140 & n23195 ) | ( n23140 & n23197 ) | ( n23195 & n23197 ) ;
  assign n23200 = ( n23195 & n23198 ) | ( n23195 & ~n23199 ) | ( n23198 & ~n23199 ) ;
  assign n23201 = ( ~n23143 & n23156 ) | ( ~n23143 & n23200 ) | ( n23156 & n23200 ) ;
  assign n23202 = ( n23143 & n23156 ) | ( n23143 & ~n23200 ) | ( n23156 & ~n23200 ) ;
  assign n23203 = ( ~n23156 & n23201 ) | ( ~n23156 & n23202 ) | ( n23201 & n23202 ) ;
  assign n23204 = n23143 & n23200 ;
  assign n23205 = n23155 & n23204 ;
  assign n23206 = n23143 | n23200 ;
  assign n23207 = n23155 | n23206 ;
  assign n23208 = n23153 & ~n23204 ;
  assign n23209 = ~n23155 & n23204 ;
  assign n23210 = ( n23207 & n23208 ) | ( n23207 & n23209 ) | ( n23208 & n23209 ) ;
  assign n23211 = n3273 & n19368 ;
  assign n23212 = n3270 | n23211 ;
  assign n23213 = ( n19882 & n23211 ) | ( n19882 & n23212 ) | ( n23211 & n23212 ) ;
  assign n23214 = n390 | n23213 ;
  assign n23215 = ( ~n19893 & n23213 ) | ( ~n19893 & n23214 ) | ( n23213 & n23214 ) ;
  assign n23216 = n3274 & ~n19701 ;
  assign n23217 = n23215 | n23216 ;
  assign n23218 = n3413 | n3424 ;
  assign n23219 = ~n1048 & n3503 ;
  assign n23220 = ~n803 & n23219 ;
  assign n23221 = ~n23218 & n23220 ;
  assign n23222 = ~n3579 & n23221 ;
  assign n23223 = ~n3589 & n23222 ;
  assign n23224 = ~n3526 & n23223 ;
  assign n23225 = ( ~n23182 & n23191 ) | ( ~n23182 & n23224 ) | ( n23191 & n23224 ) ;
  assign n23226 = ( n23182 & n23191 ) | ( n23182 & n23224 ) | ( n23191 & n23224 ) ;
  assign n23227 = ( n23182 & n23225 ) | ( n23182 & ~n23226 ) | ( n23225 & ~n23226 ) ;
  assign n23228 = ( n23193 & n23217 ) | ( n23193 & ~n23227 ) | ( n23217 & ~n23227 ) ;
  assign n23229 = ( n23193 & ~n23217 ) | ( n23193 & n23227 ) | ( ~n23217 & n23227 ) ;
  assign n23230 = ( ~n23193 & n23228 ) | ( ~n23193 & n23229 ) | ( n23228 & n23229 ) ;
  assign n23231 = n3541 & ~n20100 ;
  assign n23232 = n4039 & ~n20095 ;
  assign n23233 = n3501 & n20091 ;
  assign n23234 = n23232 | n23233 ;
  assign n23235 = n23231 | n23234 ;
  assign n23236 = n3536 & n19916 ;
  assign n23237 = n23235 | n23236 ;
  assign n23238 = ( n6269 & ~n23235 ) | ( n6269 & n23237 ) | ( ~n23235 & n23237 ) ;
  assign n23239 = ( ~n23230 & n23237 ) | ( ~n23230 & n23238 ) | ( n23237 & n23238 ) ;
  assign n23240 = ( n23230 & n23237 ) | ( n23230 & n23238 ) | ( n23237 & n23238 ) ;
  assign n23241 = ( n23230 & n23239 ) | ( n23230 & ~n23240 ) | ( n23239 & ~n23240 ) ;
  assign n23242 = ~n23199 & n23241 ;
  assign n23243 = n23199 & ~n23241 ;
  assign n23244 = n23242 | n23243 ;
  assign n23245 = ~n23210 & n23244 ;
  assign n23246 = ~n23205 & n23244 ;
  assign n23247 = ( n23205 & n23210 ) | ( n23205 & ~n23246 ) | ( n23210 & ~n23246 ) ;
  assign n23248 = ( ~n23205 & n23245 ) | ( ~n23205 & n23247 ) | ( n23245 & n23247 ) ;
  assign n23249 = x29 & ~n23237 ;
  assign n23250 = ~x29 & n23237 ;
  assign n23251 = n23249 | n23250 ;
  assign n23252 = ( x26 & ~n23230 ) | ( x26 & n23251 ) | ( ~n23230 & n23251 ) ;
  assign n23253 = n3536 & n20091 ;
  assign n23254 = n3541 | n23253 ;
  assign n23255 = ( ~n20097 & n23253 ) | ( ~n20097 & n23254 ) | ( n23253 & n23254 ) ;
  assign n23256 = n3273 & ~n19701 ;
  assign n23257 = n3270 | n23256 ;
  assign n23258 = ( n19916 & n23256 ) | ( n19916 & n23257 ) | ( n23256 & n23257 ) ;
  assign n23259 = n390 | n23258 ;
  assign n23260 = ( n19920 & n23258 ) | ( n19920 & n23259 ) | ( n23258 & n23259 ) ;
  assign n23261 = n3274 & n19882 ;
  assign n23262 = n23260 | n23261 ;
  assign n23263 = n3514 | n3530 ;
  assign n23264 = ( n6269 & n23182 ) | ( n6269 & n23263 ) | ( n23182 & n23263 ) ;
  assign n23265 = ( ~n6269 & n23182 ) | ( ~n6269 & n23263 ) | ( n23182 & n23263 ) ;
  assign n23266 = ( n6269 & ~n23264 ) | ( n6269 & n23265 ) | ( ~n23264 & n23265 ) ;
  assign n23267 = n23226 | n23266 ;
  assign n23268 = n23226 & n23266 ;
  assign n23269 = n23267 & ~n23268 ;
  assign n23270 = ( n23255 & ~n23262 ) | ( n23255 & n23269 ) | ( ~n23262 & n23269 ) ;
  assign n23271 = ( n23255 & n23262 ) | ( n23255 & ~n23269 ) | ( n23262 & ~n23269 ) ;
  assign n23272 = ( ~n23255 & n23270 ) | ( ~n23255 & n23271 ) | ( n23270 & n23271 ) ;
  assign n23273 = ( ~n23228 & n23252 ) | ( ~n23228 & n23272 ) | ( n23252 & n23272 ) ;
  assign n23274 = ( n23228 & n23252 ) | ( n23228 & n23272 ) | ( n23252 & n23272 ) ;
  assign n23275 = ( n23228 & n23273 ) | ( n23228 & ~n23274 ) | ( n23273 & ~n23274 ) ;
  assign n23276 = ( n23243 & ~n23247 ) | ( n23243 & n23275 ) | ( ~n23247 & n23275 ) ;
  assign n23277 = ( n23243 & n23247 ) | ( n23243 & ~n23275 ) | ( n23247 & ~n23275 ) ;
  assign n23278 = ( ~n23243 & n23276 ) | ( ~n23243 & n23277 ) | ( n23276 & n23277 ) ;
  assign y0 = n19903 ;
  assign y1 = n20080 ;
  assign y2 = ~n20257 ;
  assign y3 = ~n20416 ;
  assign y4 = ~n20579 ;
  assign y5 = ~n20728 ;
  assign y6 = ~n20885 ;
  assign y7 = ~n21039 ;
  assign y8 = n21187 ;
  assign y9 = n21331 ;
  assign y10 = n21473 ;
  assign y11 = n21615 ;
  assign y12 = ~n21755 ;
  assign y13 = ~n21876 ;
  assign y14 = ~n21992 ;
  assign y15 = n22105 ;
  assign y16 = ~n22215 ;
  assign y17 = n22315 ;
  assign y18 = ~n22412 ;
  assign y19 = ~n22505 ;
  assign y20 = ~n22594 ;
  assign y21 = n22679 ;
  assign y22 = n22759 ;
  assign y23 = ~n22834 ;
  assign y24 = ~n22904 ;
  assign y25 = ~n22975 ;
  assign y26 = n23037 ;
  assign y27 = ~n23096 ;
  assign y28 = ~n23151 ;
  assign y29 = n23203 ;
  assign y30 = ~n23248 ;
  assign y31 = n23278 ;
endmodule
