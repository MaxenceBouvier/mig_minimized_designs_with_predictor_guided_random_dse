module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 ;
  assign n25 = x0 | x1 ;
  assign n26 = x2 | n25 ;
  assign n27 = x3 | n26 ;
  assign n28 = x4 | n27 ;
  assign n29 = x5 | n28 ;
  assign n30 = x6 | n29 ;
  assign n31 = x7 | n30 ;
  assign n32 = x8 | n31 ;
  assign n33 = x9 | n32 ;
  assign n34 = x10 | n33 ;
  assign n35 = x11 | n34 ;
  assign n36 = x12 | n35 ;
  assign n37 = x13 | n36 ;
  assign n38 = x14 | n37 ;
  assign n39 = x15 | n38 ;
  assign n40 = ( x15 & x22 ) | ( x15 & ~n38 ) | ( x22 & ~n38 ) ;
  assign n41 = x15 | x22 ;
  assign n42 = ( n39 & n40 ) | ( n39 & ~n41 ) | ( n40 & ~n41 ) ;
  assign n43 = x18 | x19 ;
  assign n44 = x15 & ~x22 ;
  assign n45 = ( ~x22 & n38 ) | ( ~x22 & n44 ) | ( n38 & n44 ) ;
  assign n46 = x16 | n45 ;
  assign n47 = x17 | n46 ;
  assign n48 = ~x22 & n47 ;
  assign n49 = ( ~x22 & n43 ) | ( ~x22 & n48 ) | ( n43 & n48 ) ;
  assign n50 = x20 | n49 ;
  assign n51 = x20 & n49 ;
  assign n52 = n50 & ~n51 ;
  assign n53 = x21 & x22 ;
  assign n54 = x21 | x22 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = n52 & n55 ;
  assign n57 = ~n42 & n56 ;
  assign n58 = x16 & n45 ;
  assign n59 = n46 & ~n58 ;
  assign n60 = x17 & x22 ;
  assign n61 = x17 | x22 ;
  assign n62 = ~n60 & n61 ;
  assign n63 = n59 & ~n62 ;
  assign n64 = ~x18 & x19 ;
  assign n65 = x19 & n48 ;
  assign n66 = x18 & n48 ;
  assign n67 = ( n64 & ~n65 ) | ( n64 & n66 ) | ( ~n65 & n66 ) ;
  assign n68 = n63 & n67 ;
  assign n69 = n56 & n68 ;
  assign n70 = ~n57 & n69 ;
  assign n71 = x19 & x22 ;
  assign n72 = x18 & x22 ;
  assign n73 = ( n64 & ~n71 ) | ( n64 & n72 ) | ( ~n71 & n72 ) ;
  assign n74 = n63 & n73 ;
  assign n75 = x21 & ~n50 ;
  assign n76 = ~x21 & n51 ;
  assign n77 = n75 | n76 ;
  assign n78 = n52 | n77 ;
  assign n79 = n42 | n78 ;
  assign n80 = n74 & ~n79 ;
  assign n81 = n42 & ~n78 ;
  assign n82 = n43 | n48 ;
  assign n83 = x18 & x19 ;
  assign n84 = n48 & n83 ;
  assign n85 = n82 & ~n84 ;
  assign n86 = n63 & ~n85 ;
  assign n87 = n81 & n86 ;
  assign n88 = n80 | n87 ;
  assign n89 = n70 | n88 ;
  assign n90 = n59 & n62 ;
  assign n91 = n67 & n90 ;
  assign n92 = n57 & n91 ;
  assign n93 = x17 & n58 ;
  assign n94 = n47 & ~n93 ;
  assign n95 = n85 | n94 ;
  assign n96 = n57 & ~n95 ;
  assign n97 = x19 | x22 ;
  assign n98 = ~n71 & n97 ;
  assign n99 = n72 | n83 ;
  assign n100 = ( n43 & n98 ) | ( n43 & ~n99 ) | ( n98 & ~n99 ) ;
  assign n101 = n90 & ~n100 ;
  assign n102 = n81 & n101 ;
  assign n103 = n96 | n102 ;
  assign n104 = n92 | n103 ;
  assign n105 = n89 | n104 ;
  assign n106 = n52 & ~n55 ;
  assign n107 = ~n42 & n106 ;
  assign n108 = n101 & n107 ;
  assign n109 = n42 & n77 ;
  assign n110 = ~n59 & n94 ;
  assign n111 = n73 & n110 ;
  assign n112 = n109 & n111 ;
  assign n113 = ~n42 & n77 ;
  assign n114 = n74 & n113 ;
  assign n115 = n112 | n114 ;
  assign n116 = n108 | n115 ;
  assign n117 = n42 & n56 ;
  assign n118 = ~n95 & n117 ;
  assign n119 = n91 & n109 ;
  assign n120 = n118 | n119 ;
  assign n121 = n68 & ~n79 ;
  assign n122 = ~n42 & n52 ;
  assign n123 = n74 & n122 ;
  assign n124 = n121 | n123 ;
  assign n125 = n120 | n124 ;
  assign n126 = n42 & n106 ;
  assign n127 = n68 & n126 ;
  assign n128 = n67 & n110 ;
  assign n129 = n57 & n128 ;
  assign n130 = n86 & n117 ;
  assign n131 = n129 | n130 ;
  assign n132 = n127 | n131 ;
  assign n133 = n125 | n132 ;
  assign n134 = n116 | n133 ;
  assign n135 = n105 | n134 ;
  assign n136 = n107 & n111 ;
  assign n137 = n91 & n107 ;
  assign n138 = n136 | n137 ;
  assign n139 = n63 & ~n100 ;
  assign n140 = n113 & n139 ;
  assign n141 = n74 & n109 ;
  assign n142 = n140 | n141 ;
  assign n143 = n138 | n142 ;
  assign n144 = ~n100 & n110 ;
  assign n145 = n81 & n144 ;
  assign n146 = n117 & n128 ;
  assign n147 = n145 | n146 ;
  assign n148 = ~n85 & n110 ;
  assign n149 = ~n79 & n148 ;
  assign n150 = n101 & n113 ;
  assign n151 = n149 | n150 ;
  assign n152 = n147 | n151 ;
  assign n153 = n143 | n152 ;
  assign n154 = n77 & n86 ;
  assign n155 = x18 & ~n47 ;
  assign n156 = ~x18 & n93 ;
  assign n157 = n155 | n156 ;
  assign n158 = ~n98 & n157 ;
  assign n159 = n113 & n158 ;
  assign n160 = n154 | n159 ;
  assign n161 = n101 & n117 ;
  assign n162 = n68 & n81 ;
  assign n163 = n161 | n162 ;
  assign n164 = n126 & n148 ;
  assign n165 = n113 & n148 ;
  assign n166 = n164 | n165 ;
  assign n167 = n163 | n166 ;
  assign n168 = n160 | n167 ;
  assign n169 = n153 | n168 ;
  assign n170 = ~n95 & n107 ;
  assign n171 = n86 & n126 ;
  assign n172 = n170 | n171 ;
  assign n173 = n68 & n113 ;
  assign n174 = n67 & ~n94 ;
  assign n175 = ~n79 & n174 ;
  assign n176 = n74 & n117 ;
  assign n177 = n175 | n176 ;
  assign n178 = n173 | n177 ;
  assign n179 = n81 & n158 ;
  assign n180 = n107 & n128 ;
  assign n181 = n111 & n117 ;
  assign n182 = n180 | n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = n178 | n183 ;
  assign n185 = n172 | n184 ;
  assign n186 = n169 | n185 ;
  assign n187 = n135 | n186 ;
  assign n188 = n117 & n144 ;
  assign n189 = n73 & n90 ;
  assign n190 = n57 & n189 ;
  assign n191 = n188 | n190 ;
  assign n192 = ~n85 & n90 ;
  assign n193 = ~n79 & n192 ;
  assign n194 = n191 | n193 ;
  assign n195 = n81 & n189 ;
  assign n196 = n109 & n148 ;
  assign n197 = n195 | n196 ;
  assign n198 = ~n79 & n86 ;
  assign n199 = n109 & n192 ;
  assign n200 = n198 | n199 ;
  assign n201 = n197 | n200 ;
  assign n202 = n194 | n201 ;
  assign n203 = n57 & n192 ;
  assign n204 = n86 | n174 ;
  assign n205 = n107 & n204 ;
  assign n206 = n203 | n205 ;
  assign n207 = n106 & n158 ;
  assign n208 = n42 & n207 ;
  assign n209 = n109 & n174 ;
  assign n210 = n208 | n209 ;
  assign n211 = n206 | n210 ;
  assign n212 = n74 & n126 ;
  assign n213 = n126 & n144 ;
  assign n214 = ~n79 & n128 ;
  assign n215 = n213 | n214 ;
  assign n216 = n212 | n215 ;
  assign n217 = n211 | n216 ;
  assign n218 = n202 | n217 ;
  assign n219 = n187 | n218 ;
  assign n220 = ( x5 & x22 ) | ( x5 & ~n28 ) | ( x22 & ~n28 ) ;
  assign n221 = x5 | x22 ;
  assign n222 = ( n29 & n220 ) | ( n29 & ~n221 ) | ( n220 & ~n221 ) ;
  assign n223 = ( x4 & x22 ) | ( x4 & ~n27 ) | ( x22 & ~n27 ) ;
  assign n224 = x4 | x22 ;
  assign n225 = ( n28 & n223 ) | ( n28 & ~n224 ) | ( n223 & ~n224 ) ;
  assign n226 = n222 & n225 ;
  assign n227 = n222 | n225 ;
  assign n228 = ~n226 & n227 ;
  assign n229 = ( x2 & x22 ) | ( x2 & ~n25 ) | ( x22 & ~n25 ) ;
  assign n230 = x2 | x22 ;
  assign n231 = ( n26 & n229 ) | ( n26 & ~n230 ) | ( n229 & ~n230 ) ;
  assign n232 = ( x3 & x22 ) | ( x3 & ~n26 ) | ( x22 & ~n26 ) ;
  assign n233 = x3 | x22 ;
  assign n234 = ( n27 & n232 ) | ( n27 & ~n233 ) | ( n232 & ~n233 ) ;
  assign n235 = n231 | n234 ;
  assign n236 = n231 & n234 ;
  assign n237 = n235 & ~n236 ;
  assign n238 = n228 & n237 ;
  assign n239 = n74 & n81 ;
  assign n240 = n213 | n239 ;
  assign n241 = n68 & n107 ;
  assign n242 = n180 | n241 ;
  assign n243 = n191 | n242 ;
  assign n244 = n240 | n243 ;
  assign n245 = n81 & n111 ;
  assign n246 = n108 | n245 ;
  assign n247 = n91 & n106 ;
  assign n248 = n136 | n247 ;
  assign n249 = ( n74 & n106 ) | ( n74 & n248 ) | ( n106 & n248 ) ;
  assign n250 = n246 | n249 ;
  assign n251 = n77 & n144 ;
  assign n252 = n42 & n251 ;
  assign n253 = n57 & n144 ;
  assign n254 = n252 | n253 ;
  assign n255 = n250 | n254 ;
  assign n256 = n244 | n255 ;
  assign n257 = n109 & n158 ;
  assign n258 = n198 | n257 ;
  assign n259 = n117 & n174 ;
  assign n260 = n96 | n259 ;
  assign n261 = n126 & n174 ;
  assign n262 = n98 & n157 ;
  assign n263 = n57 & n262 ;
  assign n264 = n261 | n263 ;
  assign n265 = n260 | n264 ;
  assign n266 = n258 | n265 ;
  assign n267 = ~n42 & n154 ;
  assign n268 = n113 & n189 ;
  assign n269 = n267 | n268 ;
  assign n270 = n159 | n161 ;
  assign n271 = n269 | n270 ;
  assign n272 = n57 & n139 ;
  assign n273 = n80 | n272 ;
  assign n274 = n271 | n273 ;
  assign n275 = n266 | n274 ;
  assign n276 = n256 | n275 ;
  assign n277 = n111 & n126 ;
  assign n278 = n68 & n109 ;
  assign n279 = n109 & n262 ;
  assign n280 = n278 | n279 ;
  assign n281 = n277 | n280 ;
  assign n282 = n117 & n139 ;
  assign n283 = n42 & n154 ;
  assign n284 = n282 | n283 ;
  assign n285 = n281 | n284 ;
  assign n286 = ~n79 & n158 ;
  assign n287 = n107 & n174 ;
  assign n288 = n286 | n287 ;
  assign n289 = n285 | n288 ;
  assign n290 = ~n42 & n251 ;
  assign n291 = n109 & n128 ;
  assign n292 = n290 | n291 ;
  assign n293 = n109 & n189 ;
  assign n294 = n129 | n293 ;
  assign n295 = n175 | n294 ;
  assign n296 = n292 | n295 ;
  assign n297 = n107 & n139 ;
  assign n298 = n81 & n128 ;
  assign n299 = n297 | n298 ;
  assign n300 = n117 & n262 ;
  assign n301 = n91 | n174 ;
  assign n302 = n56 & n301 ;
  assign n303 = ~n42 & n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = n299 | n304 ;
  assign n306 = n296 | n305 ;
  assign n307 = n289 | n306 ;
  assign n308 = n276 | n307 ;
  assign n309 = n106 & n189 ;
  assign n310 = n81 & ~n85 ;
  assign n311 = n110 & n310 ;
  assign n312 = ~n79 & n111 ;
  assign n313 = n311 | n312 ;
  assign n314 = n309 | n313 ;
  assign n315 = n81 & n139 ;
  assign n316 = n87 | n130 ;
  assign n317 = n315 | n316 ;
  assign n318 = n314 | n317 ;
  assign n319 = n91 & n117 ;
  assign n320 = n118 | n319 ;
  assign n321 = n101 & n126 ;
  assign n322 = n113 & n262 ;
  assign n323 = n321 | n322 ;
  assign n324 = n320 | n323 ;
  assign n325 = n121 | n173 ;
  assign n326 = n207 | n325 ;
  assign n327 = n324 | n326 ;
  assign n328 = n107 & n144 ;
  assign n329 = n111 & n113 ;
  assign n330 = n328 | n329 ;
  assign n331 = ~n79 & n139 ;
  assign n332 = n149 | n331 ;
  assign n333 = n330 | n332 ;
  assign n334 = n77 & n101 ;
  assign n335 = n162 | n334 ;
  assign n336 = n126 & n139 ;
  assign n337 = n68 | n128 ;
  assign n338 = ( n126 & n336 ) | ( n126 & n337 ) | ( n336 & n337 ) ;
  assign n339 = n335 | n338 ;
  assign n340 = n333 | n339 ;
  assign n341 = n327 | n340 ;
  assign n342 = n318 | n341 ;
  assign n343 = n308 | n342 ;
  assign n344 = n126 & n262 ;
  assign n345 = n96 | n344 ;
  assign n346 = n127 | n164 ;
  assign n347 = n345 | n346 ;
  assign n348 = n268 | n329 ;
  assign n349 = n145 | n239 ;
  assign n350 = n348 | n349 ;
  assign n351 = n347 | n350 ;
  assign n352 = n56 & n74 ;
  assign n353 = n294 | n352 ;
  assign n354 = n107 & n262 ;
  assign n355 = n86 & n107 ;
  assign n356 = n354 | n355 ;
  assign n357 = n242 | n356 ;
  assign n358 = n353 | n357 ;
  assign n359 = n351 | n358 ;
  assign n360 = ~n79 & n189 ;
  assign n361 = n328 | n360 ;
  assign n362 = n126 & n192 ;
  assign n363 = n213 | n362 ;
  assign n364 = n361 | n363 ;
  assign n365 = n359 | n364 ;
  assign n366 = n175 | n336 ;
  assign n367 = n365 | n366 ;
  assign n368 = n57 & n111 ;
  assign n369 = n259 | n368 ;
  assign n370 = n118 | n277 ;
  assign n371 = n81 & n262 ;
  assign n372 = ~n79 & n144 ;
  assign n373 = n371 | n372 ;
  assign n374 = n370 | n373 ;
  assign n375 = n369 | n374 ;
  assign n376 = n248 | n312 ;
  assign n377 = n375 | n376 ;
  assign n378 = ~n95 & n126 ;
  assign n379 = n107 & n189 ;
  assign n380 = n378 | n379 ;
  assign n381 = n212 | n319 ;
  assign n382 = n380 | n381 ;
  assign n383 = ~n79 & n262 ;
  assign n384 = n195 | n383 ;
  assign n385 = ~n95 & n109 ;
  assign n386 = n279 | n385 ;
  assign n387 = n384 | n386 ;
  assign n388 = n107 & n192 ;
  assign n389 = n122 & n174 ;
  assign n390 = n388 | n389 ;
  assign n391 = n179 | n267 ;
  assign n392 = n390 | n391 ;
  assign n393 = n387 | n392 ;
  assign n394 = n382 | n393 ;
  assign n395 = n377 | n394 ;
  assign n396 = n367 | n395 ;
  assign n397 = n74 & n107 ;
  assign n398 = n261 | n397 ;
  assign n399 = n102 | n398 ;
  assign n400 = n117 & n189 ;
  assign n401 = n283 | n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = ~n42 & n207 ;
  assign n404 = ~n95 & n113 ;
  assign n405 = ~n79 & n101 ;
  assign n406 = n404 | n405 ;
  assign n407 = n403 | n406 ;
  assign n408 = n322 | n331 ;
  assign n409 = n80 | n408 ;
  assign n410 = n407 | n409 ;
  assign n411 = n402 | n410 ;
  assign n412 = n208 | n297 ;
  assign n413 = n181 | n196 ;
  assign n414 = n412 | n413 ;
  assign n415 = n140 | n170 ;
  assign n416 = n92 | n321 ;
  assign n417 = n415 | n416 ;
  assign n418 = n414 | n417 ;
  assign n419 = n107 & n148 ;
  assign n420 = n109 & n139 ;
  assign n421 = n113 & n192 ;
  assign n422 = n420 | n421 ;
  assign n423 = n419 | n422 ;
  assign n424 = n126 & n189 ;
  assign n425 = n315 | n424 ;
  assign n426 = n246 | n425 ;
  assign n427 = n423 | n426 ;
  assign n428 = n126 & n128 ;
  assign n429 = n171 | n428 ;
  assign n430 = n165 | n429 ;
  assign n431 = n199 | n430 ;
  assign n432 = n427 | n431 ;
  assign n433 = n418 | n432 ;
  assign n434 = n411 | n433 ;
  assign n435 = n396 | n434 ;
  assign n436 = n343 & n435 ;
  assign n437 = n189 | n262 ;
  assign n438 = n77 & n437 ;
  assign n439 = n81 & n174 ;
  assign n440 = n165 | n439 ;
  assign n441 = n272 | n440 ;
  assign n442 = n370 | n441 ;
  assign n443 = n57 & n101 ;
  assign n444 = n290 | n443 ;
  assign n445 = ~n78 & n91 ;
  assign n446 = n321 | n445 ;
  assign n447 = n444 | n446 ;
  assign n448 = n423 | n447 ;
  assign n449 = n442 | n448 ;
  assign n450 = n354 | n388 ;
  assign n451 = n261 | n336 ;
  assign n452 = n150 | n451 ;
  assign n453 = n450 | n452 ;
  assign n454 = n328 | n403 ;
  assign n455 = n297 | n454 ;
  assign n456 = n161 | n455 ;
  assign n457 = n453 | n456 ;
  assign n458 = n449 | n457 ;
  assign n459 = n175 | n287 ;
  assign n460 = n80 | n208 ;
  assign n461 = n459 | n460 ;
  assign n462 = n458 | n461 ;
  assign n463 = n57 & n148 ;
  assign n464 = n300 | n463 ;
  assign n465 = n57 & n86 ;
  assign n466 = n56 & n192 ;
  assign n467 = n465 | n466 ;
  assign n468 = n464 | n467 ;
  assign n469 = n117 & n148 ;
  assign n470 = n263 | n469 ;
  assign n471 = n130 | n470 ;
  assign n472 = n468 | n471 ;
  assign n473 = n140 | n159 ;
  assign n474 = n127 | n473 ;
  assign n475 = n472 | n474 ;
  assign n476 = n117 & n158 ;
  assign n477 = ~n95 & n122 ;
  assign n478 = n476 | n477 ;
  assign n479 = n380 | n478 ;
  assign n480 = n171 | n479 ;
  assign n481 = n344 | n424 ;
  assign n482 = n101 & n109 ;
  assign n483 = n385 | n482 ;
  assign n484 = n481 | n483 ;
  assign n485 = n57 & n158 ;
  assign n486 = n278 | n485 ;
  assign n487 = n164 | n195 ;
  assign n488 = n486 | n487 ;
  assign n489 = n484 | n488 ;
  assign n490 = n480 | n489 ;
  assign n491 = n256 | n490 ;
  assign n492 = n282 | n404 ;
  assign n493 = n312 | n362 ;
  assign n494 = n492 | n493 ;
  assign n495 = n214 | n428 ;
  assign n496 = n257 | n355 ;
  assign n497 = n495 | n496 ;
  assign n498 = n196 | n199 ;
  assign n499 = n497 | n498 ;
  assign n500 = n494 | n499 ;
  assign n501 = n491 | n500 ;
  assign n502 = n475 | n501 ;
  assign n503 = n462 | n502 ;
  assign n504 = n329 | n362 ;
  assign n505 = n81 & n192 ;
  assign n506 = n378 | n505 ;
  assign n507 = n173 | n286 ;
  assign n508 = n506 | n507 ;
  assign n509 = n504 | n508 ;
  assign n510 = n91 & n113 ;
  assign n511 = n80 | n510 ;
  assign n512 = n415 | n511 ;
  assign n513 = n509 | n512 ;
  assign n514 = n79 | n95 ;
  assign n515 = ~n193 & n514 ;
  assign n516 = ~n335 & n515 ;
  assign n517 = ~n280 & n516 ;
  assign n518 = n77 & n174 ;
  assign n519 = n214 | n252 ;
  assign n520 = n518 | n519 ;
  assign n521 = n293 | n371 ;
  assign n522 = n81 & ~n95 ;
  assign n523 = n239 | n522 ;
  assign n524 = n521 | n523 ;
  assign n525 = n520 | n524 ;
  assign n526 = n517 & ~n525 ;
  assign n527 = ~n513 & n526 ;
  assign n528 = n112 | n311 ;
  assign n529 = n87 | n119 ;
  assign n530 = ~n79 & n91 ;
  assign n531 = n141 | n530 ;
  assign n532 = n529 | n531 ;
  assign n533 = n528 | n532 ;
  assign n534 = n113 & n128 ;
  assign n535 = n298 | n534 ;
  assign n536 = n258 | n535 ;
  assign n537 = n533 | n536 ;
  assign n538 = n149 | n383 ;
  assign n539 = n164 | n322 ;
  assign n540 = n292 | n539 ;
  assign n541 = n538 | n540 ;
  assign n542 = n114 | n420 ;
  assign n543 = n121 | n419 ;
  assign n544 = n542 | n543 ;
  assign n545 = n268 | n360 ;
  assign n546 = n544 | n545 ;
  assign n547 = n159 | n388 ;
  assign n548 = n546 | n547 ;
  assign n549 = n541 | n548 ;
  assign n550 = n537 | n549 ;
  assign n551 = n527 & ~n550 ;
  assign n552 = n78 & n551 ;
  assign n553 = ( ~n503 & n551 ) | ( ~n503 & n552 ) | ( n551 & n552 ) ;
  assign n554 = n56 & ~n95 ;
  assign n555 = n552 & ~n554 ;
  assign n556 = ( n438 & n553 ) | ( n438 & ~n555 ) | ( n553 & ~n555 ) ;
  assign n557 = n286 | n298 ;
  assign n558 = ( n68 & ~n78 ) | ( n68 & n557 ) | ( ~n78 & n557 ) ;
  assign n559 = n556 | n558 ;
  assign n560 = n214 | n445 ;
  assign n561 = n439 | n560 ;
  assign n562 = n559 | n561 ;
  assign n563 = n146 | n282 ;
  assign n564 = n267 | n421 ;
  assign n565 = n563 | n564 ;
  assign n566 = n253 | n565 ;
  assign n567 = n165 | n404 ;
  assign n568 = n283 | n385 ;
  assign n569 = n567 | n568 ;
  assign n570 = n566 | n569 ;
  assign n571 = ( n117 & n158 ) | ( n117 & n161 ) | ( n158 & n161 ) ;
  assign n572 = n443 | n571 ;
  assign n573 = n69 | n572 ;
  assign n574 = n188 | n573 ;
  assign n575 = n272 | n329 ;
  assign n576 = n574 | n575 ;
  assign n577 = n485 | n498 ;
  assign n578 = n576 | n577 ;
  assign n579 = n570 | n578 ;
  assign n580 = n562 | n579 ;
  assign n581 = n436 & ~n580 ;
  assign n582 = ( x14 & x22 ) | ( x14 & ~n37 ) | ( x22 & ~n37 ) ;
  assign n583 = x14 | x22 ;
  assign n584 = ( n38 & n582 ) | ( n38 & ~n583 ) | ( n582 & ~n583 ) ;
  assign n585 = n581 & n584 ;
  assign n586 = ~n436 & n580 ;
  assign n587 = n343 | n435 ;
  assign n588 = n584 & ~n587 ;
  assign n589 = n586 & ~n588 ;
  assign n590 = n585 | n589 ;
  assign n591 = n438 | n579 ;
  assign n592 = n190 | n329 ;
  assign n593 = n472 | n592 ;
  assign n594 = n57 & n74 ;
  assign n595 = n400 | n594 ;
  assign n596 = n368 | n595 ;
  assign n597 = n129 | n176 ;
  assign n598 = n181 | n302 ;
  assign n599 = n597 | n598 ;
  assign n600 = n596 | n599 ;
  assign n601 = n593 | n600 ;
  assign n602 = n562 | n601 ;
  assign n603 = ~n591 & n602 ;
  assign n604 = ( x13 & x22 ) | ( x13 & ~n36 ) | ( x22 & ~n36 ) ;
  assign n605 = x13 | x22 ;
  assign n606 = ( n37 & n604 ) | ( n37 & ~n605 ) | ( n604 & ~n605 ) ;
  assign n607 = n603 & n606 ;
  assign n608 = ( x12 & x22 ) | ( x12 & ~n35 ) | ( x22 & ~n35 ) ;
  assign n609 = x12 | x22 ;
  assign n610 = ( n36 & n608 ) | ( n36 & ~n609 ) | ( n608 & ~n609 ) ;
  assign n611 = n138 | n379 ;
  assign n612 = n141 | n424 ;
  assign n613 = n115 | n612 ;
  assign n614 = n77 & n337 ;
  assign n615 = n613 | n614 ;
  assign n616 = n611 | n615 ;
  assign n617 = n106 | n251 ;
  assign n618 = n140 | n617 ;
  assign n619 = n616 | n618 ;
  assign n620 = n242 | n496 ;
  assign n621 = n429 | n620 ;
  assign n622 = n334 | n621 ;
  assign n623 = n321 | n378 ;
  assign n624 = n170 | n420 ;
  assign n625 = n623 | n624 ;
  assign n626 = n91 & n126 ;
  assign n627 = n108 | n328 ;
  assign n628 = n626 | n627 ;
  assign n629 = n625 | n628 ;
  assign n630 = n277 | n397 ;
  assign n631 = n354 | n510 ;
  assign n632 = n630 | n631 ;
  assign n633 = n212 | n518 ;
  assign n634 = n119 | n344 ;
  assign n635 = n633 | n634 ;
  assign n636 = n632 | n635 ;
  assign n637 = n547 | n636 ;
  assign n638 = n629 | n637 ;
  assign n639 = n622 | n638 ;
  assign n640 = n619 | n639 ;
  assign n641 = n610 | n640 ;
  assign n642 = ~n591 & n610 ;
  assign n643 = ( n607 & n641 ) | ( n607 & ~n642 ) | ( n641 & ~n642 ) ;
  assign n644 = ( x11 & x22 ) | ( x11 & ~n34 ) | ( x22 & ~n34 ) ;
  assign n645 = x11 | x22 ;
  assign n646 = ( n35 & n644 ) | ( n35 & ~n645 ) | ( n644 & ~n645 ) ;
  assign n647 = n640 & n646 ;
  assign n648 = ( n590 & ~n643 ) | ( n590 & n647 ) | ( ~n643 & n647 ) ;
  assign n649 = ( n590 & n643 ) | ( n590 & ~n647 ) | ( n643 & ~n647 ) ;
  assign n650 = ( ~n590 & n648 ) | ( ~n590 & n649 ) | ( n648 & n649 ) ;
  assign n651 = n580 & ~n587 ;
  assign n652 = n581 | n651 ;
  assign n653 = n580 | n606 ;
  assign n654 = n580 & n606 ;
  assign n655 = n653 & ~n654 ;
  assign n656 = n652 & n655 ;
  assign n657 = ~n436 & n587 ;
  assign n658 = ( n580 & n584 ) | ( n580 & ~n657 ) | ( n584 & ~n657 ) ;
  assign n659 = n580 | n584 ;
  assign n660 = ( n656 & ~n658 ) | ( n656 & n659 ) | ( ~n658 & n659 ) ;
  assign n661 = ~n580 & n646 ;
  assign n662 = n580 & ~n646 ;
  assign n663 = n661 | n662 ;
  assign n664 = n591 | n640 ;
  assign n665 = ~n663 & n664 ;
  assign n666 = n603 & n610 ;
  assign n667 = n665 | n666 ;
  assign n668 = n42 & n438 ;
  assign n669 = n118 | n668 ;
  assign n670 = n137 | n469 ;
  assign n671 = ( n117 & n158 ) | ( n117 & n176 ) | ( n158 & n176 ) ;
  assign n672 = n670 | n671 ;
  assign n673 = n669 | n672 ;
  assign n674 = n117 & n192 ;
  assign n675 = n145 | n674 ;
  assign n676 = n92 | n368 ;
  assign n677 = n459 | n676 ;
  assign n678 = n675 | n677 ;
  assign n679 = n119 | n505 ;
  assign n680 = n129 | n278 ;
  assign n681 = n679 | n680 ;
  assign n682 = n311 | n372 ;
  assign n683 = n681 | n682 ;
  assign n684 = n678 | n683 ;
  assign n685 = n673 | n684 ;
  assign n686 = n141 | n465 ;
  assign n687 = n70 | n315 ;
  assign n688 = n686 | n687 ;
  assign n689 = n121 | n212 ;
  assign n690 = n688 | n689 ;
  assign n691 = n196 | n421 ;
  assign n692 = n482 | n691 ;
  assign n693 = n690 | n692 ;
  assign n694 = n344 | n378 ;
  assign n695 = n181 | n694 ;
  assign n696 = n251 | n354 ;
  assign n697 = n87 | n696 ;
  assign n698 = n695 | n697 ;
  assign n699 = n214 | n286 ;
  assign n700 = n263 | n443 ;
  assign n701 = n699 | n700 ;
  assign n702 = n388 | n522 ;
  assign n703 = n172 | n702 ;
  assign n704 = n701 | n703 ;
  assign n705 = n698 | n704 ;
  assign n706 = n693 | n705 ;
  assign n707 = n282 | n405 ;
  assign n708 = n80 | n355 ;
  assign n709 = n707 | n708 ;
  assign n710 = n113 & n174 ;
  assign n711 = n253 | n710 ;
  assign n712 = n81 & n437 ;
  assign n713 = n322 | n712 ;
  assign n714 = n711 | n713 ;
  assign n715 = n709 | n714 ;
  assign n716 = n159 | n534 ;
  assign n717 = n398 | n592 ;
  assign n718 = n716 | n717 ;
  assign n719 = n245 | n259 ;
  assign n720 = n530 | n719 ;
  assign n721 = n718 | n720 ;
  assign n722 = n715 | n721 ;
  assign n723 = n706 | n722 ;
  assign n724 = n685 | n723 ;
  assign n725 = n465 | n534 ;
  assign n726 = n150 | n252 ;
  assign n727 = n725 | n726 ;
  assign n728 = n81 & n91 ;
  assign n729 = n319 | n728 ;
  assign n730 = n257 | n272 ;
  assign n731 = n729 | n730 ;
  assign n732 = n727 | n731 ;
  assign n733 = n286 | n485 ;
  assign n734 = n321 | n733 ;
  assign n735 = n282 | n403 ;
  assign n736 = n626 | n735 ;
  assign n737 = n734 | n736 ;
  assign n738 = n732 | n737 ;
  assign n739 = n372 | n419 ;
  assign n740 = n430 | n739 ;
  assign n741 = n738 | n740 ;
  assign n742 = n162 | n505 ;
  assign n743 = n482 | n510 ;
  assign n744 = n742 | n743 ;
  assign n745 = n108 | n209 ;
  assign n746 = n464 | n745 ;
  assign n747 = n120 | n412 ;
  assign n748 = n746 | n747 ;
  assign n749 = n744 | n748 ;
  assign n750 = n214 | n476 ;
  assign n751 = n469 | n750 ;
  assign n752 = n202 | n751 ;
  assign n753 = n87 | n102 ;
  assign n754 = n444 | n753 ;
  assign n755 = n752 | n754 ;
  assign n756 = n749 | n755 ;
  assign n757 = n741 | n756 ;
  assign n758 = n367 | n757 ;
  assign n759 = n724 & n758 ;
  assign n760 = ~n343 & n759 ;
  assign n761 = n584 & n760 ;
  assign n762 = n343 & ~n759 ;
  assign n763 = n724 | n758 ;
  assign n764 = ~n759 & n763 ;
  assign n765 = n343 & n764 ;
  assign n766 = ( ~n584 & n762 ) | ( ~n584 & n765 ) | ( n762 & n765 ) ;
  assign n767 = n761 | n766 ;
  assign n768 = ( x9 & x22 ) | ( x9 & ~n32 ) | ( x22 & ~n32 ) ;
  assign n769 = x9 | x22 ;
  assign n770 = ( n33 & n768 ) | ( n33 & ~n769 ) | ( n768 & ~n769 ) ;
  assign n771 = n640 & n770 ;
  assign n772 = n586 & ~n610 ;
  assign n773 = ~n580 & n587 ;
  assign n774 = n610 & n773 ;
  assign n775 = n772 | n774 ;
  assign n776 = ~n655 & n657 ;
  assign n777 = n655 & n657 ;
  assign n778 = ( n775 & ~n776 ) | ( n775 & n777 ) | ( ~n776 & n777 ) ;
  assign n779 = ( n767 & ~n771 ) | ( n767 & n778 ) | ( ~n771 & n778 ) ;
  assign n780 = ( n660 & n667 ) | ( n660 & n779 ) | ( n667 & n779 ) ;
  assign n781 = ( x10 & x22 ) | ( x10 & ~n33 ) | ( x22 & ~n33 ) ;
  assign n782 = x10 | x22 ;
  assign n783 = ( n34 & n781 ) | ( n34 & ~n782 ) | ( n781 & ~n782 ) ;
  assign n784 = ( n640 & n770 ) | ( n640 & n783 ) | ( n770 & n783 ) ;
  assign n785 = n770 & n783 ;
  assign n786 = ( ~n762 & n784 ) | ( ~n762 & n785 ) | ( n784 & n785 ) ;
  assign n787 = ( ~n770 & n771 ) | ( ~n770 & n786 ) | ( n771 & n786 ) ;
  assign n788 = ( ~n650 & n780 ) | ( ~n650 & n787 ) | ( n780 & n787 ) ;
  assign n789 = ( n650 & n780 ) | ( n650 & n787 ) | ( n780 & n787 ) ;
  assign n790 = ( n650 & n788 ) | ( n650 & ~n789 ) | ( n788 & ~n789 ) ;
  assign n791 = n603 & n646 ;
  assign n792 = ~n591 & n783 ;
  assign n793 = n640 | n783 ;
  assign n794 = ( n791 & ~n792 ) | ( n791 & n793 ) | ( ~n792 & n793 ) ;
  assign n795 = n603 & n783 ;
  assign n796 = ~n591 & n770 ;
  assign n797 = n640 | n770 ;
  assign n798 = ( n795 & ~n796 ) | ( n795 & n797 ) | ( ~n796 & n797 ) ;
  assign n799 = n343 & ~n584 ;
  assign n800 = ~n343 & n584 ;
  assign n801 = ( n764 & n799 ) | ( n764 & n800 ) | ( n799 & n800 ) ;
  assign n802 = n343 & ~n763 ;
  assign n803 = n606 | n802 ;
  assign n804 = n606 & ~n760 ;
  assign n805 = ( n801 & n803 ) | ( n801 & ~n804 ) | ( n803 & ~n804 ) ;
  assign n806 = n652 & ~n663 ;
  assign n807 = n652 & n663 ;
  assign n808 = ( n775 & ~n806 ) | ( n775 & n807 ) | ( ~n806 & n807 ) ;
  assign n809 = ( n798 & n805 ) | ( n798 & n808 ) | ( n805 & n808 ) ;
  assign n810 = ( x7 & x22 ) | ( x7 & ~n30 ) | ( x22 & ~n30 ) ;
  assign n811 = x7 | x22 ;
  assign n812 = ( n31 & n810 ) | ( n31 & ~n811 ) | ( n810 & ~n811 ) ;
  assign n813 = n640 & n812 ;
  assign n814 = n507 | n534 ;
  assign n815 = n702 | n814 ;
  assign n816 = n181 | n485 ;
  assign n817 = n239 | n674 ;
  assign n818 = n816 | n817 ;
  assign n819 = n257 | n297 ;
  assign n820 = n818 | n819 ;
  assign n821 = n815 | n820 ;
  assign n822 = n140 | n328 ;
  assign n823 = n112 | n164 ;
  assign n824 = n822 | n823 ;
  assign n825 = n57 & n204 ;
  assign n826 = n282 | n825 ;
  assign n827 = n612 | n826 ;
  assign n828 = n824 | n827 ;
  assign n829 = n176 | n241 ;
  assign n830 = n385 | n443 ;
  assign n831 = n311 | n830 ;
  assign n832 = n108 | n253 ;
  assign n833 = n80 | n162 ;
  assign n834 = n832 | n833 ;
  assign n835 = n831 | n834 ;
  assign n836 = n829 | n835 ;
  assign n837 = n828 | n836 ;
  assign n838 = n821 | n837 ;
  assign n839 = n129 | n331 ;
  assign n840 = n198 | n428 ;
  assign n841 = n839 | n840 ;
  assign n842 = n633 | n841 ;
  assign n843 = n171 | n530 ;
  assign n844 = n416 | n843 ;
  assign n845 = n114 | n137 ;
  assign n846 = n190 | n510 ;
  assign n847 = n845 | n846 ;
  assign n848 = n844 | n847 ;
  assign n849 = n317 | n441 ;
  assign n850 = n848 | n849 ;
  assign n851 = n842 | n850 ;
  assign n852 = ~n42 & n69 ;
  assign n853 = n336 | n852 ;
  assign n854 = n145 | n853 ;
  assign n855 = n175 | n344 ;
  assign n856 = n203 | n855 ;
  assign n857 = n281 | n856 ;
  assign n858 = n854 | n857 ;
  assign n859 = n252 | n291 ;
  assign n860 = n506 | n859 ;
  assign n861 = ( n113 & n157 ) | ( n113 & n179 ) | ( n157 & n179 ) ;
  assign n862 = n860 | n861 ;
  assign n863 = n149 | n420 ;
  assign n864 = n213 | n300 ;
  assign n865 = n863 | n864 ;
  assign n866 = n119 | n196 ;
  assign n867 = n515 & ~n866 ;
  assign n868 = ~n865 & n867 ;
  assign n869 = ~n862 & n868 ;
  assign n870 = ~n858 & n869 ;
  assign n871 = ~n851 & n870 ;
  assign n872 = ~n838 & n871 ;
  assign n873 = n263 | n594 ;
  assign n874 = n130 | n213 ;
  assign n875 = n873 | n874 ;
  assign n876 = n70 | n283 ;
  assign n877 = n319 | n876 ;
  assign n878 = n716 | n877 ;
  assign n879 = n875 | n878 ;
  assign n880 = n181 | n852 ;
  assign n881 = n279 | n880 ;
  assign n882 = n325 | n881 ;
  assign n883 = n92 | n510 ;
  assign n884 = n331 | n883 ;
  assign n885 = n138 | n884 ;
  assign n886 = n882 | n885 ;
  assign n887 = n879 | n886 ;
  assign n888 = n114 | n385 ;
  assign n889 = n298 | n315 ;
  assign n890 = n888 | n889 ;
  assign n891 = n519 | n890 ;
  assign n892 = n108 | n465 ;
  assign n893 = n710 | n892 ;
  assign n894 = n891 | n893 ;
  assign n895 = n351 | n894 ;
  assign n896 = n887 | n895 ;
  assign n897 = n462 | n896 ;
  assign n898 = ~n872 & n897 ;
  assign n899 = n724 & ~n898 ;
  assign n900 = ( x8 & x22 ) | ( x8 & ~n31 ) | ( x22 & ~n31 ) ;
  assign n901 = x8 | x22 ;
  assign n902 = ( n32 & n900 ) | ( n32 & ~n901 ) | ( n900 & ~n901 ) ;
  assign n903 = ( ~n640 & n812 ) | ( ~n640 & n902 ) | ( n812 & n902 ) ;
  assign n904 = n812 | n902 ;
  assign n905 = ( n899 & ~n903 ) | ( n899 & n904 ) | ( ~n903 & n904 ) ;
  assign n906 = ( n899 & n903 ) | ( n899 & n904 ) | ( n903 & n904 ) ;
  assign n907 = ( n903 & n905 ) | ( n903 & ~n906 ) | ( n905 & ~n906 ) ;
  assign n908 = ( n813 & ~n899 ) | ( n813 & n907 ) | ( ~n899 & n907 ) ;
  assign n909 = ( n794 & n809 ) | ( n794 & n908 ) | ( n809 & n908 ) ;
  assign n910 = ( n762 & n784 ) | ( n762 & ~n785 ) | ( n784 & ~n785 ) ;
  assign n911 = ( ~n784 & n786 ) | ( ~n784 & n910 ) | ( n786 & n910 ) ;
  assign n912 = ( ~n660 & n667 ) | ( ~n660 & n779 ) | ( n667 & n779 ) ;
  assign n913 = ( n660 & ~n780 ) | ( n660 & n912 ) | ( ~n780 & n912 ) ;
  assign n914 = ( n909 & ~n911 ) | ( n909 & n913 ) | ( ~n911 & n913 ) ;
  assign n915 = n872 & ~n897 ;
  assign n916 = n898 | n915 ;
  assign n917 = n724 & ~n916 ;
  assign n918 = ~n724 & n898 ;
  assign n919 = n584 & ~n918 ;
  assign n920 = n584 | n899 ;
  assign n921 = ( n917 & ~n919 ) | ( n917 & n920 ) | ( ~n919 & n920 ) ;
  assign n922 = n760 | n802 ;
  assign n923 = n610 & ~n724 ;
  assign n924 = ~n610 & n724 ;
  assign n925 = n923 | n924 ;
  assign n926 = n922 & ~n925 ;
  assign n927 = ~n343 & n764 ;
  assign n928 = n606 & ~n927 ;
  assign n929 = n606 | n765 ;
  assign n930 = ( n926 & ~n928 ) | ( n926 & n929 ) | ( ~n928 & n929 ) ;
  assign n931 = ( ~n813 & n921 ) | ( ~n813 & n930 ) | ( n921 & n930 ) ;
  assign n932 = n603 & n770 ;
  assign n933 = n640 | n902 ;
  assign n934 = ~n591 & n902 ;
  assign n935 = ( n932 & n933 ) | ( n932 & ~n934 ) | ( n933 & ~n934 ) ;
  assign n936 = n440 | n623 ;
  assign n937 = n176 | n522 ;
  assign n938 = n463 | n937 ;
  assign n939 = n936 | n938 ;
  assign n940 = n160 | n939 ;
  assign n941 = n77 & n262 ;
  assign n942 = n162 | n941 ;
  assign n943 = n197 | n942 ;
  assign n944 = n212 | n476 ;
  assign n945 = n816 | n944 ;
  assign n946 = n943 | n945 ;
  assign n947 = n207 | n510 ;
  assign n948 = ( ~n208 & n259 ) | ( ~n208 & n947 ) | ( n259 & n947 ) ;
  assign n949 = n946 | n948 ;
  assign n950 = n77 & n128 ;
  assign n951 = n300 | n950 ;
  assign n952 = n69 | n951 ;
  assign n953 = n147 | n952 ;
  assign n954 = n314 | n953 ;
  assign n955 = n949 | n954 ;
  assign n956 = n940 | n955 ;
  assign n957 = n329 | n466 ;
  assign n958 = n191 | n957 ;
  assign n959 = n149 | n282 ;
  assign n960 = n958 | n959 ;
  assign n961 = n453 | n960 ;
  assign n962 = n208 | n405 ;
  assign n963 = n92 | n267 ;
  assign n964 = n962 | n963 ;
  assign n965 = n290 | n888 ;
  assign n966 = n299 | n965 ;
  assign n967 = n964 | n966 ;
  assign n968 = n961 | n967 ;
  assign n969 = n443 | n728 ;
  assign n970 = n164 | n209 ;
  assign n971 = n969 | n970 ;
  assign n972 = n252 | n469 ;
  assign n973 = n708 | n972 ;
  assign n974 = n971 | n973 ;
  assign n975 = n331 | n383 ;
  assign n976 = n136 | n344 ;
  assign n977 = ~n119 & n514 ;
  assign n978 = ~n976 & n977 ;
  assign n979 = ~n975 & n978 ;
  assign n980 = ~n974 & n979 ;
  assign n981 = ~n968 & n980 ;
  assign n982 = ~n956 & n981 ;
  assign n983 = n399 | n953 ;
  assign n984 = n208 | n277 ;
  assign n985 = n686 | n984 ;
  assign n986 = n361 | n985 ;
  assign n987 = n297 | n319 ;
  assign n988 = n175 | n987 ;
  assign n989 = n180 | n481 ;
  assign n990 = n988 | n989 ;
  assign n991 = n986 | n990 ;
  assign n992 = n983 | n991 ;
  assign n993 = n199 | n728 ;
  assign n994 = n383 | n993 ;
  assign n995 = n336 | n866 ;
  assign n996 = n994 | n995 ;
  assign n997 = n213 | n404 ;
  assign n998 = n996 | n997 ;
  assign n999 = n992 | n998 ;
  assign n1000 = n129 | n171 ;
  assign n1001 = n572 | n829 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = n999 | n1002 ;
  assign n1004 = n253 | n354 ;
  assign n1005 = n485 | n1004 ;
  assign n1006 = n203 | n707 ;
  assign n1007 = n611 | n1006 ;
  assign n1008 = n1005 | n1007 ;
  assign n1009 = n96 | n401 ;
  assign n1010 = n463 | n873 ;
  assign n1011 = n1009 | n1010 ;
  assign n1012 = n1008 | n1011 ;
  assign n1013 = n527 & ~n1012 ;
  assign n1014 = ~n1003 & n1013 ;
  assign n1015 = n982 | n1014 ;
  assign n1016 = ~n872 & n1015 ;
  assign n1017 = ( x6 & x22 ) | ( x6 & ~n29 ) | ( x22 & ~n29 ) ;
  assign n1018 = x6 | x22 ;
  assign n1019 = ( n30 & n1017 ) | ( n30 & ~n1018 ) | ( n1017 & ~n1018 ) ;
  assign n1020 = n640 & n1019 ;
  assign n1021 = ( n982 & ~n1016 ) | ( n982 & n1020 ) | ( ~n1016 & n1020 ) ;
  assign n1022 = n343 | n783 ;
  assign n1023 = n343 & n783 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1025 = n652 & ~n1024 ;
  assign n1026 = n657 & n663 ;
  assign n1027 = n1025 | n1026 ;
  assign n1028 = ( n935 & n1021 ) | ( n935 & n1027 ) | ( n1021 & n1027 ) ;
  assign n1029 = ( ~n907 & n931 ) | ( ~n907 & n1028 ) | ( n931 & n1028 ) ;
  assign n1030 = ( n794 & n809 ) | ( n794 & ~n908 ) | ( n809 & ~n908 ) ;
  assign n1031 = ( n908 & ~n909 ) | ( n908 & n1030 ) | ( ~n909 & n1030 ) ;
  assign n1032 = ( n767 & n771 ) | ( n767 & n778 ) | ( n771 & n778 ) ;
  assign n1033 = ( n771 & n779 ) | ( n771 & ~n1032 ) | ( n779 & ~n1032 ) ;
  assign n1034 = ( n1029 & n1031 ) | ( n1029 & ~n1033 ) | ( n1031 & ~n1033 ) ;
  assign n1035 = ( n909 & n911 ) | ( n909 & ~n913 ) | ( n911 & ~n913 ) ;
  assign n1036 = ( ~n909 & n914 ) | ( ~n909 & n1035 ) | ( n914 & n1035 ) ;
  assign n1037 = n603 & n902 ;
  assign n1038 = ~n591 & n812 ;
  assign n1039 = n640 | n812 ;
  assign n1040 = ( n1037 & ~n1038 ) | ( n1037 & n1039 ) | ( ~n1038 & n1039 ) ;
  assign n1041 = n724 & n915 ;
  assign n1042 = n918 | n1041 ;
  assign n1043 = n606 | n724 ;
  assign n1044 = n606 & n724 ;
  assign n1045 = n1043 & ~n1044 ;
  assign n1046 = n1042 & n1045 ;
  assign n1047 = n724 | n916 ;
  assign n1048 = n584 & n1047 ;
  assign n1049 = n584 | n917 ;
  assign n1050 = ( n1046 & ~n1048 ) | ( n1046 & n1049 ) | ( ~n1048 & n1049 ) ;
  assign n1051 = n580 | n770 ;
  assign n1052 = n580 & n770 ;
  assign n1053 = n1051 & ~n1052 ;
  assign n1054 = n652 & n1053 ;
  assign n1055 = ( n580 & ~n657 ) | ( n580 & n783 ) | ( ~n657 & n783 ) ;
  assign n1056 = n580 | n783 ;
  assign n1057 = ( n1054 & ~n1055 ) | ( n1054 & n1056 ) | ( ~n1055 & n1056 ) ;
  assign n1058 = ( n1040 & n1050 ) | ( n1040 & n1057 ) | ( n1050 & n1057 ) ;
  assign n1059 = ( n813 & n921 ) | ( n813 & n930 ) | ( n921 & n930 ) ;
  assign n1060 = ( n813 & n931 ) | ( n813 & ~n1059 ) | ( n931 & ~n1059 ) ;
  assign n1061 = ( ~n935 & n1021 ) | ( ~n935 & n1027 ) | ( n1021 & n1027 ) ;
  assign n1062 = ( n935 & ~n1028 ) | ( n935 & n1061 ) | ( ~n1028 & n1061 ) ;
  assign n1063 = ( n1058 & ~n1060 ) | ( n1058 & n1062 ) | ( ~n1060 & n1062 ) ;
  assign n1064 = ( n907 & n931 ) | ( n907 & ~n1028 ) | ( n931 & ~n1028 ) ;
  assign n1065 = ( ~n931 & n1029 ) | ( ~n931 & n1064 ) | ( n1029 & n1064 ) ;
  assign n1066 = ( ~n798 & n805 ) | ( ~n798 & n808 ) | ( n805 & n808 ) ;
  assign n1067 = ( n798 & ~n809 ) | ( n798 & n1066 ) | ( ~n809 & n1066 ) ;
  assign n1068 = ( n1063 & ~n1065 ) | ( n1063 & n1067 ) | ( ~n1065 & n1067 ) ;
  assign n1069 = ( n1058 & n1060 ) | ( n1058 & ~n1062 ) | ( n1060 & ~n1062 ) ;
  assign n1070 = ( ~n1058 & n1063 ) | ( ~n1058 & n1069 ) | ( n1063 & n1069 ) ;
  assign n1071 = ~n646 & n762 ;
  assign n1072 = ~n343 & n646 ;
  assign n1073 = n763 & n1072 ;
  assign n1074 = n1071 | n1073 ;
  assign n1075 = n610 | n646 ;
  assign n1076 = n610 & n646 ;
  assign n1077 = n1075 & ~n1076 ;
  assign n1078 = n764 & n1077 ;
  assign n1079 = ~n1074 & n1078 ;
  assign n1080 = n1074 & ~n1078 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = ( ~n982 & n1016 ) | ( ~n982 & n1020 ) | ( n1016 & n1020 ) ;
  assign n1083 = ( n982 & n1016 ) | ( n982 & n1020 ) | ( n1016 & n1020 ) ;
  assign n1084 = ( n982 & n1082 ) | ( n982 & ~n1083 ) | ( n1082 & ~n1083 ) ;
  assign n1085 = n222 & n640 ;
  assign n1086 = n982 & n1016 ;
  assign n1087 = n982 | n1016 ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = ~n1085 & n1088 ;
  assign n1090 = n872 & ~n1015 ;
  assign n1091 = n982 & n1014 ;
  assign n1092 = ~n872 & n1091 ;
  assign n1093 = n1090 | n1092 ;
  assign n1094 = n584 & n1093 ;
  assign n1095 = ( n1085 & n1088 ) | ( n1085 & n1094 ) | ( n1088 & n1094 ) ;
  assign n1096 = n1085 | n1094 ;
  assign n1097 = ( n1089 & ~n1095 ) | ( n1089 & n1096 ) | ( ~n1095 & n1096 ) ;
  assign n1098 = ( ~n982 & n1085 ) | ( ~n982 & n1097 ) | ( n1085 & n1097 ) ;
  assign n1099 = ( n1081 & ~n1084 ) | ( n1081 & n1098 ) | ( ~n1084 & n1098 ) ;
  assign n1100 = ( ~n1040 & n1050 ) | ( ~n1040 & n1057 ) | ( n1050 & n1057 ) ;
  assign n1101 = ( n1040 & ~n1058 ) | ( n1040 & n1100 ) | ( ~n1058 & n1100 ) ;
  assign n1102 = n925 & n1042 ;
  assign n1103 = ~n916 & n1045 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = n922 & ~n1024 ;
  assign n1106 = n922 | n1074 ;
  assign n1107 = ~n1105 & n1106 ;
  assign n1108 = n657 & n1053 ;
  assign n1109 = ( n580 & n652 ) | ( n580 & n902 ) | ( n652 & n902 ) ;
  assign n1110 = n580 & n902 ;
  assign n1111 = ( n1108 & n1109 ) | ( n1108 & ~n1110 ) | ( n1109 & ~n1110 ) ;
  assign n1112 = ( n1104 & n1107 ) | ( n1104 & n1111 ) | ( n1107 & n1111 ) ;
  assign n1113 = n603 & n812 ;
  assign n1114 = ~n591 & n1019 ;
  assign n1115 = n640 | n1019 ;
  assign n1116 = ( n1113 & ~n1114 ) | ( n1113 & n1115 ) | ( ~n1114 & n1115 ) ;
  assign n1117 = n225 & n640 ;
  assign n1118 = n606 & n1093 ;
  assign n1119 = n1088 | n1118 ;
  assign n1120 = n1015 & ~n1091 ;
  assign n1121 = n584 & n1120 ;
  assign n1122 = ( n1117 & n1119 ) | ( n1117 & n1121 ) | ( n1119 & n1121 ) ;
  assign n1123 = ( n1117 & ~n1119 ) | ( n1117 & n1121 ) | ( ~n1119 & n1121 ) ;
  assign n1124 = ( n1119 & ~n1122 ) | ( n1119 & n1123 ) | ( ~n1122 & n1123 ) ;
  assign n1125 = ( ~n982 & n1117 ) | ( ~n982 & n1124 ) | ( n1117 & n1124 ) ;
  assign n1126 = n764 & n1024 ;
  assign n1127 = ~n760 & n770 ;
  assign n1128 = n770 | n802 ;
  assign n1129 = ( n1126 & ~n1127 ) | ( n1126 & n1128 ) | ( ~n1127 & n1128 ) ;
  assign n1130 = ~n916 & n925 ;
  assign n1131 = n646 & n872 ;
  assign n1132 = n646 | n872 ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = n1042 & n1133 ;
  assign n1135 = n1130 | n1134 ;
  assign n1136 = ~n580 & n812 ;
  assign n1137 = n580 & ~n812 ;
  assign n1138 = ( n652 & n1136 ) | ( n652 & n1137 ) | ( n1136 & n1137 ) ;
  assign n1139 = ( n580 & n657 ) | ( n580 & n902 ) | ( n657 & n902 ) ;
  assign n1140 = ( ~n1110 & n1138 ) | ( ~n1110 & n1139 ) | ( n1138 & n1139 ) ;
  assign n1141 = ( n1129 & n1135 ) | ( n1129 & n1140 ) | ( n1135 & n1140 ) ;
  assign n1142 = ( n1116 & n1125 ) | ( n1116 & n1141 ) | ( n1125 & n1141 ) ;
  assign n1143 = ( n1101 & n1112 ) | ( n1101 & n1142 ) | ( n1112 & n1142 ) ;
  assign n1144 = ( ~n1070 & n1099 ) | ( ~n1070 & n1143 ) | ( n1099 & n1143 ) ;
  assign n1145 = n603 & n1019 ;
  assign n1146 = n222 | n640 ;
  assign n1147 = n222 & ~n591 ;
  assign n1148 = ( n1145 & n1146 ) | ( n1145 & ~n1147 ) | ( n1146 & ~n1147 ) ;
  assign n1149 = n610 & n872 ;
  assign n1150 = n610 | n872 ;
  assign n1151 = ~n1149 & n1150 ;
  assign n1152 = n1093 & ~n1151 ;
  assign n1153 = ( ~n606 & n872 ) | ( ~n606 & n1120 ) | ( n872 & n1120 ) ;
  assign n1154 = ~n606 & n872 ;
  assign n1155 = ( n1152 & n1153 ) | ( n1152 & ~n1154 ) | ( n1153 & ~n1154 ) ;
  assign n1156 = n234 & n640 ;
  assign n1157 = n70 | n272 ;
  assign n1158 = n495 | n1157 ;
  assign n1159 = n994 | n1158 ;
  assign n1160 = n287 | n406 ;
  assign n1161 = n138 | n1160 ;
  assign n1162 = n862 | n1161 ;
  assign n1163 = n1159 | n1162 ;
  assign n1164 = n846 | n863 ;
  assign n1165 = n725 | n1164 ;
  assign n1166 = n290 | n482 ;
  assign n1167 = n310 | n1166 ;
  assign n1168 = n1165 | n1167 ;
  assign n1169 = n379 | n469 ;
  assign n1170 = n112 | n1169 ;
  assign n1171 = n277 | n385 ;
  assign n1172 = n1170 | n1171 ;
  assign n1173 = n418 | n1172 ;
  assign n1174 = n1168 | n1173 ;
  assign n1175 = n1163 | n1174 ;
  assign n1176 = n129 | n239 ;
  assign n1177 = n92 | n179 ;
  assign n1178 = n1176 | n1177 ;
  assign n1179 = n568 | n1178 ;
  assign n1180 = n95 & ~n1179 ;
  assign n1181 = ( n1175 & ~n1179 ) | ( n1175 & n1180 ) | ( ~n1179 & n1180 ) ;
  assign n1182 = n130 | n1160 ;
  assign n1183 = n727 | n1182 ;
  assign n1184 = n378 | n710 ;
  assign n1185 = n277 | n331 ;
  assign n1186 = n363 | n1185 ;
  assign n1187 = n1184 | n1186 ;
  assign n1188 = n271 | n1187 ;
  assign n1189 = n1183 | n1188 ;
  assign n1190 = n273 | n866 ;
  assign n1191 = n959 | n1190 ;
  assign n1192 = n173 | n424 ;
  assign n1193 = n200 | n1192 ;
  assign n1194 = n1191 | n1193 ;
  assign n1195 = n193 | n400 ;
  assign n1196 = ( n107 & n158 ) | ( n107 & n379 ) | ( n158 & n379 ) ;
  assign n1197 = n373 | n1196 ;
  assign n1198 = n1195 | n1197 ;
  assign n1199 = n300 | n482 ;
  assign n1200 = n384 | n1199 ;
  assign n1201 = n621 | n1200 ;
  assign n1202 = n1198 | n1201 ;
  assign n1203 = n1194 | n1202 ;
  assign n1204 = n1189 | n1203 ;
  assign n1205 = n1181 & ~n1204 ;
  assign n1206 = n982 | n1205 ;
  assign n1207 = ( n584 & n982 ) | ( n584 & n1206 ) | ( n982 & n1206 ) ;
  assign n1208 = ( n1155 & n1156 ) | ( n1155 & ~n1207 ) | ( n1156 & ~n1207 ) ;
  assign n1209 = ~n783 & n872 ;
  assign n1210 = n783 & ~n872 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = n1042 & n1211 ;
  assign n1213 = n646 | n917 ;
  assign n1214 = n646 & n1047 ;
  assign n1215 = ( n1212 & n1213 ) | ( n1212 & ~n1214 ) | ( n1213 & ~n1214 ) ;
  assign n1216 = n343 & ~n770 ;
  assign n1217 = ~n343 & n770 ;
  assign n1218 = ( n764 & n1216 ) | ( n764 & n1217 ) | ( n1216 & n1217 ) ;
  assign n1219 = ~n760 & n902 ;
  assign n1220 = n802 | n902 ;
  assign n1221 = ( n1218 & ~n1219 ) | ( n1218 & n1220 ) | ( ~n1219 & n1220 ) ;
  assign n1222 = n343 | n1019 ;
  assign n1223 = n343 & n1019 ;
  assign n1224 = n1222 & ~n1223 ;
  assign n1225 = n652 & ~n1224 ;
  assign n1226 = ( n580 & ~n657 ) | ( n580 & n812 ) | ( ~n657 & n812 ) ;
  assign n1227 = n580 | n812 ;
  assign n1228 = ( n1225 & ~n1226 ) | ( n1225 & n1227 ) | ( ~n1226 & n1227 ) ;
  assign n1229 = ( n1215 & n1221 ) | ( n1215 & n1228 ) | ( n1221 & n1228 ) ;
  assign n1230 = ( n1148 & n1208 ) | ( n1148 & n1229 ) | ( n1208 & n1229 ) ;
  assign n1231 = ( n1104 & ~n1107 ) | ( n1104 & n1111 ) | ( ~n1107 & n1111 ) ;
  assign n1232 = ( n1107 & ~n1112 ) | ( n1107 & n1231 ) | ( ~n1112 & n1231 ) ;
  assign n1233 = ( ~n1097 & n1230 ) | ( ~n1097 & n1232 ) | ( n1230 & n1232 ) ;
  assign n1234 = ( n1081 & n1084 ) | ( n1081 & ~n1098 ) | ( n1084 & ~n1098 ) ;
  assign n1235 = ( ~n1081 & n1099 ) | ( ~n1081 & n1234 ) | ( n1099 & n1234 ) ;
  assign n1236 = ( ~n1101 & n1112 ) | ( ~n1101 & n1142 ) | ( n1112 & n1142 ) ;
  assign n1237 = ( n1101 & ~n1143 ) | ( n1101 & n1236 ) | ( ~n1143 & n1236 ) ;
  assign n1238 = ( n1233 & ~n1235 ) | ( n1233 & n1237 ) | ( ~n1235 & n1237 ) ;
  assign n1239 = ( n1233 & n1235 ) | ( n1233 & ~n1237 ) | ( n1235 & ~n1237 ) ;
  assign n1240 = ( ~n1233 & n1238 ) | ( ~n1233 & n1239 ) | ( n1238 & n1239 ) ;
  assign n1241 = ( n1097 & n1230 ) | ( n1097 & n1232 ) | ( n1230 & n1232 ) ;
  assign n1242 = ( n1097 & n1233 ) | ( n1097 & ~n1241 ) | ( n1233 & ~n1241 ) ;
  assign n1243 = ( ~n1116 & n1125 ) | ( ~n1116 & n1141 ) | ( n1125 & n1141 ) ;
  assign n1244 = ( n1116 & ~n1142 ) | ( n1116 & n1243 ) | ( ~n1142 & n1243 ) ;
  assign n1245 = ( ~n1129 & n1135 ) | ( ~n1129 & n1140 ) | ( n1135 & n1140 ) ;
  assign n1246 = ( n1129 & ~n1141 ) | ( n1129 & n1245 ) | ( ~n1141 & n1245 ) ;
  assign n1247 = ~n982 & n1205 ;
  assign n1248 = ~n606 & n1247 ;
  assign n1249 = n982 & ~n1205 ;
  assign n1250 = n584 & ~n1249 ;
  assign n1251 = ~n584 & n1206 ;
  assign n1252 = ( ~n1248 & n1250 ) | ( ~n1248 & n1251 ) | ( n1250 & n1251 ) ;
  assign n1253 = n640 & ~n1252 ;
  assign n1254 = n222 & n603 ;
  assign n1255 = n225 | n640 ;
  assign n1256 = n225 & ~n591 ;
  assign n1257 = ( n1254 & n1255 ) | ( n1254 & ~n1256 ) | ( n1255 & ~n1256 ) ;
  assign n1258 = ~n343 & n902 ;
  assign n1259 = n343 & ~n902 ;
  assign n1260 = ( n764 & n1258 ) | ( n764 & n1259 ) | ( n1258 & n1259 ) ;
  assign n1261 = n802 | n812 ;
  assign n1262 = ~n760 & n812 ;
  assign n1263 = ( n1260 & n1261 ) | ( n1260 & ~n1262 ) | ( n1261 & ~n1262 ) ;
  assign n1264 = ~n770 & n872 ;
  assign n1265 = n770 & ~n872 ;
  assign n1266 = n1264 | n1265 ;
  assign n1267 = n1042 & n1266 ;
  assign n1268 = n783 & n1047 ;
  assign n1269 = n783 | n917 ;
  assign n1270 = ( n1267 & ~n1268 ) | ( n1267 & n1269 ) | ( ~n1268 & n1269 ) ;
  assign n1271 = ~n222 & n586 ;
  assign n1272 = n222 & n773 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = n222 | n1019 ;
  assign n1275 = n222 & n1019 ;
  assign n1276 = n1274 & ~n1275 ;
  assign n1277 = n657 & n1276 ;
  assign n1278 = ~n1273 & n1277 ;
  assign n1279 = n1273 & ~n1277 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = ( n1263 & n1270 ) | ( n1263 & n1280 ) | ( n1270 & n1280 ) ;
  assign n1282 = ( n1253 & n1257 ) | ( n1253 & n1281 ) | ( n1257 & n1281 ) ;
  assign n1283 = ( ~n1124 & n1246 ) | ( ~n1124 & n1282 ) | ( n1246 & n1282 ) ;
  assign n1284 = ( ~n1242 & n1244 ) | ( ~n1242 & n1283 ) | ( n1244 & n1283 ) ;
  assign n1285 = n1120 & ~n1151 ;
  assign n1286 = n1093 & ~n1133 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = ~n640 & n1252 ;
  assign n1289 = n1253 | n1288 ;
  assign n1290 = n225 & n603 ;
  assign n1291 = n234 & ~n591 ;
  assign n1292 = n234 | n640 ;
  assign n1293 = ( n1290 & ~n1291 ) | ( n1290 & n1292 ) | ( ~n1291 & n1292 ) ;
  assign n1294 = ( n1287 & ~n1289 ) | ( n1287 & n1293 ) | ( ~n1289 & n1293 ) ;
  assign n1295 = ( ~n1215 & n1221 ) | ( ~n1215 & n1228 ) | ( n1221 & n1228 ) ;
  assign n1296 = ( n1215 & ~n1229 ) | ( n1215 & n1295 ) | ( ~n1229 & n1295 ) ;
  assign n1297 = ( n1155 & n1156 ) | ( n1155 & n1207 ) | ( n1156 & n1207 ) ;
  assign n1298 = ( n1207 & n1208 ) | ( n1207 & ~n1297 ) | ( n1208 & ~n1297 ) ;
  assign n1299 = ( n1294 & n1296 ) | ( n1294 & ~n1298 ) | ( n1296 & ~n1298 ) ;
  assign n1300 = ( n1124 & n1246 ) | ( n1124 & n1282 ) | ( n1246 & n1282 ) ;
  assign n1301 = ( n1124 & n1283 ) | ( n1124 & ~n1300 ) | ( n1283 & ~n1300 ) ;
  assign n1302 = ( n1148 & ~n1208 ) | ( n1148 & n1229 ) | ( ~n1208 & n1229 ) ;
  assign n1303 = ( n1208 & ~n1230 ) | ( n1208 & n1302 ) | ( ~n1230 & n1302 ) ;
  assign n1304 = ( n1299 & ~n1301 ) | ( n1299 & n1303 ) | ( ~n1301 & n1303 ) ;
  assign n1305 = ( n1299 & n1301 ) | ( n1299 & ~n1303 ) | ( n1301 & ~n1303 ) ;
  assign n1306 = ( ~n1299 & n1304 ) | ( ~n1299 & n1305 ) | ( n1304 & n1305 ) ;
  assign n1307 = n1120 & ~n1133 ;
  assign n1308 = n1093 & ~n1211 ;
  assign n1309 = n1307 | n1308 ;
  assign n1310 = ~n610 & n1247 ;
  assign n1311 = n606 & ~n1249 ;
  assign n1312 = ~n606 & n1206 ;
  assign n1313 = ( ~n1310 & n1311 ) | ( ~n1310 & n1312 ) | ( n1311 & n1312 ) ;
  assign n1314 = n228 & n652 ;
  assign n1315 = ~n1273 & n1314 ;
  assign n1316 = n1273 & ~n1314 ;
  assign n1317 = n1315 | n1316 ;
  assign n1318 = ( n1309 & ~n1313 ) | ( n1309 & n1317 ) | ( ~n1313 & n1317 ) ;
  assign n1319 = n872 & n902 ;
  assign n1320 = n872 | n902 ;
  assign n1321 = ~n1319 & n1320 ;
  assign n1322 = n1042 & n1321 ;
  assign n1323 = n770 & n1047 ;
  assign n1324 = n770 | n917 ;
  assign n1325 = ( n1322 & ~n1323 ) | ( n1322 & n1324 ) | ( ~n1323 & n1324 ) ;
  assign n1326 = n922 & n1224 ;
  assign n1327 = n812 & ~n927 ;
  assign n1328 = n765 | n812 ;
  assign n1329 = ( n1326 & ~n1327 ) | ( n1326 & n1328 ) | ( ~n1327 & n1328 ) ;
  assign n1330 = ~n646 & n1247 ;
  assign n1331 = ~n610 & n1206 ;
  assign n1332 = n610 & ~n1249 ;
  assign n1333 = ( ~n1330 & n1331 ) | ( ~n1330 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = n234 & n657 ;
  assign n1335 = n586 & ~n1334 ;
  assign n1336 = ~n1333 & n1335 ;
  assign n1337 = ( n1325 & n1329 ) | ( n1325 & n1336 ) | ( n1329 & n1336 ) ;
  assign n1338 = ( n1263 & ~n1270 ) | ( n1263 & n1280 ) | ( ~n1270 & n1280 ) ;
  assign n1339 = ( n1270 & ~n1281 ) | ( n1270 & n1338 ) | ( ~n1281 & n1338 ) ;
  assign n1340 = ( n1318 & n1337 ) | ( n1318 & n1339 ) | ( n1337 & n1339 ) ;
  assign n1341 = ( n1253 & ~n1257 ) | ( n1253 & n1281 ) | ( ~n1257 & n1281 ) ;
  assign n1342 = ( n1257 & ~n1282 ) | ( n1257 & n1341 ) | ( ~n1282 & n1341 ) ;
  assign n1343 = ( n1294 & ~n1296 ) | ( n1294 & n1298 ) | ( ~n1296 & n1298 ) ;
  assign n1344 = ( ~n1294 & n1299 ) | ( ~n1294 & n1343 ) | ( n1299 & n1343 ) ;
  assign n1345 = ( n1340 & n1342 ) | ( n1340 & ~n1344 ) | ( n1342 & ~n1344 ) ;
  assign n1346 = n764 & n1224 ;
  assign n1347 = n222 | n802 ;
  assign n1348 = n222 & ~n760 ;
  assign n1349 = ( n1346 & n1347 ) | ( n1346 & ~n1348 ) | ( n1347 & ~n1348 ) ;
  assign n1350 = n724 | n812 ;
  assign n1351 = n724 & n812 ;
  assign n1352 = n1350 & ~n1351 ;
  assign n1353 = n1042 & n1352 ;
  assign n1354 = n902 | n917 ;
  assign n1355 = n902 & n1047 ;
  assign n1356 = ( n1353 & n1354 ) | ( n1353 & ~n1355 ) | ( n1354 & ~n1355 ) ;
  assign n1357 = n1093 & ~n1266 ;
  assign n1358 = n1120 & ~n1211 ;
  assign n1359 = n1357 | n1358 ;
  assign n1360 = ( n1349 & n1356 ) | ( n1349 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1361 = n234 & n603 ;
  assign n1362 = ( n1325 & ~n1329 ) | ( n1325 & n1336 ) | ( ~n1329 & n1336 ) ;
  assign n1363 = ( n1329 & ~n1337 ) | ( n1329 & n1362 ) | ( ~n1337 & n1362 ) ;
  assign n1364 = ( n1360 & n1361 ) | ( n1360 & n1363 ) | ( n1361 & n1363 ) ;
  assign n1365 = ( n1287 & n1289 ) | ( n1287 & n1293 ) | ( n1289 & n1293 ) ;
  assign n1366 = ( n1289 & n1294 ) | ( n1289 & ~n1365 ) | ( n1294 & ~n1365 ) ;
  assign n1367 = ( ~n1318 & n1337 ) | ( ~n1318 & n1339 ) | ( n1337 & n1339 ) ;
  assign n1368 = ( n1318 & ~n1340 ) | ( n1318 & n1367 ) | ( ~n1340 & n1367 ) ;
  assign n1369 = ( n1364 & ~n1366 ) | ( n1364 & n1368 ) | ( ~n1366 & n1368 ) ;
  assign n1370 = ( n1364 & n1366 ) | ( n1364 & ~n1368 ) | ( n1366 & ~n1368 ) ;
  assign n1371 = ( ~n1364 & n1369 ) | ( ~n1364 & n1370 ) | ( n1369 & n1370 ) ;
  assign n1372 = ( n225 & n580 ) | ( n225 & ~n657 ) | ( n580 & ~n657 ) ;
  assign n1373 = ( n225 & n580 ) | ( n225 & n657 ) | ( n580 & n657 ) ;
  assign n1374 = ~n1372 & n1373 ;
  assign n1375 = n234 | n651 ;
  assign n1376 = n234 & ~n581 ;
  assign n1377 = ( n1374 & n1375 ) | ( n1374 & ~n1376 ) | ( n1375 & ~n1376 ) ;
  assign n1378 = ~n916 & n1352 ;
  assign n1379 = n724 | n1019 ;
  assign n1380 = n724 & n1019 ;
  assign n1381 = n1379 & ~n1380 ;
  assign n1382 = n1042 & n1381 ;
  assign n1383 = n1378 | n1382 ;
  assign n1384 = ~n783 & n1247 ;
  assign n1385 = ~n646 & n1206 ;
  assign n1386 = n646 & ~n1249 ;
  assign n1387 = ( ~n1384 & n1385 ) | ( ~n1384 & n1386 ) | ( n1385 & n1386 ) ;
  assign n1388 = n1120 & ~n1266 ;
  assign n1389 = n1093 & ~n1321 ;
  assign n1390 = n1388 | n1389 ;
  assign n1391 = ( n1383 & ~n1387 ) | ( n1383 & n1390 ) | ( ~n1387 & n1390 ) ;
  assign n1392 = n1333 & ~n1335 ;
  assign n1393 = n1336 | n1392 ;
  assign n1394 = ( n1377 & n1391 ) | ( n1377 & ~n1393 ) | ( n1391 & ~n1393 ) ;
  assign n1395 = ( n1360 & n1361 ) | ( n1360 & ~n1363 ) | ( n1361 & ~n1363 ) ;
  assign n1396 = ( n1363 & ~n1364 ) | ( n1363 & n1395 ) | ( ~n1364 & n1395 ) ;
  assign n1397 = ( n1309 & n1313 ) | ( n1309 & n1317 ) | ( n1313 & n1317 ) ;
  assign n1398 = ( n1313 & n1318 ) | ( n1313 & ~n1397 ) | ( n1318 & ~n1397 ) ;
  assign n1399 = ( n1394 & n1396 ) | ( n1394 & ~n1398 ) | ( n1396 & ~n1398 ) ;
  assign n1400 = ( ~n1349 & n1356 ) | ( ~n1349 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1401 = ( n1349 & ~n1360 ) | ( n1349 & n1400 ) | ( ~n1360 & n1400 ) ;
  assign n1402 = ~n770 & n1247 ;
  assign n1403 = n783 & ~n1249 ;
  assign n1404 = ~n783 & n1206 ;
  assign n1405 = ( ~n1402 & n1403 ) | ( ~n1402 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1406 = n234 & n764 ;
  assign n1407 = n762 & ~n1406 ;
  assign n1408 = ~n1405 & n1407 ;
  assign n1409 = ~n222 & n343 ;
  assign n1410 = n222 & ~n343 ;
  assign n1411 = ( n764 & n1409 ) | ( n764 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1412 = n225 & ~n760 ;
  assign n1413 = n225 | n802 ;
  assign n1414 = ( n1411 & ~n1412 ) | ( n1411 & n1413 ) | ( ~n1412 & n1413 ) ;
  assign n1415 = ( n1334 & n1408 ) | ( n1334 & n1414 ) | ( n1408 & n1414 ) ;
  assign n1416 = ( n1377 & ~n1391 ) | ( n1377 & n1393 ) | ( ~n1391 & n1393 ) ;
  assign n1417 = ( ~n1377 & n1394 ) | ( ~n1377 & n1416 ) | ( n1394 & n1416 ) ;
  assign n1418 = ( n1401 & n1415 ) | ( n1401 & ~n1417 ) | ( n1415 & ~n1417 ) ;
  assign n1419 = ( ~n1394 & n1396 ) | ( ~n1394 & n1398 ) | ( n1396 & n1398 ) ;
  assign n1420 = ( ~n1396 & n1399 ) | ( ~n1396 & n1419 ) | ( n1399 & n1419 ) ;
  assign n1421 = ~n1418 & n1420 ;
  assign n1422 = n1418 & ~n1420 ;
  assign n1423 = ~n812 & n872 ;
  assign n1424 = n812 & ~n872 ;
  assign n1425 = n1423 | n1424 ;
  assign n1426 = n1093 & ~n1425 ;
  assign n1427 = n1120 & ~n1321 ;
  assign n1428 = n1426 | n1427 ;
  assign n1429 = ~n225 & n343 ;
  assign n1430 = n225 & ~n343 ;
  assign n1431 = ( n764 & n1429 ) | ( n764 & n1430 ) | ( n1429 & n1430 ) ;
  assign n1432 = n234 | n802 ;
  assign n1433 = n234 & ~n760 ;
  assign n1434 = ( n1431 & n1432 ) | ( n1431 & ~n1433 ) | ( n1432 & ~n1433 ) ;
  assign n1435 = ~n916 & n1381 ;
  assign n1436 = n222 & n872 ;
  assign n1437 = n222 | n872 ;
  assign n1438 = ~n1436 & n1437 ;
  assign n1439 = n1042 & n1438 ;
  assign n1440 = n1435 | n1439 ;
  assign n1441 = ( n1428 & n1434 ) | ( n1428 & n1440 ) | ( n1434 & n1440 ) ;
  assign n1442 = ( n1383 & n1387 ) | ( n1383 & ~n1390 ) | ( n1387 & ~n1390 ) ;
  assign n1443 = ( ~n1383 & n1391 ) | ( ~n1383 & n1442 ) | ( n1391 & n1442 ) ;
  assign n1444 = ( n1334 & ~n1408 ) | ( n1334 & n1414 ) | ( ~n1408 & n1414 ) ;
  assign n1445 = ( n1408 & ~n1415 ) | ( n1408 & n1444 ) | ( ~n1415 & n1444 ) ;
  assign n1446 = ( n1441 & ~n1443 ) | ( n1441 & n1445 ) | ( ~n1443 & n1445 ) ;
  assign n1447 = n872 & ~n1019 ;
  assign n1448 = ~n872 & n1019 ;
  assign n1449 = n1447 | n1448 ;
  assign n1450 = n1093 & ~n1449 ;
  assign n1451 = n1120 & ~n1425 ;
  assign n1452 = n1450 | n1451 ;
  assign n1453 = n225 & n872 ;
  assign n1454 = n225 | n872 ;
  assign n1455 = ~n1453 & n1454 ;
  assign n1456 = n1042 & n1455 ;
  assign n1457 = n222 | n917 ;
  assign n1458 = n222 & n1047 ;
  assign n1459 = ( n1456 & n1457 ) | ( n1456 & ~n1458 ) | ( n1457 & ~n1458 ) ;
  assign n1460 = ~n902 & n1247 ;
  assign n1461 = n770 & ~n1249 ;
  assign n1462 = ~n770 & n1206 ;
  assign n1463 = ( ~n1460 & n1461 ) | ( ~n1460 & n1462 ) | ( n1461 & n1462 ) ;
  assign n1464 = ( n1452 & n1459 ) | ( n1452 & ~n1463 ) | ( n1459 & ~n1463 ) ;
  assign n1465 = n1405 & ~n1407 ;
  assign n1466 = n1408 | n1465 ;
  assign n1467 = ( ~n1428 & n1434 ) | ( ~n1428 & n1440 ) | ( n1434 & n1440 ) ;
  assign n1468 = ( n1428 & ~n1441 ) | ( n1428 & n1467 ) | ( ~n1441 & n1467 ) ;
  assign n1469 = ( n1464 & ~n1466 ) | ( n1464 & n1468 ) | ( ~n1466 & n1468 ) ;
  assign n1470 = ( ~n1441 & n1443 ) | ( ~n1441 & n1445 ) | ( n1443 & n1445 ) ;
  assign n1471 = ( ~n1445 & n1446 ) | ( ~n1445 & n1470 ) | ( n1446 & n1470 ) ;
  assign n1472 = ~n222 & n1247 ;
  assign n1473 = n1019 & ~n1249 ;
  assign n1474 = ~n1019 & n1206 ;
  assign n1475 = ( ~n1472 & n1473 ) | ( ~n1472 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ~n234 & n1016 ;
  assign n1477 = n1092 | n1476 ;
  assign n1478 = ~n1475 & n1477 ;
  assign n1479 = ~n1019 & n1247 ;
  assign n1480 = n812 & ~n1249 ;
  assign n1481 = ~n812 & n1206 ;
  assign n1482 = ( ~n1479 & n1480 ) | ( ~n1479 & n1481 ) | ( n1480 & n1481 ) ;
  assign n1483 = n1120 & ~n1438 ;
  assign n1484 = n1093 & ~n1455 ;
  assign n1485 = n1483 | n1484 ;
  assign n1486 = ( n1478 & ~n1482 ) | ( n1478 & n1485 ) | ( ~n1482 & n1485 ) ;
  assign n1487 = n234 & ~n916 ;
  assign n1488 = n225 | n982 ;
  assign n1489 = n234 & ~n1205 ;
  assign n1490 = n1488 & ~n1489 ;
  assign n1491 = n234 & ~n1120 ;
  assign n1492 = n1490 | n1491 ;
  assign n1493 = n222 & n1206 ;
  assign n1494 = n222 | n982 ;
  assign n1495 = ( n1492 & ~n1493 ) | ( n1492 & n1494 ) | ( ~n1493 & n1494 ) ;
  assign n1496 = n1120 & ~n1455 ;
  assign n1497 = n234 & ~n1090 ;
  assign n1498 = n234 | n1092 ;
  assign n1499 = ( n1496 & ~n1497 ) | ( n1496 & n1498 ) | ( ~n1497 & n1498 ) ;
  assign n1500 = n1475 & n1476 ;
  assign n1501 = n1475 | n1476 ;
  assign n1502 = ~n1500 & n1501 ;
  assign n1503 = ( n1495 & ~n1499 ) | ( n1495 & n1502 ) | ( ~n1499 & n1502 ) ;
  assign n1504 = ( n1478 & n1482 ) | ( n1478 & ~n1485 ) | ( n1482 & ~n1485 ) ;
  assign n1505 = ( ~n1478 & n1486 ) | ( ~n1478 & n1504 ) | ( n1486 & n1504 ) ;
  assign n1506 = ( ~n1487 & n1503 ) | ( ~n1487 & n1505 ) | ( n1503 & n1505 ) ;
  assign n1507 = n1093 & ~n1438 ;
  assign n1508 = n1120 & ~n1449 ;
  assign n1509 = n1507 | n1508 ;
  assign n1510 = ~n225 & n724 ;
  assign n1511 = n225 & ~n724 ;
  assign n1512 = ( ~n916 & n1510 ) | ( ~n916 & n1511 ) | ( n1510 & n1511 ) ;
  assign n1513 = n234 | n1041 ;
  assign n1514 = n234 & ~n918 ;
  assign n1515 = ( n1512 & n1513 ) | ( n1512 & ~n1514 ) | ( n1513 & ~n1514 ) ;
  assign n1516 = ~n812 & n1247 ;
  assign n1517 = ~n902 & n1206 ;
  assign n1518 = n902 & ~n1249 ;
  assign n1519 = ( ~n1516 & n1517 ) | ( ~n1516 & n1518 ) | ( n1517 & n1518 ) ;
  assign n1520 = n899 & ~n1487 ;
  assign n1521 = ~n1519 & n1520 ;
  assign n1522 = n1519 & ~n1520 ;
  assign n1523 = n1521 | n1522 ;
  assign n1524 = ( n1509 & ~n1515 ) | ( n1509 & n1523 ) | ( ~n1515 & n1523 ) ;
  assign n1525 = ( n1509 & n1515 ) | ( n1509 & ~n1523 ) | ( n1515 & ~n1523 ) ;
  assign n1526 = ( ~n1509 & n1524 ) | ( ~n1509 & n1525 ) | ( n1524 & n1525 ) ;
  assign n1527 = ( ~n1486 & n1506 ) | ( ~n1486 & n1526 ) | ( n1506 & n1526 ) ;
  assign n1528 = ( n1452 & ~n1459 ) | ( n1452 & n1463 ) | ( ~n1459 & n1463 ) ;
  assign n1529 = ( ~n1452 & n1464 ) | ( ~n1452 & n1528 ) | ( n1464 & n1528 ) ;
  assign n1530 = n1527 | n1529 ;
  assign n1531 = ( n1464 & n1466 ) | ( n1464 & ~n1468 ) | ( n1466 & ~n1468 ) ;
  assign n1532 = ( ~n1464 & n1469 ) | ( ~n1464 & n1531 ) | ( n1469 & n1531 ) ;
  assign n1533 = n1406 | n1521 ;
  assign n1534 = n1525 | n1533 ;
  assign n1535 = ~n1532 & n1534 ;
  assign n1536 = n1530 & ~n1535 ;
  assign n1537 = ( n1406 & n1521 ) | ( n1406 & n1525 ) | ( n1521 & n1525 ) ;
  assign n1538 = n1527 & n1529 ;
  assign n1539 = n1532 & ~n1537 ;
  assign n1540 = ( ~n1537 & n1538 ) | ( ~n1537 & n1539 ) | ( n1538 & n1539 ) ;
  assign n1541 = n1536 | n1540 ;
  assign n1542 = ( ~n1469 & n1471 ) | ( ~n1469 & n1541 ) | ( n1471 & n1541 ) ;
  assign n1543 = ( n1401 & ~n1415 ) | ( n1401 & n1417 ) | ( ~n1415 & n1417 ) ;
  assign n1544 = ( ~n1401 & n1418 ) | ( ~n1401 & n1543 ) | ( n1418 & n1543 ) ;
  assign n1545 = ( ~n1446 & n1542 ) | ( ~n1446 & n1544 ) | ( n1542 & n1544 ) ;
  assign n1546 = ~n1422 & n1545 ;
  assign n1547 = n1421 | n1546 ;
  assign n1548 = ( n1371 & ~n1399 ) | ( n1371 & n1547 ) | ( ~n1399 & n1547 ) ;
  assign n1549 = ( n1340 & ~n1342 ) | ( n1340 & n1344 ) | ( ~n1342 & n1344 ) ;
  assign n1550 = ( ~n1340 & n1345 ) | ( ~n1340 & n1549 ) | ( n1345 & n1549 ) ;
  assign n1551 = ( ~n1369 & n1548 ) | ( ~n1369 & n1550 ) | ( n1548 & n1550 ) ;
  assign n1552 = ( n1306 & ~n1345 ) | ( n1306 & n1551 ) | ( ~n1345 & n1551 ) ;
  assign n1553 = ( n1242 & n1244 ) | ( n1242 & n1283 ) | ( n1244 & n1283 ) ;
  assign n1554 = ( n1242 & n1284 ) | ( n1242 & ~n1553 ) | ( n1284 & ~n1553 ) ;
  assign n1555 = ( ~n1304 & n1552 ) | ( ~n1304 & n1554 ) | ( n1552 & n1554 ) ;
  assign n1556 = ( n1240 & ~n1284 ) | ( n1240 & n1555 ) | ( ~n1284 & n1555 ) ;
  assign n1557 = ( n1070 & n1099 ) | ( n1070 & n1143 ) | ( n1099 & n1143 ) ;
  assign n1558 = ( n1070 & n1144 ) | ( n1070 & ~n1557 ) | ( n1144 & ~n1557 ) ;
  assign n1559 = ( ~n1238 & n1556 ) | ( ~n1238 & n1558 ) | ( n1556 & n1558 ) ;
  assign n1560 = ( n1063 & n1065 ) | ( n1063 & ~n1067 ) | ( n1065 & ~n1067 ) ;
  assign n1561 = ( ~n1063 & n1068 ) | ( ~n1063 & n1560 ) | ( n1068 & n1560 ) ;
  assign n1562 = ( ~n1144 & n1559 ) | ( ~n1144 & n1561 ) | ( n1559 & n1561 ) ;
  assign n1563 = ( n1029 & ~n1031 ) | ( n1029 & n1033 ) | ( ~n1031 & n1033 ) ;
  assign n1564 = ( ~n1029 & n1034 ) | ( ~n1029 & n1563 ) | ( n1034 & n1563 ) ;
  assign n1565 = ( ~n1068 & n1562 ) | ( ~n1068 & n1564 ) | ( n1562 & n1564 ) ;
  assign n1566 = ( ~n1034 & n1036 ) | ( ~n1034 & n1565 ) | ( n1036 & n1565 ) ;
  assign n1567 = ( n790 & ~n914 ) | ( n790 & n1566 ) | ( ~n914 & n1566 ) ;
  assign n1568 = n640 & n1077 ;
  assign n1569 = n586 | n1568 ;
  assign n1570 = ~n655 & n664 ;
  assign n1571 = n584 & n603 ;
  assign n1572 = n1570 | n1571 ;
  assign n1573 = ( n649 & ~n1569 ) | ( n649 & n1572 ) | ( ~n1569 & n1572 ) ;
  assign n1574 = ( n649 & n1569 ) | ( n649 & ~n1572 ) | ( n1569 & ~n1572 ) ;
  assign n1575 = ( ~n649 & n1573 ) | ( ~n649 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1576 = ( ~n788 & n1567 ) | ( ~n788 & n1575 ) | ( n1567 & n1575 ) ;
  assign n1577 = n584 & n606 ;
  assign n1578 = n640 & n1577 ;
  assign n1579 = ~n1576 & n1578 ;
  assign n1580 = n173 | n373 ;
  assign n1581 = n1011 | n1580 ;
  assign n1582 = n165 | n331 ;
  assign n1583 = n495 | n1582 ;
  assign n1584 = n252 | n728 ;
  assign n1585 = n188 | n1584 ;
  assign n1586 = n1583 | n1585 ;
  assign n1587 = n296 | n1586 ;
  assign n1588 = n1581 | n1587 ;
  assign n1589 = n379 | n626 ;
  assign n1590 = n180 | n522 ;
  assign n1591 = n1589 | n1590 ;
  assign n1592 = n575 | n1591 ;
  assign n1593 = n240 | n534 ;
  assign n1594 = n193 | n710 ;
  assign n1595 = n391 | n1594 ;
  assign n1596 = n1593 | n1595 ;
  assign n1597 = n1592 | n1596 ;
  assign n1598 = n211 | n546 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = ~n828 & n977 ;
  assign n1601 = ~n949 & n1600 ;
  assign n1602 = ~n1599 & n1601 ;
  assign n1603 = ~n1588 & n1602 ;
  assign n1604 = n584 & n591 ;
  assign n1605 = ( n38 & n584 ) | ( n38 & n606 ) | ( n584 & n606 ) ;
  assign n1606 = ~n1577 & n1605 ;
  assign n1607 = ( n640 & ~n1075 ) | ( n640 & n1606 ) | ( ~n1075 & n1606 ) ;
  assign n1608 = ~n1075 & n1606 ;
  assign n1609 = ( n1604 & n1607 ) | ( n1604 & ~n1608 ) | ( n1607 & ~n1608 ) ;
  assign n1610 = ( ~n1573 & n1576 ) | ( ~n1573 & n1609 ) | ( n1576 & n1609 ) ;
  assign n1611 = ( n1573 & n1576 ) | ( n1573 & ~n1609 ) | ( n1576 & ~n1609 ) ;
  assign n1612 = ( ~n1576 & n1610 ) | ( ~n1576 & n1611 ) | ( n1610 & n1611 ) ;
  assign n1613 = n400 | n710 ;
  assign n1614 = n254 | n1613 ;
  assign n1615 = n479 | n1614 ;
  assign n1616 = n313 | n1615 ;
  assign n1617 = n239 | n957 ;
  assign n1618 = n669 | n719 ;
  assign n1619 = n1617 | n1618 ;
  assign n1620 = n456 | n1619 ;
  assign n1621 = n1616 | n1620 ;
  assign n1622 = n136 | n199 ;
  assign n1623 = n149 | n594 ;
  assign n1624 = n1622 | n1623 ;
  assign n1625 = n731 | n846 ;
  assign n1626 = n1624 | n1625 ;
  assign n1627 = n242 | n408 ;
  assign n1628 = n116 | n1627 ;
  assign n1629 = n690 | n1628 ;
  assign n1630 = n1626 | n1629 ;
  assign n1631 = n171 | n439 ;
  assign n1632 = n626 | n1631 ;
  assign n1633 = n419 | n1632 ;
  assign n1634 = n209 | n261 ;
  assign n1635 = n176 | n371 ;
  assign n1636 = n1634 | n1635 ;
  assign n1637 = n1633 | n1636 ;
  assign n1638 = n69 | n278 ;
  assign n1639 = n405 | n1638 ;
  assign n1640 = n290 | n505 ;
  assign n1641 = n1639 | n1640 ;
  assign n1642 = n198 | n282 ;
  assign n1643 = n56 & n148 ;
  assign n1644 = n159 | n1643 ;
  assign n1645 = n1642 | n1644 ;
  assign n1646 = n179 | n421 ;
  assign n1647 = n545 | n1646 ;
  assign n1648 = n1645 | n1647 ;
  assign n1649 = n1641 | n1648 ;
  assign n1650 = n1637 | n1649 ;
  assign n1651 = n1630 | n1650 ;
  assign n1652 = n1621 | n1651 ;
  assign n1653 = ( n788 & n1567 ) | ( n788 & n1575 ) | ( n1567 & n1575 ) ;
  assign n1654 = ( n788 & n1576 ) | ( n788 & ~n1653 ) | ( n1576 & ~n1653 ) ;
  assign n1655 = n87 | n199 ;
  assign n1656 = n121 | n145 ;
  assign n1657 = n478 | n1656 ;
  assign n1658 = n1655 | n1657 ;
  assign n1659 = n681 | n1658 ;
  assign n1660 = n879 | n1659 ;
  assign n1661 = n377 | n1660 ;
  assign n1662 = n463 | n832 ;
  assign n1663 = n824 | n1662 ;
  assign n1664 = n734 | n1663 ;
  assign n1665 = n968 | n1664 ;
  assign n1666 = n1661 | n1665 ;
  assign n1667 = ( n790 & n914 ) | ( n790 & ~n1566 ) | ( n914 & ~n1566 ) ;
  assign n1668 = ( ~n790 & n1567 ) | ( ~n790 & n1667 ) | ( n1567 & n1667 ) ;
  assign n1669 = n181 | n531 ;
  assign n1670 = n296 | n1633 ;
  assign n1671 = n268 | n469 ;
  assign n1672 = n197 | n1671 ;
  assign n1673 = n1614 | n1672 ;
  assign n1674 = n145 | n424 ;
  assign n1675 = n336 | n420 ;
  assign n1676 = n1674 | n1675 ;
  assign n1677 = n130 | n482 ;
  assign n1678 = n415 | n1677 ;
  assign n1679 = n1676 | n1678 ;
  assign n1680 = n1673 | n1679 ;
  assign n1681 = n1670 | n1680 ;
  assign n1682 = n1669 | n1681 ;
  assign n1683 = n127 | n150 ;
  assign n1684 = n679 | n1683 ;
  assign n1685 = n382 | n1684 ;
  assign n1686 = n70 | n190 ;
  assign n1687 = n421 | n485 ;
  assign n1688 = n1686 | n1687 ;
  assign n1689 = n831 | n1688 ;
  assign n1690 = n305 | n1689 ;
  assign n1691 = n1685 | n1690 ;
  assign n1692 = n102 | n312 ;
  assign n1693 = n179 | n1692 ;
  assign n1694 = n315 | n368 ;
  assign n1695 = n970 | n1694 ;
  assign n1696 = n1693 | n1695 ;
  assign n1697 = n240 | n407 ;
  assign n1698 = n1696 | n1697 ;
  assign n1699 = n289 | n1698 ;
  assign n1700 = n1691 | n1699 ;
  assign n1701 = n1682 | n1700 ;
  assign n1702 = n162 | n241 ;
  assign n1703 = n371 | n1702 ;
  assign n1704 = n1681 | n1703 ;
  assign n1705 = n154 | n277 ;
  assign n1706 = n450 | n1705 ;
  assign n1707 = ~n686 & n977 ;
  assign n1708 = ~n89 & n1707 ;
  assign n1709 = ~n1706 & n1708 ;
  assign n1710 = n278 | n321 ;
  assign n1711 = n534 | n1710 ;
  assign n1712 = n1709 & ~n1711 ;
  assign n1713 = n173 | n975 ;
  assign n1714 = n206 | n1713 ;
  assign n1715 = n137 | n263 ;
  assign n1716 = n454 | n1715 ;
  assign n1717 = n572 | n1694 ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = n1714 | n1718 ;
  assign n1720 = n1626 | n1719 ;
  assign n1721 = n1712 & ~n1720 ;
  assign n1722 = ~n1704 & n1721 ;
  assign n1723 = n87 | n362 ;
  assign n1724 = n161 | n420 ;
  assign n1725 = n1723 | n1724 ;
  assign n1726 = n114 | n279 ;
  assign n1727 = n348 | n1726 ;
  assign n1728 = n1725 | n1727 ;
  assign n1729 = n92 | n355 ;
  assign n1730 = n312 | n1729 ;
  assign n1731 = n835 | n1730 ;
  assign n1732 = n1728 | n1731 ;
  assign n1733 = n424 | n719 ;
  assign n1734 = n1593 | n1733 ;
  assign n1735 = n1639 | n1734 ;
  assign n1736 = n153 | n1735 ;
  assign n1737 = n1732 | n1736 ;
  assign n1738 = n1588 | n1737 ;
  assign n1739 = n139 & n458 ;
  assign n1740 = n1738 | n1739 ;
  assign n1741 = n146 | n300 ;
  assign n1742 = n259 | n268 ;
  assign n1743 = n1741 | n1742 ;
  assign n1744 = n408 | n624 ;
  assign n1745 = n1743 | n1744 ;
  assign n1746 = n455 | n1745 ;
  assign n1747 = n42 & n52 ;
  assign n1748 = n86 & n1747 ;
  assign n1749 = n312 | n1748 ;
  assign n1750 = n163 | n1749 ;
  assign n1751 = n194 | n1750 ;
  assign n1752 = n179 | n290 ;
  assign n1753 = n258 | n1634 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1751 | n1754 ;
  assign n1756 = n1746 | n1755 ;
  assign n1757 = n57 & n174 ;
  assign n1758 = n360 | n1757 ;
  assign n1759 = n338 | n1758 ;
  assign n1760 = n969 | n1759 ;
  assign n1761 = n568 | n632 ;
  assign n1762 = n1669 | n1761 ;
  assign n1763 = n1760 | n1762 ;
  assign n1764 = n685 | n1763 ;
  assign n1765 = n1756 | n1764 ;
  assign n1766 = n373 | n463 ;
  assign n1767 = n89 | n441 ;
  assign n1768 = n1766 | n1767 ;
  assign n1769 = n404 | n505 ;
  assign n1770 = n522 | n1769 ;
  assign n1771 = n596 | n1770 ;
  assign n1772 = n163 | n445 ;
  assign n1773 = n1771 | n1772 ;
  assign n1774 = n1768 | n1773 ;
  assign n1775 = n203 | n538 ;
  assign n1776 = n102 | n485 ;
  assign n1777 = n1775 | n1776 ;
  assign n1778 = n263 | n405 ;
  assign n1779 = n889 | n1778 ;
  assign n1780 = n1777 | n1779 ;
  assign n1781 = n1774 | n1780 ;
  assign n1782 = n283 | n311 ;
  assign n1783 = n178 | n1782 ;
  assign n1784 = n453 | n1783 ;
  assign n1785 = n287 | n419 ;
  assign n1786 = n1184 | n1785 ;
  assign n1787 = n743 | n1786 ;
  assign n1788 = n1745 | n1787 ;
  assign n1789 = n1784 | n1788 ;
  assign n1790 = ~n256 & n1600 ;
  assign n1791 = ~n1789 & n1790 ;
  assign n1792 = ~n1781 & n1791 ;
  assign n1793 = n692 | n964 ;
  assign n1794 = n1766 | n1793 ;
  assign n1795 = n291 | n852 ;
  assign n1796 = n334 | n383 ;
  assign n1797 = n1795 | n1796 ;
  assign n1798 = n681 | n1797 ;
  assign n1799 = n815 | n1798 ;
  assign n1800 = n1794 | n1799 ;
  assign n1801 = n1763 | n1800 ;
  assign n1802 = n1621 | n1801 ;
  assign n1803 = ( n1369 & n1548 ) | ( n1369 & ~n1550 ) | ( n1548 & ~n1550 ) ;
  assign n1804 = ( ~n1548 & n1551 ) | ( ~n1548 & n1803 ) | ( n1551 & n1803 ) ;
  assign n1805 = ~n1802 & n1804 ;
  assign n1806 = n119 | n422 ;
  assign n1807 = n530 | n594 ;
  assign n1808 = n291 | n1807 ;
  assign n1809 = n1806 | n1808 ;
  assign n1810 = n96 | n287 ;
  assign n1811 = n163 | n1589 ;
  assign n1812 = n1810 | n1811 ;
  assign n1813 = n147 | n754 ;
  assign n1814 = n1812 | n1813 ;
  assign n1815 = n1809 | n1814 ;
  assign n1816 = n845 | n1758 ;
  assign n1817 = n816 | n1816 ;
  assign n1818 = n298 | n319 ;
  assign n1819 = n713 | n1818 ;
  assign n1820 = n1817 | n1819 ;
  assign n1821 = n165 | n245 ;
  assign n1822 = n140 | n400 ;
  assign n1823 = n321 | n1822 ;
  assign n1824 = n1821 | n1823 ;
  assign n1825 = n136 | n209 ;
  assign n1826 = n272 | n1825 ;
  assign n1827 = n68 & n106 ;
  assign n1828 = n312 | n1827 ;
  assign n1829 = n1826 | n1828 ;
  assign n1830 = n74 & ~n78 ;
  assign n1831 = n199 | n1830 ;
  assign n1832 = n263 | n267 ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = n1829 | n1833 ;
  assign n1835 = n1824 | n1834 ;
  assign n1836 = n1820 | n1835 ;
  assign n1837 = n1815 | n1836 ;
  assign n1838 = ( ~n1306 & n1345 ) | ( ~n1306 & n1551 ) | ( n1345 & n1551 ) ;
  assign n1839 = ( ~n1551 & n1552 ) | ( ~n1551 & n1838 ) | ( n1552 & n1838 ) ;
  assign n1840 = ( n1805 & ~n1837 ) | ( n1805 & n1839 ) | ( ~n1837 & n1839 ) ;
  assign n1841 = ( n1304 & n1552 ) | ( n1304 & ~n1554 ) | ( n1552 & ~n1554 ) ;
  assign n1842 = ( ~n1552 & n1555 ) | ( ~n1552 & n1841 ) | ( n1555 & n1841 ) ;
  assign n1843 = ( n1792 & n1840 ) | ( n1792 & n1842 ) | ( n1840 & n1842 ) ;
  assign n1844 = ( ~n1240 & n1284 ) | ( ~n1240 & n1555 ) | ( n1284 & n1555 ) ;
  assign n1845 = ( ~n1555 & n1556 ) | ( ~n1555 & n1844 ) | ( n1556 & n1844 ) ;
  assign n1846 = ( ~n1765 & n1843 ) | ( ~n1765 & n1845 ) | ( n1843 & n1845 ) ;
  assign n1847 = ( n1238 & n1556 ) | ( n1238 & ~n1558 ) | ( n1556 & ~n1558 ) ;
  assign n1848 = ( ~n1556 & n1559 ) | ( ~n1556 & n1847 ) | ( n1559 & n1847 ) ;
  assign n1849 = ( ~n1740 & n1846 ) | ( ~n1740 & n1848 ) | ( n1846 & n1848 ) ;
  assign n1850 = n329 | n682 ;
  assign n1851 = n612 | n675 ;
  assign n1852 = n1850 | n1851 ;
  assign n1853 = n458 | n1852 ;
  assign n1854 = n293 | n391 ;
  assign n1855 = n241 | n363 ;
  assign n1856 = n1854 | n1855 ;
  assign n1857 = n1820 | n1856 ;
  assign n1858 = n188 | n397 ;
  assign n1859 = n951 | n1858 ;
  assign n1860 = n842 | n1859 ;
  assign n1861 = n1771 | n1860 ;
  assign n1862 = n1857 | n1861 ;
  assign n1863 = n1853 | n1862 ;
  assign n1864 = ( n1144 & n1559 ) | ( n1144 & n1561 ) | ( n1559 & n1561 ) ;
  assign n1865 = ( n1144 & n1562 ) | ( n1144 & ~n1864 ) | ( n1562 & ~n1864 ) ;
  assign n1866 = ( n1849 & ~n1863 ) | ( n1849 & n1865 ) | ( ~n1863 & n1865 ) ;
  assign n1867 = n360 | n372 ;
  assign n1868 = n838 | n1867 ;
  assign n1869 = n354 | n362 ;
  assign n1870 = n259 | n419 ;
  assign n1871 = n1869 | n1870 ;
  assign n1872 = n261 | n298 ;
  assign n1873 = ( ~n42 & n52 ) | ( ~n42 & n189 ) | ( n52 & n189 ) ;
  assign n1874 = ( n188 & n189 ) | ( n188 & ~n1873 ) | ( n189 & ~n1873 ) ;
  assign n1875 = n1872 | n1874 ;
  assign n1876 = n572 | n843 ;
  assign n1877 = n1875 | n1876 ;
  assign n1878 = n1871 | n1877 ;
  assign n1879 = n133 | n1878 ;
  assign n1880 = n1163 | n1879 ;
  assign n1881 = n1868 | n1880 ;
  assign n1882 = ( n1068 & n1562 ) | ( n1068 & ~n1564 ) | ( n1562 & ~n1564 ) ;
  assign n1883 = ( ~n1562 & n1565 ) | ( ~n1562 & n1882 ) | ( n1565 & n1882 ) ;
  assign n1884 = ( n1866 & ~n1881 ) | ( n1866 & n1883 ) | ( ~n1881 & n1883 ) ;
  assign n1885 = ( n1034 & ~n1036 ) | ( n1034 & n1565 ) | ( ~n1036 & n1565 ) ;
  assign n1886 = ( ~n1565 & n1566 ) | ( ~n1565 & n1885 ) | ( n1566 & n1885 ) ;
  assign n1887 = ( n1722 & n1884 ) | ( n1722 & n1886 ) | ( n1884 & n1886 ) ;
  assign n1888 = ( n1668 & ~n1701 ) | ( n1668 & n1887 ) | ( ~n1701 & n1887 ) ;
  assign n1889 = ( n1654 & ~n1666 ) | ( n1654 & n1888 ) | ( ~n1666 & n1888 ) ;
  assign n1890 = ( n1612 & ~n1652 ) | ( n1612 & n1889 ) | ( ~n1652 & n1889 ) ;
  assign n1891 = ( n1579 & n1603 ) | ( n1579 & n1890 ) | ( n1603 & n1890 ) ;
  assign n1892 = ( ~n1579 & n1603 ) | ( ~n1579 & n1890 ) | ( n1603 & n1890 ) ;
  assign n1893 = ( n1579 & ~n1891 ) | ( n1579 & n1892 ) | ( ~n1891 & n1892 ) ;
  assign n1894 = ( n1668 & n1701 ) | ( n1668 & ~n1887 ) | ( n1701 & ~n1887 ) ;
  assign n1895 = ( ~n1668 & n1888 ) | ( ~n1668 & n1894 ) | ( n1888 & n1894 ) ;
  assign n1896 = ( n1866 & n1881 ) | ( n1866 & ~n1883 ) | ( n1881 & ~n1883 ) ;
  assign n1897 = ( ~n1866 & n1884 ) | ( ~n1866 & n1896 ) | ( n1884 & n1896 ) ;
  assign n1898 = ( n1849 & n1863 ) | ( n1849 & ~n1865 ) | ( n1863 & ~n1865 ) ;
  assign n1899 = ( ~n1849 & n1866 ) | ( ~n1849 & n1898 ) | ( n1866 & n1898 ) ;
  assign n1900 = ( ~n1792 & n1840 ) | ( ~n1792 & n1842 ) | ( n1840 & n1842 ) ;
  assign n1901 = ( n1792 & ~n1843 ) | ( n1792 & n1900 ) | ( ~n1843 & n1900 ) ;
  assign n1902 = ( n1805 & n1837 ) | ( n1805 & ~n1839 ) | ( n1837 & ~n1839 ) ;
  assign n1903 = ( ~n1805 & n1840 ) | ( ~n1805 & n1902 ) | ( n1840 & n1902 ) ;
  assign n1904 = ~n1901 & n1903 ;
  assign n1905 = ( n1765 & n1843 ) | ( n1765 & ~n1845 ) | ( n1843 & ~n1845 ) ;
  assign n1906 = ( ~n1843 & n1846 ) | ( ~n1843 & n1905 ) | ( n1846 & n1905 ) ;
  assign n1907 = n1904 | n1906 ;
  assign n1908 = ( n1740 & ~n1846 ) | ( n1740 & n1848 ) | ( ~n1846 & n1848 ) ;
  assign n1909 = ( ~n1848 & n1849 ) | ( ~n1848 & n1908 ) | ( n1849 & n1908 ) ;
  assign n1910 = n1907 & n1909 ;
  assign n1911 = n1899 | n1910 ;
  assign n1912 = n1897 & n1911 ;
  assign n1913 = ( n1722 & n1884 ) | ( n1722 & ~n1886 ) | ( n1884 & ~n1886 ) ;
  assign n1914 = ( n1886 & ~n1887 ) | ( n1886 & n1913 ) | ( ~n1887 & n1913 ) ;
  assign n1915 = ~n1912 & n1914 ;
  assign n1916 = n1895 & ~n1915 ;
  assign n1917 = ( n1654 & n1666 ) | ( n1654 & ~n1888 ) | ( n1666 & ~n1888 ) ;
  assign n1918 = ( ~n1654 & n1889 ) | ( ~n1654 & n1917 ) | ( n1889 & n1917 ) ;
  assign n1919 = n1916 | n1918 ;
  assign n1920 = ( n1612 & n1652 ) | ( n1612 & ~n1889 ) | ( n1652 & ~n1889 ) ;
  assign n1921 = ( ~n1612 & n1890 ) | ( ~n1612 & n1920 ) | ( n1890 & n1920 ) ;
  assign n1922 = n1919 & n1921 ;
  assign n1923 = n1893 & n1922 ;
  assign n1924 = n1802 & ~n1804 ;
  assign n1925 = n1805 | n1924 ;
  assign n1926 = n1903 & n1925 ;
  assign n1927 = n1901 & ~n1926 ;
  assign n1928 = n1906 & ~n1927 ;
  assign n1929 = n1909 | n1928 ;
  assign n1930 = n1899 & n1929 ;
  assign n1931 = n1897 | n1930 ;
  assign n1932 = ~n1914 & n1931 ;
  assign n1933 = n1895 | n1932 ;
  assign n1934 = n1918 & n1933 ;
  assign n1935 = n1921 | n1934 ;
  assign n1936 = ( n1893 & ~n1922 ) | ( n1893 & n1935 ) | ( ~n1922 & n1935 ) ;
  assign n1937 = n1893 & n1935 ;
  assign n1938 = ( n1923 & n1936 ) | ( n1923 & ~n1937 ) | ( n1936 & ~n1937 ) ;
  assign n1939 = n225 & n236 ;
  assign n1940 = ( n28 & ~n222 ) | ( n28 & n235 ) | ( ~n222 & n235 ) ;
  assign n1941 = ( n228 & n1939 ) | ( n228 & ~n1940 ) | ( n1939 & ~n1940 ) ;
  assign n1942 = n1918 & n1941 ;
  assign n1943 = ( n225 & n236 ) | ( n225 & ~n237 ) | ( n236 & ~n237 ) ;
  assign n1944 = ~n1939 & n1943 ;
  assign n1945 = n1921 & n1944 ;
  assign n1946 = n1942 | n1945 ;
  assign n1947 = ~n228 & n237 ;
  assign n1948 = ~n1893 & n1947 ;
  assign n1949 = n1946 | n1948 ;
  assign n1950 = ( n238 & ~n1938 ) | ( n238 & n1949 ) | ( ~n1938 & n1949 ) ;
  assign n1951 = n222 | n1949 ;
  assign n1952 = ~n1950 & n1951 ;
  assign n1953 = ( ~n1949 & n1950 ) | ( ~n1949 & n1951 ) | ( n1950 & n1951 ) ;
  assign n1954 = ( ~n222 & n1952 ) | ( ~n222 & n1953 ) | ( n1952 & n1953 ) ;
  assign n1955 = ~n1919 & n1921 ;
  assign n1956 = ( n1919 & n1921 ) | ( n1919 & ~n1934 ) | ( n1921 & ~n1934 ) ;
  assign n1957 = n1921 & ~n1934 ;
  assign n1958 = ( n1955 & n1956 ) | ( n1955 & ~n1957 ) | ( n1956 & ~n1957 ) ;
  assign n1959 = n1895 & n1941 ;
  assign n1960 = n1918 & n1944 ;
  assign n1961 = n1959 | n1960 ;
  assign n1962 = n1921 & n1947 ;
  assign n1963 = n1961 | n1962 ;
  assign n1964 = ( n238 & n1958 ) | ( n238 & n1963 ) | ( n1958 & n1963 ) ;
  assign n1965 = n222 & ~n1963 ;
  assign n1966 = n1964 | n1965 ;
  assign n1967 = ( n1963 & ~n1964 ) | ( n1963 & n1965 ) | ( ~n1964 & n1965 ) ;
  assign n1968 = ( ~n222 & n1966 ) | ( ~n222 & n1967 ) | ( n1966 & n1967 ) ;
  assign n1969 = n1916 & n1918 ;
  assign n1970 = ( ~n1916 & n1918 ) | ( ~n1916 & n1933 ) | ( n1918 & n1933 ) ;
  assign n1971 = ( ~n1934 & n1969 ) | ( ~n1934 & n1970 ) | ( n1969 & n1970 ) ;
  assign n1972 = ~n1914 & n1941 ;
  assign n1973 = n1895 & n1944 ;
  assign n1974 = n1972 | n1973 ;
  assign n1975 = n1918 & n1947 ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = ( n238 & n1971 ) | ( n238 & n1976 ) | ( n1971 & n1976 ) ;
  assign n1978 = n222 & ~n1976 ;
  assign n1979 = n1977 | n1978 ;
  assign n1980 = ( n1976 & ~n1977 ) | ( n1976 & n1978 ) | ( ~n1977 & n1978 ) ;
  assign n1981 = ( ~n222 & n1979 ) | ( ~n222 & n1980 ) | ( n1979 & n1980 ) ;
  assign n1982 = x7 & x8 ;
  assign n1983 = x7 | x8 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = n1276 & n1984 ;
  assign n1986 = n1897 | n1911 ;
  assign n1987 = ( n1897 & ~n1911 ) | ( n1897 & n1930 ) | ( ~n1911 & n1930 ) ;
  assign n1988 = ( ~n1931 & n1986 ) | ( ~n1931 & n1987 ) | ( n1986 & n1987 ) ;
  assign n1989 = n812 & n1275 ;
  assign n1990 = n812 | n1274 ;
  assign n1991 = ( n1984 & n1989 ) | ( n1984 & ~n1990 ) | ( n1989 & ~n1990 ) ;
  assign n1992 = n1909 & n1991 ;
  assign n1993 = ( n812 & n1275 ) | ( n812 & ~n1276 ) | ( n1275 & ~n1276 ) ;
  assign n1994 = ~n1989 & n1993 ;
  assign n1995 = n1899 & n1994 ;
  assign n1996 = n1992 | n1995 ;
  assign n1997 = n1276 & ~n1984 ;
  assign n1998 = n1897 & n1997 ;
  assign n1999 = n1996 | n1998 ;
  assign n2000 = ( n1985 & n1988 ) | ( n1985 & n1999 ) | ( n1988 & n1999 ) ;
  assign n2001 = n902 | n1999 ;
  assign n2002 = ~n2000 & n2001 ;
  assign n2003 = ( ~n1999 & n2000 ) | ( ~n1999 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2004 = ( ~n902 & n2002 ) | ( ~n902 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2005 = n1077 & n1925 ;
  assign n2006 = ~n770 & n902 ;
  assign n2007 = n770 & ~n902 ;
  assign n2008 = n2006 | n2007 ;
  assign n2009 = n646 & ~n783 ;
  assign n2010 = ~n646 & n783 ;
  assign n2011 = ( n2008 & n2009 ) | ( n2008 & n2010 ) | ( n2009 & n2010 ) ;
  assign n2012 = n2008 & ~n2011 ;
  assign n2013 = n1906 & n2012 ;
  assign n2014 = n2011 | n2013 ;
  assign n2015 = ( n1904 & ~n1906 ) | ( n1904 & n1927 ) | ( ~n1906 & n1927 ) ;
  assign n2016 = ~n1904 & n1928 ;
  assign n2017 = n2015 | n2016 ;
  assign n2018 = ( n2013 & n2014 ) | ( n2013 & ~n2017 ) | ( n2014 & ~n2017 ) ;
  assign n2019 = ~n646 & n902 ;
  assign n2020 = ( n770 & n783 ) | ( n770 & ~n902 ) | ( n783 & ~n902 ) ;
  assign n2021 = n646 | n2020 ;
  assign n2022 = n902 | n2020 ;
  assign n2023 = ( n2019 & n2021 ) | ( n2019 & ~n2022 ) | ( n2021 & ~n2022 ) ;
  assign n2024 = n1903 & n2023 ;
  assign n2025 = ~n2008 & n2022 ;
  assign n2026 = ~n785 & n2025 ;
  assign n2027 = ~n1901 & n2026 ;
  assign n2028 = n2024 | n2027 ;
  assign n2029 = n2018 | n2028 ;
  assign n2030 = n1903 & n2026 ;
  assign n2031 = ~n1901 & n2012 ;
  assign n2032 = n2030 | n2031 ;
  assign n2033 = n1903 & ~n1925 ;
  assign n2034 = n1901 & ~n2033 ;
  assign n2035 = ~n1901 & n2033 ;
  assign n2036 = n2034 | n2035 ;
  assign n2037 = n1925 & n2023 ;
  assign n2038 = n2011 | n2037 ;
  assign n2039 = ( ~n2036 & n2037 ) | ( ~n2036 & n2038 ) | ( n2037 & n2038 ) ;
  assign n2040 = n2032 | n2039 ;
  assign n2041 = n1903 | n1925 ;
  assign n2042 = ~n1926 & n2041 ;
  assign n2043 = n1925 & n2026 ;
  assign n2044 = n2011 | n2043 ;
  assign n2045 = ( n2042 & n2043 ) | ( n2042 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2046 = n1903 & n2012 ;
  assign n2047 = n2045 | n2046 ;
  assign n2048 = n1925 & n2008 ;
  assign n2049 = n646 & n2048 ;
  assign n2050 = ( n646 & n2047 ) | ( n646 & n2049 ) | ( n2047 & n2049 ) ;
  assign n2051 = n2040 | n2050 ;
  assign n2052 = n646 & n2051 ;
  assign n2053 = ( n2005 & n2029 ) | ( n2005 & ~n2052 ) | ( n2029 & ~n2052 ) ;
  assign n2054 = ( n2005 & ~n2029 ) | ( n2005 & n2052 ) | ( ~n2029 & n2052 ) ;
  assign n2055 = ( ~n2005 & n2053 ) | ( ~n2005 & n2054 ) | ( n2053 & n2054 ) ;
  assign n2056 = n1899 & n1910 ;
  assign n2057 = ( n1899 & ~n1910 ) | ( n1899 & n1929 ) | ( ~n1910 & n1929 ) ;
  assign n2058 = ( ~n1930 & n2056 ) | ( ~n1930 & n2057 ) | ( n2056 & n2057 ) ;
  assign n2059 = n1906 & n1991 ;
  assign n2060 = n1909 & n1994 ;
  assign n2061 = n2059 | n2060 ;
  assign n2062 = n1899 & n1997 ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = ( n1985 & n2058 ) | ( n1985 & n2063 ) | ( n2058 & n2063 ) ;
  assign n2065 = n902 & ~n2063 ;
  assign n2066 = n2064 | n2065 ;
  assign n2067 = ( n2063 & ~n2064 ) | ( n2063 & n2065 ) | ( ~n2064 & n2065 ) ;
  assign n2068 = ( ~n902 & n2066 ) | ( ~n902 & n2067 ) | ( n2066 & n2067 ) ;
  assign n2069 = n2040 & n2050 ;
  assign n2070 = n2051 & ~n2069 ;
  assign n2071 = ( ~n1909 & n1927 ) | ( ~n1909 & n2015 ) | ( n1927 & n2015 ) ;
  assign n2072 = ( n1909 & n1927 ) | ( n1909 & n2015 ) | ( n1927 & n2015 ) ;
  assign n2073 = ( n1909 & n2071 ) | ( n1909 & ~n2072 ) | ( n2071 & ~n2072 ) ;
  assign n2074 = ~n1901 & n1991 ;
  assign n2075 = n1906 & n1994 ;
  assign n2076 = n2074 | n2075 ;
  assign n2077 = n1909 & n1997 ;
  assign n2078 = n2076 | n2077 ;
  assign n2079 = ( n1985 & n2073 ) | ( n1985 & n2078 ) | ( n2073 & n2078 ) ;
  assign n2080 = n902 & ~n2078 ;
  assign n2081 = n2079 | n2080 ;
  assign n2082 = ( n2078 & ~n2079 ) | ( n2078 & n2080 ) | ( ~n2079 & n2080 ) ;
  assign n2083 = ( ~n902 & n2081 ) | ( ~n902 & n2082 ) | ( n2081 & n2082 ) ;
  assign n2084 = ~n2047 & n2049 ;
  assign n2085 = n2047 & ~n2049 ;
  assign n2086 = n2084 | n2085 ;
  assign n2087 = n1903 & n1991 ;
  assign n2088 = ~n1901 & n1994 ;
  assign n2089 = n2087 | n2088 ;
  assign n2090 = n1906 & n1997 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = n1985 & ~n2017 ;
  assign n2093 = n2091 | n2092 ;
  assign n2094 = n1985 & ~n2036 ;
  assign n2095 = n1903 & n1994 ;
  assign n2096 = ~n1901 & n1997 ;
  assign n2097 = n2095 | n2096 ;
  assign n2098 = n1925 & n1991 ;
  assign n2099 = n2097 | n2098 ;
  assign n2100 = n2094 | n2099 ;
  assign n2101 = n1276 & n1925 ;
  assign n2102 = n1925 & n1994 ;
  assign n2103 = n1985 | n2102 ;
  assign n2104 = ( n2042 & n2102 ) | ( n2042 & n2103 ) | ( n2102 & n2103 ) ;
  assign n2105 = n1903 & n1997 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n2101 | n2106 ;
  assign n2108 = n2100 | n2107 ;
  assign n2109 = n902 & n2108 ;
  assign n2110 = ( n2048 & n2093 ) | ( n2048 & ~n2109 ) | ( n2093 & ~n2109 ) ;
  assign n2111 = ( n2048 & ~n2093 ) | ( n2048 & n2109 ) | ( ~n2093 & n2109 ) ;
  assign n2112 = ( ~n2048 & n2110 ) | ( ~n2048 & n2111 ) | ( n2110 & n2111 ) ;
  assign n2113 = n902 & ~n2108 ;
  assign n2114 = ( n2048 & ~n2112 ) | ( n2048 & n2113 ) | ( ~n2112 & n2113 ) ;
  assign n2115 = ( n2083 & n2086 ) | ( n2083 & n2114 ) | ( n2086 & n2114 ) ;
  assign n2116 = ( n2068 & n2070 ) | ( n2068 & n2115 ) | ( n2070 & n2115 ) ;
  assign n2117 = ( n2004 & n2055 ) | ( n2004 & n2116 ) | ( n2055 & n2116 ) ;
  assign n2118 = ( ~n2004 & n2055 ) | ( ~n2004 & n2116 ) | ( n2055 & n2116 ) ;
  assign n2119 = ( n2004 & ~n2117 ) | ( n2004 & n2118 ) | ( ~n2117 & n2118 ) ;
  assign n2120 = ~n1895 & n1915 ;
  assign n2121 = ( n1895 & n1915 ) | ( n1895 & n1932 ) | ( n1915 & n1932 ) ;
  assign n2122 = ( n1933 & n2120 ) | ( n1933 & ~n2121 ) | ( n2120 & ~n2121 ) ;
  assign n2123 = n1897 & n1941 ;
  assign n2124 = ~n1914 & n1944 ;
  assign n2125 = n2123 | n2124 ;
  assign n2126 = n1895 & n1947 ;
  assign n2127 = n2125 | n2126 ;
  assign n2128 = ( n238 & ~n2122 ) | ( n238 & n2127 ) | ( ~n2122 & n2127 ) ;
  assign n2129 = n222 | n2127 ;
  assign n2130 = ~n2128 & n2129 ;
  assign n2131 = ( ~n2127 & n2128 ) | ( ~n2127 & n2129 ) | ( n2128 & n2129 ) ;
  assign n2132 = ( ~n222 & n2130 ) | ( ~n222 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2133 = n1912 & n1914 ;
  assign n2134 = ( ~n1912 & n1914 ) | ( ~n1912 & n1931 ) | ( n1914 & n1931 ) ;
  assign n2135 = n1914 & n1931 ;
  assign n2136 = ( n2133 & n2134 ) | ( n2133 & ~n2135 ) | ( n2134 & ~n2135 ) ;
  assign n2137 = n1899 & n1941 ;
  assign n2138 = n1897 & n1944 ;
  assign n2139 = n2137 | n2138 ;
  assign n2140 = ~n1914 & n1947 ;
  assign n2141 = n2139 | n2140 ;
  assign n2142 = ( n238 & ~n2136 ) | ( n238 & n2141 ) | ( ~n2136 & n2141 ) ;
  assign n2143 = n222 | n2141 ;
  assign n2144 = ~n2142 & n2143 ;
  assign n2145 = ( ~n2141 & n2142 ) | ( ~n2141 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2146 = ( ~n222 & n2144 ) | ( ~n222 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2147 = n1909 & n1941 ;
  assign n2148 = n1899 & n1944 ;
  assign n2149 = n2147 | n2148 ;
  assign n2150 = n1897 & n1947 ;
  assign n2151 = n2149 | n2150 ;
  assign n2152 = ( n238 & n1988 ) | ( n238 & n2151 ) | ( n1988 & n2151 ) ;
  assign n2153 = n222 | n2151 ;
  assign n2154 = ~n2152 & n2153 ;
  assign n2155 = ( ~n2151 & n2152 ) | ( ~n2151 & n2153 ) | ( n2152 & n2153 ) ;
  assign n2156 = ( ~n222 & n2154 ) | ( ~n222 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = n1906 & n1941 ;
  assign n2158 = n1909 & n1944 ;
  assign n2159 = n2157 | n2158 ;
  assign n2160 = n1899 & n1947 ;
  assign n2161 = n2159 | n2160 ;
  assign n2162 = ( n238 & n2058 ) | ( n238 & n2161 ) | ( n2058 & n2161 ) ;
  assign n2163 = n222 & ~n2161 ;
  assign n2164 = n2162 | n2163 ;
  assign n2165 = ( n2161 & ~n2162 ) | ( n2161 & n2163 ) | ( ~n2162 & n2163 ) ;
  assign n2166 = ( ~n222 & n2164 ) | ( ~n222 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = ~n902 & n2100 ;
  assign n2168 = ( n902 & n2100 ) | ( n902 & n2107 ) | ( n2100 & n2107 ) ;
  assign n2169 = n2100 & n2107 ;
  assign n2170 = ( n2167 & n2168 ) | ( n2167 & ~n2169 ) | ( n2168 & ~n2169 ) ;
  assign n2171 = ~n1901 & n1941 ;
  assign n2172 = n1906 & n1944 ;
  assign n2173 = n2171 | n2172 ;
  assign n2174 = n1909 & n1947 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = ( n238 & n2073 ) | ( n238 & n2175 ) | ( n2073 & n2175 ) ;
  assign n2177 = n222 & ~n2175 ;
  assign n2178 = n2176 | n2177 ;
  assign n2179 = ( n2175 & ~n2176 ) | ( n2175 & n2177 ) | ( ~n2176 & n2177 ) ;
  assign n2180 = ( ~n222 & n2178 ) | ( ~n222 & n2179 ) | ( n2178 & n2179 ) ;
  assign n2181 = n902 & n2101 ;
  assign n2182 = ~n2106 & n2181 ;
  assign n2183 = n2106 & ~n2181 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = n1903 & n1941 ;
  assign n2186 = ~n1901 & n1944 ;
  assign n2187 = n2185 | n2186 ;
  assign n2188 = n1906 & n1947 ;
  assign n2189 = n2187 | n2188 ;
  assign n2190 = n238 & ~n2017 ;
  assign n2191 = n2189 | n2190 ;
  assign n2192 = n237 & n1925 ;
  assign n2193 = n222 & n2192 ;
  assign n2194 = n1903 & n1947 ;
  assign n2195 = n238 | n2194 ;
  assign n2196 = ( n2042 & n2194 ) | ( n2042 & n2195 ) | ( n2194 & n2195 ) ;
  assign n2197 = n1925 & n1944 ;
  assign n2198 = n2196 | n2197 ;
  assign n2199 = n2193 | n2198 ;
  assign n2200 = n238 & ~n2036 ;
  assign n2201 = n1903 & n1944 ;
  assign n2202 = ~n1901 & n1947 ;
  assign n2203 = n2201 | n2202 ;
  assign n2204 = n1925 & n1941 ;
  assign n2205 = n2203 | n2204 ;
  assign n2206 = n2200 | n2205 ;
  assign n2207 = ( n222 & n2199 ) | ( n222 & n2206 ) | ( n2199 & n2206 ) ;
  assign n2208 = ( n222 & n2193 ) | ( n222 & n2207 ) | ( n2193 & n2207 ) ;
  assign n2209 = ( n2101 & n2191 ) | ( n2101 & ~n2208 ) | ( n2191 & ~n2208 ) ;
  assign n2210 = ( n2101 & ~n2191 ) | ( n2101 & n2208 ) | ( ~n2191 & n2208 ) ;
  assign n2211 = ( ~n2101 & n2209 ) | ( ~n2101 & n2210 ) | ( n2209 & n2210 ) ;
  assign n2212 = n222 & ~n2207 ;
  assign n2213 = ( n2101 & ~n2211 ) | ( n2101 & n2212 ) | ( ~n2211 & n2212 ) ;
  assign n2214 = ( n2180 & n2184 ) | ( n2180 & n2213 ) | ( n2184 & n2213 ) ;
  assign n2215 = ( n2166 & n2170 ) | ( n2166 & n2214 ) | ( n2170 & n2214 ) ;
  assign n2216 = ( n2112 & n2156 ) | ( n2112 & n2215 ) | ( n2156 & n2215 ) ;
  assign n2217 = ( ~n2083 & n2086 ) | ( ~n2083 & n2114 ) | ( n2086 & n2114 ) ;
  assign n2218 = ( n2083 & ~n2115 ) | ( n2083 & n2217 ) | ( ~n2115 & n2217 ) ;
  assign n2219 = ( n2146 & n2216 ) | ( n2146 & n2218 ) | ( n2216 & n2218 ) ;
  assign n2220 = ( n2068 & ~n2070 ) | ( n2068 & n2115 ) | ( ~n2070 & n2115 ) ;
  assign n2221 = ( n2070 & ~n2116 ) | ( n2070 & n2220 ) | ( ~n2116 & n2220 ) ;
  assign n2222 = ( n2132 & n2219 ) | ( n2132 & n2221 ) | ( n2219 & n2221 ) ;
  assign n2223 = ( n1981 & n2119 ) | ( n1981 & n2222 ) | ( n2119 & n2222 ) ;
  assign n2224 = n2011 & n2073 ;
  assign n2225 = ~n1901 & n2023 ;
  assign n2226 = n1909 & n2012 ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = ( ~n646 & n2224 ) | ( ~n646 & n2227 ) | ( n2224 & n2227 ) ;
  assign n2229 = n1906 & n2026 ;
  assign n2230 = n646 & ~n2227 ;
  assign n2231 = n2229 | n2230 ;
  assign n2232 = ( n2224 & n2229 ) | ( n2224 & n2230 ) | ( n2229 & n2230 ) ;
  assign n2233 = ( n2228 & n2231 ) | ( n2228 & ~n2232 ) | ( n2231 & ~n2232 ) ;
  assign n2234 = n606 | n1075 ;
  assign n2235 = ( n606 & n1075 ) | ( n606 & n1077 ) | ( n1075 & n1077 ) ;
  assign n2236 = n2234 & ~n2235 ;
  assign n2237 = n1925 & n2236 ;
  assign n2238 = n1077 & n1606 ;
  assign n2239 = n2237 | n2238 ;
  assign n2240 = ( n2042 & n2237 ) | ( n2042 & n2239 ) | ( n2237 & n2239 ) ;
  assign n2241 = n1077 & ~n1606 ;
  assign n2242 = n1903 & n2241 ;
  assign n2243 = n2240 | n2242 ;
  assign n2244 = n584 & n2005 ;
  assign n2245 = n2243 | n2244 ;
  assign n2246 = n2243 & n2244 ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = n646 & ~n2051 ;
  assign n2249 = ( n2005 & ~n2055 ) | ( n2005 & n2248 ) | ( ~n2055 & n2248 ) ;
  assign n2250 = ( n2233 & n2247 ) | ( n2233 & n2249 ) | ( n2247 & n2249 ) ;
  assign n2251 = ( ~n2233 & n2247 ) | ( ~n2233 & n2249 ) | ( n2247 & n2249 ) ;
  assign n2252 = ( n2233 & ~n2250 ) | ( n2233 & n2251 ) | ( ~n2250 & n2251 ) ;
  assign n2253 = n1899 & n1991 ;
  assign n2254 = n1897 & n1994 ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = ~n1914 & n1997 ;
  assign n2257 = n2255 | n2256 ;
  assign n2258 = ( n1985 & ~n2136 ) | ( n1985 & n2257 ) | ( ~n2136 & n2257 ) ;
  assign n2259 = n902 | n2257 ;
  assign n2260 = ~n2258 & n2259 ;
  assign n2261 = ( ~n2257 & n2258 ) | ( ~n2257 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2262 = ( ~n902 & n2260 ) | ( ~n902 & n2261 ) | ( n2260 & n2261 ) ;
  assign n2263 = ( n2117 & n2252 ) | ( n2117 & n2262 ) | ( n2252 & n2262 ) ;
  assign n2264 = ( n2117 & ~n2252 ) | ( n2117 & n2262 ) | ( ~n2252 & n2262 ) ;
  assign n2265 = ( n2252 & ~n2263 ) | ( n2252 & n2264 ) | ( ~n2263 & n2264 ) ;
  assign n2266 = ( n1968 & n2223 ) | ( n1968 & n2265 ) | ( n2223 & n2265 ) ;
  assign n2267 = n1897 & n1991 ;
  assign n2268 = ~n1914 & n1994 ;
  assign n2269 = n2267 | n2268 ;
  assign n2270 = n1895 & n1997 ;
  assign n2271 = n2269 | n2270 ;
  assign n2272 = ( n1985 & ~n2122 ) | ( n1985 & n2271 ) | ( ~n2122 & n2271 ) ;
  assign n2273 = n902 | n2271 ;
  assign n2274 = ~n2272 & n2273 ;
  assign n2275 = ( ~n2271 & n2272 ) | ( ~n2271 & n2273 ) | ( n2272 & n2273 ) ;
  assign n2276 = ( ~n902 & n2274 ) | ( ~n902 & n2275 ) | ( n2274 & n2275 ) ;
  assign n2277 = ~n2036 & n2238 ;
  assign n2278 = n1903 & n2236 ;
  assign n2279 = ~n1901 & n2241 ;
  assign n2280 = n2278 | n2279 ;
  assign n2281 = ~n584 & n1076 ;
  assign n2282 = ( n1606 & ~n2234 ) | ( n1606 & n2281 ) | ( ~n2234 & n2281 ) ;
  assign n2283 = n1925 & n2282 ;
  assign n2284 = n2280 | n2283 ;
  assign n2285 = n2277 | n2284 ;
  assign n2286 = ~n584 & n2285 ;
  assign n2287 = n2005 | n2243 ;
  assign n2288 = ( n584 & n2285 ) | ( n584 & n2287 ) | ( n2285 & n2287 ) ;
  assign n2289 = n2285 & n2287 ;
  assign n2290 = ( n2286 & n2288 ) | ( n2286 & ~n2289 ) | ( n2288 & ~n2289 ) ;
  assign n2291 = n1906 & n2023 ;
  assign n2292 = n1909 & n2026 ;
  assign n2293 = n2291 | n2292 ;
  assign n2294 = n1899 & n2012 ;
  assign n2295 = n2293 | n2294 ;
  assign n2296 = ( n2011 & n2058 ) | ( n2011 & n2295 ) | ( n2058 & n2295 ) ;
  assign n2297 = n646 & ~n2295 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = ( n2295 & ~n2296 ) | ( n2295 & n2297 ) | ( ~n2296 & n2297 ) ;
  assign n2300 = ( ~n646 & n2298 ) | ( ~n646 & n2299 ) | ( n2298 & n2299 ) ;
  assign n2301 = ( n2250 & ~n2290 ) | ( n2250 & n2300 ) | ( ~n2290 & n2300 ) ;
  assign n2302 = ( n2250 & n2290 ) | ( n2250 & n2300 ) | ( n2290 & n2300 ) ;
  assign n2303 = ( n2290 & n2301 ) | ( n2290 & ~n2302 ) | ( n2301 & ~n2302 ) ;
  assign n2304 = ( n2263 & n2276 ) | ( n2263 & n2303 ) | ( n2276 & n2303 ) ;
  assign n2305 = ( ~n2263 & n2276 ) | ( ~n2263 & n2303 ) | ( n2276 & n2303 ) ;
  assign n2306 = ( n2263 & ~n2304 ) | ( n2263 & n2305 ) | ( ~n2304 & n2305 ) ;
  assign n2307 = ( n1954 & n2266 ) | ( n1954 & n2306 ) | ( n2266 & n2306 ) ;
  assign n2308 = ( ~n1954 & n2266 ) | ( ~n1954 & n2306 ) | ( n2266 & n2306 ) ;
  assign n2309 = ( n1954 & ~n2307 ) | ( n1954 & n2308 ) | ( ~n2307 & n2308 ) ;
  assign n2310 = ( x0 & x1 ) | ( x0 & ~x2 ) | ( x1 & ~x2 ) ;
  assign n2311 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n2312 = n2310 & n2311 ;
  assign n2313 = x0 & ~n2312 ;
  assign n2314 = n511 | n853 ;
  assign n2315 = n958 | n2314 ;
  assign n2316 = n427 | n2315 ;
  assign n2317 = n1820 | n2316 ;
  assign n2318 = n1189 | n2317 ;
  assign n2319 = n173 | n214 ;
  assign n2320 = n127 | n2319 ;
  assign n2321 = n356 | n2320 ;
  assign n2322 = n736 | n2321 ;
  assign n2323 = n1586 | n1693 ;
  assign n2324 = n2322 | n2323 ;
  assign n2325 = n2318 | n2324 ;
  assign n2326 = n1891 & ~n2325 ;
  assign n2327 = n127 | n321 ;
  assign n2328 = n1724 | n2327 ;
  assign n2329 = n180 | n257 ;
  assign n2330 = n240 | n2329 ;
  assign n2331 = n2328 | n2330 ;
  assign n2332 = n400 | n1692 ;
  assign n2333 = n2331 | n2332 ;
  assign n2334 = n678 | n1172 ;
  assign n2335 = n2333 | n2334 ;
  assign n2336 = n722 | n2335 ;
  assign n2337 = n203 | n1632 ;
  assign n2338 = n196 | n360 ;
  assign n2339 = n745 | n2338 ;
  assign n2340 = n69 | n463 ;
  assign n2341 = n170 | n2340 ;
  assign n2342 = n2339 | n2341 ;
  assign n2343 = n2337 | n2342 ;
  assign n2344 = n297 | n362 ;
  assign n2345 = n279 | n2344 ;
  assign n2346 = n1795 | n2345 ;
  assign n2347 = n372 | n1757 ;
  assign n2348 = n1752 | n2347 ;
  assign n2349 = n567 | n2348 ;
  assign n2350 = n2346 | n2349 ;
  assign n2351 = n2343 | n2350 ;
  assign n2352 = n2336 | n2351 ;
  assign n2353 = n2326 & ~n2352 ;
  assign n2354 = n538 | n671 ;
  assign n2355 = n1655 | n2354 ;
  assign n2356 = n515 & ~n880 ;
  assign n2357 = ~n1642 & n2356 ;
  assign n2358 = ~n2355 & n2357 ;
  assign n2359 = n1689 | n1771 ;
  assign n2360 = n2358 & ~n2359 ;
  assign n2361 = ~n639 & n2360 ;
  assign n2362 = ~n556 & n2361 ;
  assign n2363 = n2353 & n2362 ;
  assign n2364 = n2353 | n2362 ;
  assign n2365 = ~n2363 & n2364 ;
  assign n2366 = ~n2326 & n2352 ;
  assign n2367 = n2353 | n2366 ;
  assign n2368 = ~n1891 & n2325 ;
  assign n2369 = n2326 | n2368 ;
  assign n2370 = n1893 & ~n1922 ;
  assign n2371 = n2369 & ~n2370 ;
  assign n2372 = n2367 | n2371 ;
  assign n2373 = ~n2365 & n2372 ;
  assign n2374 = ~n1893 & n1935 ;
  assign n2375 = n2369 | n2374 ;
  assign n2376 = n2367 & n2375 ;
  assign n2377 = ~n2365 & n2376 ;
  assign n2378 = ( n2365 & ~n2372 ) | ( n2365 & n2376 ) | ( ~n2372 & n2376 ) ;
  assign n2379 = ( n2373 & ~n2377 ) | ( n2373 & n2378 ) | ( ~n2377 & n2378 ) ;
  assign n2380 = n2312 & ~n2365 ;
  assign n2381 = ~x0 & x1 ;
  assign n2382 = n2367 & n2381 ;
  assign n2383 = n2380 | n2382 ;
  assign n2384 = ( n2313 & ~n2379 ) | ( n2313 & n2383 ) | ( ~n2379 & n2383 ) ;
  assign n2385 = n231 & ~n2383 ;
  assign n2386 = n2384 | n2385 ;
  assign n2387 = ( n2383 & ~n2384 ) | ( n2383 & n2385 ) | ( ~n2384 & n2385 ) ;
  assign n2388 = ( ~n231 & n2386 ) | ( ~n231 & n2387 ) | ( n2386 & n2387 ) ;
  assign n2389 = x2 & ~n25 ;
  assign n2390 = n2369 & n2389 ;
  assign n2391 = n2388 & ~n2390 ;
  assign n2392 = n2367 & n2371 ;
  assign n2393 = ( n2367 & ~n2371 ) | ( n2367 & n2375 ) | ( ~n2371 & n2375 ) ;
  assign n2394 = ( ~n2376 & n2392 ) | ( ~n2376 & n2393 ) | ( n2392 & n2393 ) ;
  assign n2395 = n2369 & n2381 ;
  assign n2396 = n2312 & n2367 ;
  assign n2397 = n2395 | n2396 ;
  assign n2398 = ( n2313 & n2394 ) | ( n2313 & n2397 ) | ( n2394 & n2397 ) ;
  assign n2399 = n231 & ~n2397 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = ( n2397 & ~n2398 ) | ( n2397 & n2399 ) | ( ~n2398 & n2399 ) ;
  assign n2402 = ( ~n231 & n2400 ) | ( ~n231 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2403 = ~n1893 & n2389 ;
  assign n2404 = n2402 & ~n2403 ;
  assign n2405 = ( ~n1968 & n2223 ) | ( ~n1968 & n2265 ) | ( n2223 & n2265 ) ;
  assign n2406 = ( n1968 & ~n2266 ) | ( n1968 & n2405 ) | ( ~n2266 & n2405 ) ;
  assign n2407 = n2369 & n2370 ;
  assign n2408 = ( ~n2369 & n2370 ) | ( ~n2369 & n2374 ) | ( n2370 & n2374 ) ;
  assign n2409 = n2369 & ~n2374 ;
  assign n2410 = ( ~n2407 & n2408 ) | ( ~n2407 & n2409 ) | ( n2408 & n2409 ) ;
  assign n2411 = ~n1893 & n2381 ;
  assign n2412 = n2312 & n2369 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = ( n2313 & ~n2410 ) | ( n2313 & n2413 ) | ( ~n2410 & n2413 ) ;
  assign n2415 = n231 & ~n2413 ;
  assign n2416 = n2414 | n2415 ;
  assign n2417 = ( n2413 & ~n2414 ) | ( n2413 & n2415 ) | ( ~n2414 & n2415 ) ;
  assign n2418 = ( ~n231 & n2416 ) | ( ~n231 & n2417 ) | ( n2416 & n2417 ) ;
  assign n2419 = n1921 & n2389 ;
  assign n2420 = n2418 & ~n2419 ;
  assign n2421 = n1958 & n2313 ;
  assign n2422 = n231 & n2421 ;
  assign n2423 = n1918 & n2381 ;
  assign n2424 = n1921 & n2312 ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = ( ~n231 & n2421 ) | ( ~n231 & n2425 ) | ( n2421 & n2425 ) ;
  assign n2427 = n231 & ~n2389 ;
  assign n2428 = ( n231 & ~n1895 ) | ( n231 & n2427 ) | ( ~n1895 & n2427 ) ;
  assign n2429 = ~n2425 & n2428 ;
  assign n2430 = ( ~n2422 & n2426 ) | ( ~n2422 & n2429 ) | ( n2426 & n2429 ) ;
  assign n2431 = ( ~n2146 & n2216 ) | ( ~n2146 & n2218 ) | ( n2216 & n2218 ) ;
  assign n2432 = ( n2146 & ~n2219 ) | ( n2146 & n2431 ) | ( ~n2219 & n2431 ) ;
  assign n2433 = n1971 & n2313 ;
  assign n2434 = n231 & n2433 ;
  assign n2435 = n1895 & n2381 ;
  assign n2436 = n1918 & n2312 ;
  assign n2437 = n2435 | n2436 ;
  assign n2438 = ( ~n231 & n2433 ) | ( ~n231 & n2437 ) | ( n2433 & n2437 ) ;
  assign n2439 = ( n231 & n1914 ) | ( n231 & n2427 ) | ( n1914 & n2427 ) ;
  assign n2440 = ~n2437 & n2439 ;
  assign n2441 = ( ~n2434 & n2438 ) | ( ~n2434 & n2440 ) | ( n2438 & n2440 ) ;
  assign n2442 = ~n2122 & n2313 ;
  assign n2443 = n231 & n2442 ;
  assign n2444 = ~n1914 & n2381 ;
  assign n2445 = n1895 & n2312 ;
  assign n2446 = n2444 | n2445 ;
  assign n2447 = ( ~n231 & n2442 ) | ( ~n231 & n2446 ) | ( n2442 & n2446 ) ;
  assign n2448 = ( n231 & ~n1897 ) | ( n231 & n2427 ) | ( ~n1897 & n2427 ) ;
  assign n2449 = ~n2446 & n2448 ;
  assign n2450 = ( ~n2443 & n2447 ) | ( ~n2443 & n2449 ) | ( n2447 & n2449 ) ;
  assign n2451 = ( ~n2166 & n2170 ) | ( ~n2166 & n2214 ) | ( n2170 & n2214 ) ;
  assign n2452 = ( n2166 & ~n2215 ) | ( n2166 & n2451 ) | ( ~n2215 & n2451 ) ;
  assign n2453 = n1988 & n2313 ;
  assign n2454 = n231 & n2453 ;
  assign n2455 = n1899 & n2381 ;
  assign n2456 = n1897 & n2312 ;
  assign n2457 = n2455 | n2456 ;
  assign n2458 = ( ~n231 & n2453 ) | ( ~n231 & n2457 ) | ( n2453 & n2457 ) ;
  assign n2459 = ( n231 & ~n1909 ) | ( n231 & n2427 ) | ( ~n1909 & n2427 ) ;
  assign n2460 = ~n2457 & n2459 ;
  assign n2461 = ( ~n2454 & n2458 ) | ( ~n2454 & n2460 ) | ( n2458 & n2460 ) ;
  assign n2462 = n2058 & n2313 ;
  assign n2463 = n231 & n2462 ;
  assign n2464 = n1909 & n2381 ;
  assign n2465 = n1899 & n2312 ;
  assign n2466 = n2464 | n2465 ;
  assign n2467 = ( ~n231 & n2462 ) | ( ~n231 & n2466 ) | ( n2462 & n2466 ) ;
  assign n2468 = ( n231 & ~n1906 ) | ( n231 & n2427 ) | ( ~n1906 & n2427 ) ;
  assign n2469 = ~n2466 & n2468 ;
  assign n2470 = ( ~n2463 & n2467 ) | ( ~n2463 & n2469 ) | ( n2467 & n2469 ) ;
  assign n2471 = ~n222 & n2206 ;
  assign n2472 = n2199 & n2206 ;
  assign n2473 = ( n2207 & n2471 ) | ( n2207 & ~n2472 ) | ( n2471 & ~n2472 ) ;
  assign n2474 = n1903 & n2389 ;
  assign n2475 = ~n1901 & n2381 ;
  assign n2476 = n2474 | n2475 ;
  assign n2477 = n1906 & n2312 ;
  assign n2478 = n2476 | n2477 ;
  assign n2479 = ~n2017 & n2313 ;
  assign n2480 = n2478 | n2479 ;
  assign n2481 = n2193 & n2198 ;
  assign n2482 = n2199 & ~n2481 ;
  assign n2483 = ( n231 & n2480 ) | ( n231 & n2482 ) | ( n2480 & n2482 ) ;
  assign n2484 = n231 & ~n2041 ;
  assign n2485 = n1901 | n2192 ;
  assign n2486 = ( n2192 & n2484 ) | ( n2192 & n2485 ) | ( n2484 & n2485 ) ;
  assign n2487 = ( n231 & n2480 ) | ( n231 & ~n2486 ) | ( n2480 & ~n2486 ) ;
  assign n2488 = n2483 & ~n2487 ;
  assign n2489 = n2480 & n2486 ;
  assign n2490 = ~n231 & n2482 ;
  assign n2491 = ( ~n231 & n2489 ) | ( ~n231 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = n1906 & n2381 ;
  assign n2493 = n1909 & n2312 ;
  assign n2494 = n2492 | n2493 ;
  assign n2495 = n2073 & n2313 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = ~n2491 & n2496 ;
  assign n2498 = ~n2480 & n2486 ;
  assign n2499 = ( n231 & n1901 ) | ( n231 & n2427 ) | ( n1901 & n2427 ) ;
  assign n2500 = n2482 & n2499 ;
  assign n2501 = ( n2498 & n2499 ) | ( n2498 & n2500 ) | ( n2499 & n2500 ) ;
  assign n2502 = n2496 | n2501 ;
  assign n2503 = ( n2488 & ~n2497 ) | ( n2488 & n2502 ) | ( ~n2497 & n2502 ) ;
  assign n2504 = ( n2470 & n2473 ) | ( n2470 & n2503 ) | ( n2473 & n2503 ) ;
  assign n2505 = ( n2211 & n2461 ) | ( n2211 & n2504 ) | ( n2461 & n2504 ) ;
  assign n2506 = ~n2136 & n2313 ;
  assign n2507 = n1897 & n2381 ;
  assign n2508 = ~n1914 & n2312 ;
  assign n2509 = n2507 | n2508 ;
  assign n2510 = n1899 & ~n2389 ;
  assign n2511 = ( n1899 & n2509 ) | ( n1899 & ~n2510 ) | ( n2509 & ~n2510 ) ;
  assign n2512 = n2506 | n2511 ;
  assign n2513 = n231 & ~n2512 ;
  assign n2514 = ~n231 & n2512 ;
  assign n2515 = n2513 | n2514 ;
  assign n2516 = ( ~n2180 & n2184 ) | ( ~n2180 & n2213 ) | ( n2184 & n2213 ) ;
  assign n2517 = ( n2180 & ~n2214 ) | ( n2180 & n2516 ) | ( ~n2214 & n2516 ) ;
  assign n2518 = ( n2505 & n2515 ) | ( n2505 & n2517 ) | ( n2515 & n2517 ) ;
  assign n2519 = ( n2450 & n2452 ) | ( n2450 & n2518 ) | ( n2452 & n2518 ) ;
  assign n2520 = ( ~n2112 & n2156 ) | ( ~n2112 & n2215 ) | ( n2156 & n2215 ) ;
  assign n2521 = ( n2112 & ~n2216 ) | ( n2112 & n2520 ) | ( ~n2216 & n2520 ) ;
  assign n2522 = ( n2441 & n2519 ) | ( n2441 & n2521 ) | ( n2519 & n2521 ) ;
  assign n2523 = ( n2430 & n2432 ) | ( n2430 & n2522 ) | ( n2432 & n2522 ) ;
  assign n2524 = ( ~n2132 & n2219 ) | ( ~n2132 & n2221 ) | ( n2219 & n2221 ) ;
  assign n2525 = ( n2132 & ~n2222 ) | ( n2132 & n2524 ) | ( ~n2222 & n2524 ) ;
  assign n2526 = n1921 & n2381 ;
  assign n2527 = ~n1893 & n2312 ;
  assign n2528 = n2526 | n2527 ;
  assign n2529 = ( ~n1938 & n2313 ) | ( ~n1938 & n2528 ) | ( n2313 & n2528 ) ;
  assign n2530 = n231 | n2528 ;
  assign n2531 = ~n2529 & n2530 ;
  assign n2532 = ( ~n2528 & n2529 ) | ( ~n2528 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2533 = ( ~n231 & n2531 ) | ( ~n231 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2534 = n1918 & n2389 ;
  assign n2535 = n2533 & ~n2534 ;
  assign n2536 = ( n2523 & n2525 ) | ( n2523 & n2535 ) | ( n2525 & n2535 ) ;
  assign n2537 = ( ~n1981 & n2119 ) | ( ~n1981 & n2222 ) | ( n2119 & n2222 ) ;
  assign n2538 = ( n1981 & ~n2223 ) | ( n1981 & n2537 ) | ( ~n2223 & n2537 ) ;
  assign n2539 = ( n2420 & n2536 ) | ( n2420 & n2538 ) | ( n2536 & n2538 ) ;
  assign n2540 = ( n2404 & n2406 ) | ( n2404 & n2539 ) | ( n2406 & n2539 ) ;
  assign n2541 = ( n2309 & n2391 ) | ( n2309 & n2540 ) | ( n2391 & n2540 ) ;
  assign n2542 = ( ~n2309 & n2391 ) | ( ~n2309 & n2540 ) | ( n2391 & n2540 ) ;
  assign n2543 = ( n2309 & ~n2541 ) | ( n2309 & n2542 ) | ( ~n2541 & n2542 ) ;
  assign n2544 = n219 & n2543 ;
  assign n2545 = n863 | n984 ;
  assign n2546 = n530 | n674 ;
  assign n2547 = n597 | n2546 ;
  assign n2548 = n2545 | n2547 ;
  assign n2549 = n315 | n521 ;
  assign n2550 = n1583 | n2549 ;
  assign n2551 = n2548 | n2550 ;
  assign n2552 = n996 | n2551 ;
  assign n2553 = n150 | n259 ;
  assign n2554 = n754 | n2553 ;
  assign n2555 = n2552 | n2554 ;
  assign n2556 = n1715 | n2329 ;
  assign n2557 = n141 | n372 ;
  assign n2558 = n254 | n2557 ;
  assign n2559 = n2556 | n2558 ;
  assign n2560 = n239 | n1757 ;
  assign n2561 = n368 | n2560 ;
  assign n2562 = n2559 | n2561 ;
  assign n2563 = n944 | n1646 ;
  assign n2564 = n188 | n203 ;
  assign n2565 = n888 | n2564 ;
  assign n2566 = n2563 | n2565 ;
  assign n2567 = n286 | n450 ;
  assign n2568 = n744 | n2567 ;
  assign n2569 = n2566 | n2568 ;
  assign n2570 = n1829 | n2569 ;
  assign n2571 = n2562 | n2570 ;
  assign n2572 = n2555 | n2571 ;
  assign n2573 = n1921 & n1941 ;
  assign n2574 = ~n1893 & n1944 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = n1947 & n2369 ;
  assign n2577 = n2575 | n2576 ;
  assign n2578 = ( n238 & ~n2410 ) | ( n238 & n2577 ) | ( ~n2410 & n2577 ) ;
  assign n2579 = n222 & ~n2577 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = ( n2577 & ~n2578 ) | ( n2577 & n2579 ) | ( ~n2578 & n2579 ) ;
  assign n2582 = ( ~n222 & n2580 ) | ( ~n222 & n2581 ) | ( n2580 & n2581 ) ;
  assign n2583 = ~n1914 & n1991 ;
  assign n2584 = n1895 & n1994 ;
  assign n2585 = n2583 | n2584 ;
  assign n2586 = n1918 & n1997 ;
  assign n2587 = n2585 | n2586 ;
  assign n2588 = ( n1971 & n1985 ) | ( n1971 & n2587 ) | ( n1985 & n2587 ) ;
  assign n2589 = n902 & ~n2587 ;
  assign n2590 = n2588 | n2589 ;
  assign n2591 = ( n2587 & ~n2588 ) | ( n2587 & n2589 ) | ( ~n2588 & n2589 ) ;
  assign n2592 = ( ~n902 & n2590 ) | ( ~n902 & n2591 ) | ( n2590 & n2591 ) ;
  assign n2593 = n2285 | n2287 ;
  assign n2594 = ( n584 & n1925 ) | ( n584 & n2593 ) | ( n1925 & n2593 ) ;
  assign n2595 = n1903 & n2282 ;
  assign n2596 = ~n1901 & n2236 ;
  assign n2597 = n2595 | n2596 ;
  assign n2598 = n1906 & n2241 ;
  assign n2599 = n2597 | n2598 ;
  assign n2600 = ~n2017 & n2238 ;
  assign n2601 = n2599 | n2600 ;
  assign n2602 = n1925 & n2593 ;
  assign n2603 = ( ~n2594 & n2601 ) | ( ~n2594 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = ( n2594 & n2601 ) | ( n2594 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2605 = ( n2594 & n2603 ) | ( n2594 & ~n2604 ) | ( n2603 & ~n2604 ) ;
  assign n2606 = n1909 & n2023 ;
  assign n2607 = n1899 & n2026 ;
  assign n2608 = n2606 | n2607 ;
  assign n2609 = n1897 & n2012 ;
  assign n2610 = n2608 | n2609 ;
  assign n2611 = ( n1988 & n2011 ) | ( n1988 & n2610 ) | ( n2011 & n2610 ) ;
  assign n2612 = n646 | n2610 ;
  assign n2613 = ~n2611 & n2612 ;
  assign n2614 = ( ~n2610 & n2611 ) | ( ~n2610 & n2612 ) | ( n2611 & n2612 ) ;
  assign n2615 = ( ~n646 & n2613 ) | ( ~n646 & n2614 ) | ( n2613 & n2614 ) ;
  assign n2616 = ( n2302 & ~n2605 ) | ( n2302 & n2615 ) | ( ~n2605 & n2615 ) ;
  assign n2617 = ( n2302 & n2605 ) | ( n2302 & n2615 ) | ( n2605 & n2615 ) ;
  assign n2618 = ( n2605 & n2616 ) | ( n2605 & ~n2617 ) | ( n2616 & ~n2617 ) ;
  assign n2619 = ( n2304 & n2592 ) | ( n2304 & n2618 ) | ( n2592 & n2618 ) ;
  assign n2620 = ( ~n2304 & n2592 ) | ( ~n2304 & n2618 ) | ( n2592 & n2618 ) ;
  assign n2621 = ( n2304 & ~n2619 ) | ( n2304 & n2620 ) | ( ~n2619 & n2620 ) ;
  assign n2622 = ( n2307 & n2582 ) | ( n2307 & n2621 ) | ( n2582 & n2621 ) ;
  assign n2623 = ( n2307 & ~n2582 ) | ( n2307 & n2621 ) | ( ~n2582 & n2621 ) ;
  assign n2624 = ( n2582 & ~n2622 ) | ( n2582 & n2623 ) | ( ~n2622 & n2623 ) ;
  assign n2625 = n207 | n251 ;
  assign n2626 = n976 | n2625 ;
  assign n2627 = n1589 | n2626 ;
  assign n2628 = n576 | n1005 ;
  assign n2629 = n613 | n2628 ;
  assign n2630 = n2627 | n2629 ;
  assign n2631 = n475 | n622 ;
  assign n2632 = n2630 | n2631 ;
  assign n2633 = n2363 & ~n2632 ;
  assign n2634 = ( n556 & ~n2363 ) | ( n556 & n2632 ) | ( ~n2363 & n2632 ) ;
  assign n2635 = n2633 | n2634 ;
  assign n2636 = n2373 & ~n2635 ;
  assign n2637 = n2365 & ~n2376 ;
  assign n2638 = ( n2373 & n2635 ) | ( n2373 & n2637 ) | ( n2635 & n2637 ) ;
  assign n2639 = n2635 | n2637 ;
  assign n2640 = ( n2636 & ~n2638 ) | ( n2636 & n2639 ) | ( ~n2638 & n2639 ) ;
  assign n2641 = n2312 & n2635 ;
  assign n2642 = ~n2365 & n2381 ;
  assign n2643 = n2641 | n2642 ;
  assign n2644 = ( n2313 & ~n2640 ) | ( n2313 & n2643 ) | ( ~n2640 & n2643 ) ;
  assign n2645 = n231 | n2643 ;
  assign n2646 = ~n2644 & n2645 ;
  assign n2647 = ( ~n2643 & n2644 ) | ( ~n2643 & n2645 ) | ( n2644 & n2645 ) ;
  assign n2648 = ( ~n231 & n2646 ) | ( ~n231 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2649 = n2367 & n2389 ;
  assign n2650 = n2648 & ~n2649 ;
  assign n2651 = ( n2541 & n2624 ) | ( n2541 & n2650 ) | ( n2624 & n2650 ) ;
  assign n2652 = ( n2541 & ~n2624 ) | ( n2541 & n2650 ) | ( ~n2624 & n2650 ) ;
  assign n2653 = ( n2624 & ~n2651 ) | ( n2624 & n2652 ) | ( ~n2651 & n2652 ) ;
  assign n2654 = ( n2544 & n2572 ) | ( n2544 & n2653 ) | ( n2572 & n2653 ) ;
  assign n2655 = n106 & n204 ;
  assign n2656 = n636 | n2655 ;
  assign n2657 = n146 | n616 ;
  assign n2658 = n2656 | n2657 ;
  assign n2659 = n601 | n2658 ;
  assign n2660 = n556 | n2659 ;
  assign n2661 = ~n2633 & n2660 ;
  assign n2662 = n2373 | n2635 ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = n2635 & ~n2637 ;
  assign n2665 = ( n2661 & ~n2662 ) | ( n2661 & n2664 ) | ( ~n2662 & n2664 ) ;
  assign n2666 = n2661 | n2664 ;
  assign n2667 = ( n2663 & n2665 ) | ( n2663 & ~n2666 ) | ( n2665 & ~n2666 ) ;
  assign n2668 = n2312 & n2661 ;
  assign n2669 = n2381 & n2635 ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = ( n2313 & n2667 ) | ( n2313 & n2670 ) | ( n2667 & n2670 ) ;
  assign n2672 = n231 | n2670 ;
  assign n2673 = ~n2671 & n2672 ;
  assign n2674 = ( ~n2670 & n2671 ) | ( ~n2670 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2675 = ( ~n231 & n2673 ) | ( ~n231 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = ~n2365 & n2389 ;
  assign n2677 = n2675 & ~n2676 ;
  assign n2678 = n1944 & n2369 ;
  assign n2679 = n238 | n2678 ;
  assign n2680 = ( n2394 & n2678 ) | ( n2394 & n2679 ) | ( n2678 & n2679 ) ;
  assign n2681 = ~n1893 & n1941 ;
  assign n2682 = n1947 & n2367 ;
  assign n2683 = n2681 | n2682 ;
  assign n2684 = ( n222 & n2680 ) | ( n222 & n2683 ) | ( n2680 & n2683 ) ;
  assign n2685 = n222 | n2680 ;
  assign n2686 = ( ~n222 & n2680 ) | ( ~n222 & n2683 ) | ( n2680 & n2683 ) ;
  assign n2687 = ( ~n2684 & n2685 ) | ( ~n2684 & n2686 ) | ( n2685 & n2686 ) ;
  assign n2688 = n1895 & n1991 ;
  assign n2689 = n1918 & n1994 ;
  assign n2690 = n2688 | n2689 ;
  assign n2691 = n1921 & n1997 ;
  assign n2692 = n2690 | n2691 ;
  assign n2693 = ( n1958 & n1985 ) | ( n1958 & n2692 ) | ( n1985 & n2692 ) ;
  assign n2694 = n902 & ~n2692 ;
  assign n2695 = n2693 | n2694 ;
  assign n2696 = ( n2692 & ~n2693 ) | ( n2692 & n2694 ) | ( ~n2693 & n2694 ) ;
  assign n2697 = ( ~n902 & n2695 ) | ( ~n902 & n2696 ) | ( n2695 & n2696 ) ;
  assign n2698 = ~n1925 & n2593 ;
  assign n2699 = n2601 | n2698 ;
  assign n2700 = ( n584 & n1903 ) | ( n584 & n2699 ) | ( n1903 & n2699 ) ;
  assign n2701 = ~n1901 & n2282 ;
  assign n2702 = n1906 & n2236 ;
  assign n2703 = n2701 | n2702 ;
  assign n2704 = n1909 & n2241 ;
  assign n2705 = n2703 | n2704 ;
  assign n2706 = n2073 & n2238 ;
  assign n2707 = n2705 | n2706 ;
  assign n2708 = n1903 & n2699 ;
  assign n2709 = ( ~n2700 & n2707 ) | ( ~n2700 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2710 = ( n2700 & n2707 ) | ( n2700 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2711 = ( n2700 & n2709 ) | ( n2700 & ~n2710 ) | ( n2709 & ~n2710 ) ;
  assign n2712 = n1899 & n2023 ;
  assign n2713 = n1897 & n2026 ;
  assign n2714 = n2712 | n2713 ;
  assign n2715 = ~n1914 & n2012 ;
  assign n2716 = n2714 | n2715 ;
  assign n2717 = ( n2011 & ~n2136 ) | ( n2011 & n2716 ) | ( ~n2136 & n2716 ) ;
  assign n2718 = n646 | n2716 ;
  assign n2719 = ~n2717 & n2718 ;
  assign n2720 = ( ~n2716 & n2717 ) | ( ~n2716 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2721 = ( ~n646 & n2719 ) | ( ~n646 & n2720 ) | ( n2719 & n2720 ) ;
  assign n2722 = ( n2617 & ~n2711 ) | ( n2617 & n2721 ) | ( ~n2711 & n2721 ) ;
  assign n2723 = ( n2617 & n2711 ) | ( n2617 & n2721 ) | ( n2711 & n2721 ) ;
  assign n2724 = ( n2711 & n2722 ) | ( n2711 & ~n2723 ) | ( n2722 & ~n2723 ) ;
  assign n2725 = ( n2619 & n2697 ) | ( n2619 & n2724 ) | ( n2697 & n2724 ) ;
  assign n2726 = ( ~n2619 & n2697 ) | ( ~n2619 & n2724 ) | ( n2697 & n2724 ) ;
  assign n2727 = ( n2619 & ~n2725 ) | ( n2619 & n2726 ) | ( ~n2725 & n2726 ) ;
  assign n2728 = ( ~n2622 & n2687 ) | ( ~n2622 & n2727 ) | ( n2687 & n2727 ) ;
  assign n2729 = ( n2622 & n2687 ) | ( n2622 & n2727 ) | ( n2687 & n2727 ) ;
  assign n2730 = ( n2622 & n2728 ) | ( n2622 & ~n2729 ) | ( n2728 & ~n2729 ) ;
  assign n2731 = ( n2651 & n2677 ) | ( n2651 & n2730 ) | ( n2677 & n2730 ) ;
  assign n2732 = ( n2651 & ~n2677 ) | ( n2651 & n2730 ) | ( ~n2677 & n2730 ) ;
  assign n2733 = ( n2677 & ~n2731 ) | ( n2677 & n2732 ) | ( ~n2731 & n2732 ) ;
  assign n2734 = n1000 | n1674 ;
  assign n2735 = n277 | n521 ;
  assign n2736 = n311 | n2735 ;
  assign n2737 = n2734 | n2736 ;
  assign n2738 = n146 | n261 ;
  assign n2739 = n127 | n728 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n1166 | n2740 ;
  assign n2742 = n316 | n547 ;
  assign n2743 = n2741 | n2742 ;
  assign n2744 = n2737 | n2743 ;
  assign n2745 = n195 | n378 ;
  assign n2746 = n492 | n2745 ;
  assign n2747 = n2744 | n2746 ;
  assign n2748 = n1170 | n1594 ;
  assign n2749 = n300 | n328 ;
  assign n2750 = n428 | n485 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n1806 | n2347 ;
  assign n2753 = n2751 | n2752 ;
  assign n2754 = n2748 | n2753 ;
  assign n2755 = n278 | n443 ;
  assign n2756 = n496 | n2755 ;
  assign n2757 = n2346 | n2756 ;
  assign n2758 = n327 | n2757 ;
  assign n2759 = n256 | n2758 ;
  assign n2760 = n2754 | n2759 ;
  assign n2761 = n2747 | n2760 ;
  assign n2762 = ( ~n2654 & n2733 ) | ( ~n2654 & n2761 ) | ( n2733 & n2761 ) ;
  assign n2763 = n365 | n1175 ;
  assign n2764 = n2661 & n2662 ;
  assign n2765 = ~n553 & n2764 ;
  assign n2766 = ( n553 & ~n2666 ) | ( n553 & n2764 ) | ( ~n2666 & n2764 ) ;
  assign n2767 = ~n553 & n2666 ;
  assign n2768 = ( ~n2765 & n2766 ) | ( ~n2765 & n2767 ) | ( n2766 & n2767 ) ;
  assign n2769 = ~n553 & n2312 ;
  assign n2770 = n2381 | n2769 ;
  assign n2771 = ( n2661 & n2769 ) | ( n2661 & n2770 ) | ( n2769 & n2770 ) ;
  assign n2772 = ( n2313 & ~n2768 ) | ( n2313 & n2771 ) | ( ~n2768 & n2771 ) ;
  assign n2773 = n231 & ~n2771 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = ( n2771 & ~n2772 ) | ( n2771 & n2773 ) | ( ~n2772 & n2773 ) ;
  assign n2776 = ( ~n231 & n2774 ) | ( ~n231 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2777 = n2389 & n2635 ;
  assign n2778 = n2776 & ~n2777 ;
  assign n2779 = n238 & ~n2379 ;
  assign n2780 = n222 & n2779 ;
  assign n2781 = n1941 & n2369 ;
  assign n2782 = n1944 & n2367 ;
  assign n2783 = n2781 | n2782 ;
  assign n2784 = n1947 & ~n2365 ;
  assign n2785 = n2783 | n2784 ;
  assign n2786 = ( ~n222 & n2779 ) | ( ~n222 & n2785 ) | ( n2779 & n2785 ) ;
  assign n2787 = n222 & ~n2785 ;
  assign n2788 = ( ~n2780 & n2786 ) | ( ~n2780 & n2787 ) | ( n2786 & n2787 ) ;
  assign n2789 = n1918 & n1991 ;
  assign n2790 = n1921 & n1994 ;
  assign n2791 = n2789 | n2790 ;
  assign n2792 = ~n1893 & n1997 ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = ( ~n1938 & n1985 ) | ( ~n1938 & n2793 ) | ( n1985 & n2793 ) ;
  assign n2795 = n902 | n2793 ;
  assign n2796 = ~n2794 & n2795 ;
  assign n2797 = ( ~n2793 & n2794 ) | ( ~n2793 & n2795 ) | ( n2794 & n2795 ) ;
  assign n2798 = ( ~n902 & n2796 ) | ( ~n902 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2799 = n1897 & n2023 ;
  assign n2800 = ~n1914 & n2026 ;
  assign n2801 = n2799 | n2800 ;
  assign n2802 = n1895 & n2012 ;
  assign n2803 = n2801 | n2802 ;
  assign n2804 = ( n2011 & ~n2122 ) | ( n2011 & n2803 ) | ( ~n2122 & n2803 ) ;
  assign n2805 = n646 | n2803 ;
  assign n2806 = ~n2804 & n2805 ;
  assign n2807 = ( ~n2803 & n2804 ) | ( ~n2803 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2808 = ( ~n646 & n2806 ) | ( ~n646 & n2807 ) | ( n2806 & n2807 ) ;
  assign n2809 = ( ~n1903 & n2699 ) | ( ~n1903 & n2707 ) | ( n2699 & n2707 ) ;
  assign n2810 = ( n584 & n1901 ) | ( n584 & ~n2809 ) | ( n1901 & ~n2809 ) ;
  assign n2811 = n1906 & n2282 ;
  assign n2812 = n1909 & n2236 ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = n1899 & n2241 ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = n2058 & n2238 ;
  assign n2817 = n2815 | n2816 ;
  assign n2818 = n1901 & ~n2809 ;
  assign n2819 = ( ~n2810 & n2817 ) | ( ~n2810 & n2818 ) | ( n2817 & n2818 ) ;
  assign n2820 = ( n2810 & n2817 ) | ( n2810 & n2818 ) | ( n2817 & n2818 ) ;
  assign n2821 = ( n2810 & n2819 ) | ( n2810 & ~n2820 ) | ( n2819 & ~n2820 ) ;
  assign n2822 = ( n2723 & n2808 ) | ( n2723 & n2821 ) | ( n2808 & n2821 ) ;
  assign n2823 = ( ~n2723 & n2808 ) | ( ~n2723 & n2821 ) | ( n2808 & n2821 ) ;
  assign n2824 = ( n2723 & ~n2822 ) | ( n2723 & n2823 ) | ( ~n2822 & n2823 ) ;
  assign n2825 = ( n2725 & n2798 ) | ( n2725 & n2824 ) | ( n2798 & n2824 ) ;
  assign n2826 = ( ~n2725 & n2798 ) | ( ~n2725 & n2824 ) | ( n2798 & n2824 ) ;
  assign n2827 = ( n2725 & ~n2825 ) | ( n2725 & n2826 ) | ( ~n2825 & n2826 ) ;
  assign n2828 = ( ~n2729 & n2788 ) | ( ~n2729 & n2827 ) | ( n2788 & n2827 ) ;
  assign n2829 = ( n2729 & n2788 ) | ( n2729 & n2827 ) | ( n2788 & n2827 ) ;
  assign n2830 = ( n2729 & n2828 ) | ( n2729 & ~n2829 ) | ( n2828 & ~n2829 ) ;
  assign n2831 = ( n2731 & ~n2778 ) | ( n2731 & n2830 ) | ( ~n2778 & n2830 ) ;
  assign n2832 = ( n2731 & n2778 ) | ( n2731 & n2830 ) | ( n2778 & n2830 ) ;
  assign n2833 = ( n2778 & n2831 ) | ( n2778 & ~n2832 ) | ( n2831 & ~n2832 ) ;
  assign n2834 = ( ~n2654 & n2763 ) | ( ~n2654 & n2833 ) | ( n2763 & n2833 ) ;
  assign n2835 = ( n2654 & n2763 ) | ( n2654 & n2833 ) | ( n2763 & n2833 ) ;
  assign n2836 = ( n2654 & n2834 ) | ( n2654 & ~n2835 ) | ( n2834 & ~n2835 ) ;
  assign n2837 = n2762 & n2836 ;
  assign n2838 = n2762 | n2836 ;
  assign n2839 = ~n2837 & n2838 ;
  assign n2840 = ~x22 & x23 ;
  assign n2841 = x22 & ~x23 ;
  assign n2842 = n2840 | n2841 ;
  assign n2843 = ( n2762 & n2836 ) | ( n2762 & n2842 ) | ( n2836 & n2842 ) ;
  assign n2844 = n553 & ~n2764 ;
  assign n2845 = n300 | n319 ;
  assign n2846 = n130 | n443 ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = n177 | n1656 ;
  assign n2849 = n2847 | n2848 ;
  assign n2850 = n566 | n2849 ;
  assign n2851 = n719 | n2850 ;
  assign n2852 = n465 | n880 ;
  assign n2853 = n752 | n2852 ;
  assign n2854 = n2851 | n2853 ;
  assign n2855 = n1781 | n2854 ;
  assign n2856 = n1181 & ~n2855 ;
  assign n2857 = n664 & n2856 ;
  assign n2858 = n2844 & ~n2857 ;
  assign n2859 = ~n2844 & n2857 ;
  assign n2860 = ~n2767 & n2859 ;
  assign n2861 = n2858 | n2860 ;
  assign n2862 = n2312 & ~n2857 ;
  assign n2863 = ~n553 & n2381 ;
  assign n2864 = n2862 | n2863 ;
  assign n2865 = ( n2313 & n2861 ) | ( n2313 & n2864 ) | ( n2861 & n2864 ) ;
  assign n2866 = n231 | n2864 ;
  assign n2867 = ~n2865 & n2866 ;
  assign n2868 = ( ~n2864 & n2865 ) | ( ~n2864 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2869 = ( ~n231 & n2867 ) | ( ~n231 & n2868 ) | ( n2867 & n2868 ) ;
  assign n2870 = n2389 & n2661 ;
  assign n2871 = n2869 & ~n2870 ;
  assign n2872 = n238 & ~n2640 ;
  assign n2873 = n222 & n2872 ;
  assign n2874 = n1944 & ~n2365 ;
  assign n2875 = n1941 & n2367 ;
  assign n2876 = n2874 | n2875 ;
  assign n2877 = n1947 & n2635 ;
  assign n2878 = n2876 | n2877 ;
  assign n2879 = ( ~n222 & n2872 ) | ( ~n222 & n2878 ) | ( n2872 & n2878 ) ;
  assign n2880 = n222 & ~n2878 ;
  assign n2881 = ( ~n2873 & n2879 ) | ( ~n2873 & n2880 ) | ( n2879 & n2880 ) ;
  assign n2882 = ~n1914 & n2023 ;
  assign n2883 = n1895 & n2026 ;
  assign n2884 = n2882 | n2883 ;
  assign n2885 = n1918 & n2012 ;
  assign n2886 = n2884 | n2885 ;
  assign n2887 = ( n1971 & n2011 ) | ( n1971 & n2886 ) | ( n2011 & n2886 ) ;
  assign n2888 = n646 & ~n2886 ;
  assign n2889 = n2887 | n2888 ;
  assign n2890 = ( n2886 & ~n2887 ) | ( n2886 & n2888 ) | ( ~n2887 & n2888 ) ;
  assign n2891 = ( ~n646 & n2889 ) | ( ~n646 & n2890 ) | ( n2889 & n2890 ) ;
  assign n2892 = ( n1901 & n2809 ) | ( n1901 & n2817 ) | ( n2809 & n2817 ) ;
  assign n2893 = ( ~n584 & n1906 ) | ( ~n584 & n2892 ) | ( n1906 & n2892 ) ;
  assign n2894 = n1909 & n2282 ;
  assign n2895 = n1899 & n2236 ;
  assign n2896 = n2894 | n2895 ;
  assign n2897 = n1897 & n2241 ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = n1988 & n2238 ;
  assign n2900 = n2898 | n2899 ;
  assign n2901 = n1906 | n2892 ;
  assign n2902 = ( n2893 & n2900 ) | ( n2893 & ~n2901 ) | ( n2900 & ~n2901 ) ;
  assign n2903 = ( n2893 & ~n2900 ) | ( n2893 & n2901 ) | ( ~n2900 & n2901 ) ;
  assign n2904 = ( ~n2893 & n2902 ) | ( ~n2893 & n2903 ) | ( n2902 & n2903 ) ;
  assign n2905 = ( n2822 & n2891 ) | ( n2822 & n2904 ) | ( n2891 & n2904 ) ;
  assign n2906 = ( ~n2822 & n2891 ) | ( ~n2822 & n2904 ) | ( n2891 & n2904 ) ;
  assign n2907 = ( n2822 & ~n2905 ) | ( n2822 & n2906 ) | ( ~n2905 & n2906 ) ;
  assign n2908 = n1921 & n1991 ;
  assign n2909 = ~n1893 & n1994 ;
  assign n2910 = n2908 | n2909 ;
  assign n2911 = n1997 & n2369 ;
  assign n2912 = n2910 | n2911 ;
  assign n2913 = ( n1985 & ~n2410 ) | ( n1985 & n2912 ) | ( ~n2410 & n2912 ) ;
  assign n2914 = n902 & ~n2912 ;
  assign n2915 = n2913 | n2914 ;
  assign n2916 = ( n2912 & ~n2913 ) | ( n2912 & n2914 ) | ( ~n2913 & n2914 ) ;
  assign n2917 = ( ~n902 & n2915 ) | ( ~n902 & n2916 ) | ( n2915 & n2916 ) ;
  assign n2918 = ( n2825 & ~n2907 ) | ( n2825 & n2917 ) | ( ~n2907 & n2917 ) ;
  assign n2919 = ( n2825 & n2907 ) | ( n2825 & n2917 ) | ( n2907 & n2917 ) ;
  assign n2920 = ( n2907 & n2918 ) | ( n2907 & ~n2919 ) | ( n2918 & ~n2919 ) ;
  assign n2921 = ( n2829 & n2881 ) | ( n2829 & n2920 ) | ( n2881 & n2920 ) ;
  assign n2922 = ( ~n2829 & n2881 ) | ( ~n2829 & n2920 ) | ( n2881 & n2920 ) ;
  assign n2923 = ( n2829 & ~n2921 ) | ( n2829 & n2922 ) | ( ~n2921 & n2922 ) ;
  assign n2924 = ( n2832 & n2871 ) | ( n2832 & n2923 ) | ( n2871 & n2923 ) ;
  assign n2925 = ( ~n2832 & n2871 ) | ( ~n2832 & n2923 ) | ( n2871 & n2923 ) ;
  assign n2926 = ( n2832 & ~n2924 ) | ( n2832 & n2925 ) | ( ~n2924 & n2925 ) ;
  assign n2927 = n208 | n1858 ;
  assign n2928 = n976 | n1195 ;
  assign n2929 = n2339 | n2928 ;
  assign n2930 = n2927 | n2929 ;
  assign n2931 = n1170 | n1726 ;
  assign n2932 = n2930 | n2931 ;
  assign n2933 = n2744 | n2932 ;
  assign n2934 = n415 | n864 ;
  assign n2935 = n720 | n2934 ;
  assign n2936 = n1719 | n2935 ;
  assign n2937 = n2933 | n2936 ;
  assign n2938 = ( n2835 & n2926 ) | ( n2835 & n2937 ) | ( n2926 & n2937 ) ;
  assign n2939 = ( ~n2835 & n2926 ) | ( ~n2835 & n2937 ) | ( n2926 & n2937 ) ;
  assign n2940 = ( n2835 & ~n2938 ) | ( n2835 & n2939 ) | ( ~n2938 & n2939 ) ;
  assign n2941 = ~n2843 & n2940 ;
  assign n2942 = n2843 & ~n2940 ;
  assign n2943 = n2941 | n2942 ;
  assign n2944 = ( n2842 & n2843 ) | ( n2842 & n2940 ) | ( n2843 & n2940 ) ;
  assign n2945 = n2767 | n2858 ;
  assign n2946 = n2381 & ~n2857 ;
  assign n2947 = n2313 | n2946 ;
  assign n2948 = ( n2945 & n2946 ) | ( n2945 & n2947 ) | ( n2946 & n2947 ) ;
  assign n2949 = ~n553 & n2389 ;
  assign n2950 = ( n231 & n2948 ) | ( n231 & ~n2949 ) | ( n2948 & ~n2949 ) ;
  assign n2951 = ( n231 & n2948 ) | ( n231 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2952 = n2950 & ~n2951 ;
  assign n2953 = ~n1893 & n1991 ;
  assign n2954 = n1994 & n2369 ;
  assign n2955 = n2953 | n2954 ;
  assign n2956 = n1997 & n2367 ;
  assign n2957 = n2955 | n2956 ;
  assign n2958 = ( n1985 & n2394 ) | ( n1985 & n2957 ) | ( n2394 & n2957 ) ;
  assign n2959 = n902 & ~n2957 ;
  assign n2960 = n2958 | n2959 ;
  assign n2961 = ( n2957 & ~n2958 ) | ( n2957 & n2959 ) | ( ~n2958 & n2959 ) ;
  assign n2962 = ( ~n902 & n2960 ) | ( ~n902 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2963 = n1895 & n2023 ;
  assign n2964 = n1918 & n2026 ;
  assign n2965 = n2963 | n2964 ;
  assign n2966 = n1921 & n2012 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = ( n1958 & n2011 ) | ( n1958 & n2967 ) | ( n2011 & n2967 ) ;
  assign n2969 = n646 & ~n2967 ;
  assign n2970 = n2968 | n2969 ;
  assign n2971 = ( n2967 & ~n2968 ) | ( n2967 & n2969 ) | ( ~n2968 & n2969 ) ;
  assign n2972 = ( ~n646 & n2970 ) | ( ~n646 & n2971 ) | ( n2970 & n2971 ) ;
  assign n2973 = ( ~n1906 & n2892 ) | ( ~n1906 & n2900 ) | ( n2892 & n2900 ) ;
  assign n2974 = ( ~n584 & n1909 ) | ( ~n584 & n2973 ) | ( n1909 & n2973 ) ;
  assign n2975 = n1899 & n2282 ;
  assign n2976 = n1897 & n2236 ;
  assign n2977 = n2975 | n2976 ;
  assign n2978 = ~n1914 & n2241 ;
  assign n2979 = n2977 | n2978 ;
  assign n2980 = ~n2136 & n2238 ;
  assign n2981 = n2979 | n2980 ;
  assign n2982 = n1909 | n2973 ;
  assign n2983 = ( n2974 & n2981 ) | ( n2974 & ~n2982 ) | ( n2981 & ~n2982 ) ;
  assign n2984 = ( n2974 & ~n2981 ) | ( n2974 & n2982 ) | ( ~n2981 & n2982 ) ;
  assign n2985 = ( ~n2974 & n2983 ) | ( ~n2974 & n2984 ) | ( n2983 & n2984 ) ;
  assign n2986 = ( n2905 & n2972 ) | ( n2905 & n2985 ) | ( n2972 & n2985 ) ;
  assign n2987 = ( ~n2905 & n2972 ) | ( ~n2905 & n2985 ) | ( n2972 & n2985 ) ;
  assign n2988 = ( n2905 & ~n2986 ) | ( n2905 & n2987 ) | ( ~n2986 & n2987 ) ;
  assign n2989 = ( n2919 & n2962 ) | ( n2919 & n2988 ) | ( n2962 & n2988 ) ;
  assign n2990 = ( ~n2919 & n2962 ) | ( ~n2919 & n2988 ) | ( n2962 & n2988 ) ;
  assign n2991 = ( n2919 & ~n2989 ) | ( n2919 & n2990 ) | ( ~n2989 & n2990 ) ;
  assign n2992 = n1941 & ~n2365 ;
  assign n2993 = n1944 & n2635 ;
  assign n2994 = n2992 | n2993 ;
  assign n2995 = n1947 & n2661 ;
  assign n2996 = n2994 | n2995 ;
  assign n2997 = ( n238 & n2667 ) | ( n238 & n2996 ) | ( n2667 & n2996 ) ;
  assign n2998 = n222 | n2996 ;
  assign n2999 = ~n2997 & n2998 ;
  assign n3000 = ( ~n2996 & n2997 ) | ( ~n2996 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3001 = ( ~n222 & n2999 ) | ( ~n222 & n3000 ) | ( n2999 & n3000 ) ;
  assign n3002 = ( n2921 & ~n2991 ) | ( n2921 & n3001 ) | ( ~n2991 & n3001 ) ;
  assign n3003 = ( n2921 & n2991 ) | ( n2921 & n3001 ) | ( n2991 & n3001 ) ;
  assign n3004 = ( n2991 & n3002 ) | ( n2991 & ~n3003 ) | ( n3002 & ~n3003 ) ;
  assign n3005 = ( n2924 & n2952 ) | ( n2924 & n3004 ) | ( n2952 & n3004 ) ;
  assign n3006 = ( ~n2924 & n2952 ) | ( ~n2924 & n3004 ) | ( n2952 & n3004 ) ;
  assign n3007 = ( n2924 & ~n3005 ) | ( n2924 & n3006 ) | ( ~n3005 & n3006 ) ;
  assign n3008 = n245 | n328 ;
  assign n3009 = n1004 | n3008 ;
  assign n3010 = n261 | n1590 ;
  assign n3011 = n3009 | n3010 ;
  assign n3012 = n141 | n176 ;
  assign n3013 = n188 | n3012 ;
  assign n3014 = n199 | n390 ;
  assign n3015 = n3013 | n3014 ;
  assign n3016 = n3011 | n3015 ;
  assign n3017 = n360 | n624 ;
  assign n3018 = n369 | n3017 ;
  assign n3019 = n3016 | n3018 ;
  assign n3020 = n741 | n3019 ;
  assign n3021 = n135 | n3020 ;
  assign n3022 = ( n2938 & ~n3007 ) | ( n2938 & n3021 ) | ( ~n3007 & n3021 ) ;
  assign n3023 = ( n2938 & n3007 ) | ( n2938 & n3021 ) | ( n3007 & n3021 ) ;
  assign n3024 = ( n3007 & n3022 ) | ( n3007 & ~n3023 ) | ( n3022 & ~n3023 ) ;
  assign n3025 = n2944 | n3024 ;
  assign n3026 = n2944 & n3024 ;
  assign n3027 = n3025 & ~n3026 ;
  assign n3028 = n1918 & n2023 ;
  assign n3029 = n1921 & n2026 ;
  assign n3030 = n3028 | n3029 ;
  assign n3031 = ~n1893 & n2012 ;
  assign n3032 = n3030 | n3031 ;
  assign n3033 = ( ~n1938 & n2011 ) | ( ~n1938 & n3032 ) | ( n2011 & n3032 ) ;
  assign n3034 = n646 | n3032 ;
  assign n3035 = ~n3033 & n3034 ;
  assign n3036 = ( ~n3032 & n3033 ) | ( ~n3032 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3037 = ( ~n646 & n3035 ) | ( ~n646 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3038 = ( ~n1909 & n2973 ) | ( ~n1909 & n2981 ) | ( n2973 & n2981 ) ;
  assign n3039 = ( ~n584 & n1899 ) | ( ~n584 & n3038 ) | ( n1899 & n3038 ) ;
  assign n3040 = n1895 & n2241 ;
  assign n3041 = n1897 & n2282 ;
  assign n3042 = ~n1914 & n2236 ;
  assign n3043 = n3041 | n3042 ;
  assign n3044 = n3040 | n3043 ;
  assign n3045 = ~n2122 & n2238 ;
  assign n3046 = n3044 | n3045 ;
  assign n3047 = n1899 | n3038 ;
  assign n3048 = ( n3039 & n3046 ) | ( n3039 & ~n3047 ) | ( n3046 & ~n3047 ) ;
  assign n3049 = ( n3039 & ~n3046 ) | ( n3039 & n3047 ) | ( ~n3046 & n3047 ) ;
  assign n3050 = ( ~n3039 & n3048 ) | ( ~n3039 & n3049 ) | ( n3048 & n3049 ) ;
  assign n3051 = ( n2986 & n3037 ) | ( n2986 & n3050 ) | ( n3037 & n3050 ) ;
  assign n3052 = ( ~n2986 & n3037 ) | ( ~n2986 & n3050 ) | ( n3037 & n3050 ) ;
  assign n3053 = ( n2986 & ~n3051 ) | ( n2986 & n3052 ) | ( ~n3051 & n3052 ) ;
  assign n3054 = n1991 & n2369 ;
  assign n3055 = n1994 & n2367 ;
  assign n3056 = n3054 | n3055 ;
  assign n3057 = n1997 & ~n2365 ;
  assign n3058 = n3056 | n3057 ;
  assign n3059 = ( n1985 & ~n2379 ) | ( n1985 & n3058 ) | ( ~n2379 & n3058 ) ;
  assign n3060 = n902 & ~n3058 ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = ( n3058 & ~n3059 ) | ( n3058 & n3060 ) | ( ~n3059 & n3060 ) ;
  assign n3063 = ( ~n902 & n3061 ) | ( ~n902 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3064 = ( n2989 & ~n3053 ) | ( n2989 & n3063 ) | ( ~n3053 & n3063 ) ;
  assign n3065 = ( n2989 & n3053 ) | ( n2989 & n3063 ) | ( n3053 & n3063 ) ;
  assign n3066 = ( n3053 & n3064 ) | ( n3053 & ~n3065 ) | ( n3064 & ~n3065 ) ;
  assign n3067 = ~n553 & n1947 ;
  assign n3068 = n222 & n3067 ;
  assign n3069 = n1941 & n2635 ;
  assign n3070 = n1944 & n2661 ;
  assign n3071 = n3069 | n3070 ;
  assign n3072 = n238 | n3071 ;
  assign n3073 = ( ~n2768 & n3071 ) | ( ~n2768 & n3072 ) | ( n3071 & n3072 ) ;
  assign n3074 = ( ~n222 & n3067 ) | ( ~n222 & n3073 ) | ( n3067 & n3073 ) ;
  assign n3075 = n222 & ~n3073 ;
  assign n3076 = ( ~n3068 & n3074 ) | ( ~n3068 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = n2844 | n2857 ;
  assign n3078 = n2389 & ~n2857 ;
  assign n3079 = ( n231 & n2313 ) | ( n231 & n3077 ) | ( n2313 & n3077 ) ;
  assign n3080 = ( ~n3077 & n3078 ) | ( ~n3077 & n3079 ) | ( n3078 & n3079 ) ;
  assign n3081 = n2313 & ~n3079 ;
  assign n3082 = ( n231 & ~n3080 ) | ( n231 & n3081 ) | ( ~n3080 & n3081 ) ;
  assign n3083 = ( ~n3066 & n3076 ) | ( ~n3066 & n3082 ) | ( n3076 & n3082 ) ;
  assign n3084 = ( n3066 & n3076 ) | ( n3066 & n3082 ) | ( n3076 & n3082 ) ;
  assign n3085 = ( n3066 & n3083 ) | ( n3066 & ~n3084 ) | ( n3083 & ~n3084 ) ;
  assign n3086 = ( n3003 & n3005 ) | ( n3003 & n3085 ) | ( n3005 & n3085 ) ;
  assign n3087 = ( n3003 & ~n3005 ) | ( n3003 & n3085 ) | ( ~n3005 & n3085 ) ;
  assign n3088 = ( n3005 & ~n3086 ) | ( n3005 & n3087 ) | ( ~n3086 & n3087 ) ;
  assign n3089 = n166 | n742 ;
  assign n3090 = n2561 | n2927 ;
  assign n3091 = n3089 | n3090 ;
  assign n3092 = n296 | n3091 ;
  assign n3093 = n114 | n485 ;
  assign n3094 = n193 | n3093 ;
  assign n3095 = n528 | n854 ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = n3092 | n3096 ;
  assign n3098 = n704 | n1626 ;
  assign n3099 = n1189 | n3098 ;
  assign n3100 = n3097 | n3099 ;
  assign n3101 = ( n3023 & ~n3088 ) | ( n3023 & n3100 ) | ( ~n3088 & n3100 ) ;
  assign n3102 = ( n3023 & n3088 ) | ( n3023 & n3100 ) | ( n3088 & n3100 ) ;
  assign n3103 = ( n3088 & n3101 ) | ( n3088 & ~n3102 ) | ( n3101 & ~n3102 ) ;
  assign n3104 = n3025 | n3103 ;
  assign n3105 = n2837 & n2940 ;
  assign n3106 = n3024 & n3105 ;
  assign n3107 = n2842 | n3106 ;
  assign n3108 = ( n3025 & ~n3103 ) | ( n3025 & n3107 ) | ( ~n3103 & n3107 ) ;
  assign n3109 = ~n3103 & n3107 ;
  assign n3110 = ( n3104 & ~n3108 ) | ( n3104 & n3109 ) | ( ~n3108 & n3109 ) ;
  assign n3111 = n1947 & ~n2857 ;
  assign n3112 = ~n553 & n1944 ;
  assign n3113 = n3111 | n3112 ;
  assign n3114 = n1941 & n2661 ;
  assign n3115 = n3113 | n3114 ;
  assign n3116 = n238 | n3115 ;
  assign n3117 = ( n2861 & n3115 ) | ( n2861 & n3116 ) | ( n3115 & n3116 ) ;
  assign n3118 = n222 & ~n3117 ;
  assign n3119 = ~n222 & n3117 ;
  assign n3120 = n3118 | n3119 ;
  assign n3121 = n1994 & ~n2365 ;
  assign n3122 = n1991 & n2367 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = n1997 & n2635 ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = ( n1985 & ~n2640 ) | ( n1985 & n3125 ) | ( ~n2640 & n3125 ) ;
  assign n3127 = n902 | n3125 ;
  assign n3128 = ~n3126 & n3127 ;
  assign n3129 = ( ~n3125 & n3126 ) | ( ~n3125 & n3127 ) | ( n3126 & n3127 ) ;
  assign n3130 = ( ~n902 & n3128 ) | ( ~n902 & n3129 ) | ( n3128 & n3129 ) ;
  assign n3131 = n1921 & n2023 ;
  assign n3132 = ~n1893 & n2026 ;
  assign n3133 = n3131 | n3132 ;
  assign n3134 = n2012 & n2369 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = ( n2011 & ~n2410 ) | ( n2011 & n3135 ) | ( ~n2410 & n3135 ) ;
  assign n3137 = n646 & ~n3135 ;
  assign n3138 = n3136 | n3137 ;
  assign n3139 = ( n3135 & ~n3136 ) | ( n3135 & n3137 ) | ( ~n3136 & n3137 ) ;
  assign n3140 = ( ~n646 & n3138 ) | ( ~n646 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3141 = ( ~n1899 & n3038 ) | ( ~n1899 & n3046 ) | ( n3038 & n3046 ) ;
  assign n3142 = n584 & ~n3141 ;
  assign n3143 = n584 & ~n1897 ;
  assign n3144 = ~n1914 & n2282 ;
  assign n3145 = n1895 & n2236 ;
  assign n3146 = n3144 | n3145 ;
  assign n3147 = n1918 & n2241 ;
  assign n3148 = n3146 | n3147 ;
  assign n3149 = n1971 & n2238 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = ( n231 & n3143 ) | ( n231 & ~n3150 ) | ( n3143 & ~n3150 ) ;
  assign n3152 = ( ~n231 & n3143 ) | ( ~n231 & n3150 ) | ( n3143 & n3150 ) ;
  assign n3153 = ( ~n3143 & n3151 ) | ( ~n3143 & n3152 ) | ( n3151 & n3152 ) ;
  assign n3154 = ( n3140 & n3142 ) | ( n3140 & n3153 ) | ( n3142 & n3153 ) ;
  assign n3155 = ( ~n3140 & n3142 ) | ( ~n3140 & n3153 ) | ( n3142 & n3153 ) ;
  assign n3156 = ( n3140 & ~n3154 ) | ( n3140 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = ( n3051 & n3130 ) | ( n3051 & n3156 ) | ( n3130 & n3156 ) ;
  assign n3158 = ( ~n3051 & n3130 ) | ( ~n3051 & n3156 ) | ( n3130 & n3156 ) ;
  assign n3159 = ( n3051 & ~n3157 ) | ( n3051 & n3158 ) | ( ~n3157 & n3158 ) ;
  assign n3160 = ( n3065 & n3120 ) | ( n3065 & n3159 ) | ( n3120 & n3159 ) ;
  assign n3161 = ( ~n3065 & n3120 ) | ( ~n3065 & n3159 ) | ( n3120 & n3159 ) ;
  assign n3162 = ( n3065 & ~n3160 ) | ( n3065 & n3161 ) | ( ~n3160 & n3161 ) ;
  assign n3163 = ( n3084 & n3086 ) | ( n3084 & n3162 ) | ( n3086 & n3162 ) ;
  assign n3164 = ( n3084 & ~n3086 ) | ( n3084 & n3162 ) | ( ~n3086 & n3162 ) ;
  assign n3165 = ( n3086 & ~n3163 ) | ( n3086 & n3164 ) | ( ~n3163 & n3164 ) ;
  assign n3166 = n198 | n1590 ;
  assign n3167 = n1775 | n3166 ;
  assign n3168 = n300 | n362 ;
  assign n3169 = n197 | n3168 ;
  assign n3170 = n407 | n3169 ;
  assign n3171 = n3167 | n3170 ;
  assign n3172 = n894 | n3171 ;
  assign n3173 = n685 | n3172 ;
  assign n3174 = n1835 | n3173 ;
  assign n3175 = ( n3102 & ~n3165 ) | ( n3102 & n3174 ) | ( ~n3165 & n3174 ) ;
  assign n3176 = ( n3102 & n3165 ) | ( n3102 & n3174 ) | ( n3165 & n3174 ) ;
  assign n3177 = ( n3165 & n3175 ) | ( n3165 & ~n3176 ) | ( n3175 & ~n3176 ) ;
  assign n3178 = n3107 | n3177 ;
  assign n3179 = ( n2842 & n3103 ) | ( n2842 & n3104 ) | ( n3103 & n3104 ) ;
  assign n3180 = ( n3107 & ~n3177 ) | ( n3107 & n3179 ) | ( ~n3177 & n3179 ) ;
  assign n3181 = ~n3177 & n3179 ;
  assign n3182 = ( n3178 & ~n3180 ) | ( n3178 & n3181 ) | ( ~n3180 & n3181 ) ;
  assign n3183 = n584 | n3150 ;
  assign n3184 = ~n3152 & n3183 ;
  assign n3185 = n584 & ~n1914 ;
  assign n3186 = ( ~n231 & n3184 ) | ( ~n231 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3187 = ( n231 & n3184 ) | ( n231 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3188 = ( n231 & n3186 ) | ( n231 & ~n3187 ) | ( n3186 & ~n3187 ) ;
  assign n3189 = ~n1893 & n2023 ;
  assign n3190 = n2026 & n2369 ;
  assign n3191 = n3189 | n3190 ;
  assign n3192 = n2012 & n2367 ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = ( n2011 & n2394 ) | ( n2011 & n3193 ) | ( n2394 & n3193 ) ;
  assign n3195 = n646 & ~n3193 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = ( n3193 & ~n3194 ) | ( n3193 & n3195 ) | ( ~n3194 & n3195 ) ;
  assign n3198 = ( ~n646 & n3196 ) | ( ~n646 & n3197 ) | ( n3196 & n3197 ) ;
  assign n3199 = n1895 & n2282 ;
  assign n3200 = n1918 & n2236 ;
  assign n3201 = n3199 | n3200 ;
  assign n3202 = n1921 & n2241 ;
  assign n3203 = n3201 | n3202 ;
  assign n3204 = ( n1958 & n2238 ) | ( n1958 & n3203 ) | ( n2238 & n3203 ) ;
  assign n3205 = n584 | n3203 ;
  assign n3206 = ~n3204 & n3205 ;
  assign n3207 = ( ~n3203 & n3204 ) | ( ~n3203 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3208 = ( ~n584 & n3206 ) | ( ~n584 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3209 = ( n3188 & n3198 ) | ( n3188 & n3208 ) | ( n3198 & n3208 ) ;
  assign n3210 = ( ~n3188 & n3198 ) | ( ~n3188 & n3208 ) | ( n3198 & n3208 ) ;
  assign n3211 = ( n3188 & ~n3209 ) | ( n3188 & n3210 ) | ( ~n3209 & n3210 ) ;
  assign n3212 = n1991 & ~n2365 ;
  assign n3213 = n1994 & n2635 ;
  assign n3214 = n3212 | n3213 ;
  assign n3215 = n1997 & n2661 ;
  assign n3216 = n3214 | n3215 ;
  assign n3217 = ( n1985 & n2667 ) | ( n1985 & n3216 ) | ( n2667 & n3216 ) ;
  assign n3218 = n902 | n3216 ;
  assign n3219 = ~n3217 & n3218 ;
  assign n3220 = ( ~n3216 & n3217 ) | ( ~n3216 & n3218 ) | ( n3217 & n3218 ) ;
  assign n3221 = ( ~n902 & n3219 ) | ( ~n902 & n3220 ) | ( n3219 & n3220 ) ;
  assign n3222 = ( n3154 & ~n3211 ) | ( n3154 & n3221 ) | ( ~n3211 & n3221 ) ;
  assign n3223 = ( n3154 & n3211 ) | ( n3154 & n3221 ) | ( n3211 & n3221 ) ;
  assign n3224 = ( n3211 & n3222 ) | ( n3211 & ~n3223 ) | ( n3222 & ~n3223 ) ;
  assign n3225 = n1944 & ~n2857 ;
  assign n3226 = n222 & n3225 ;
  assign n3227 = ~n553 & n1941 ;
  assign n3228 = n238 | n3227 ;
  assign n3229 = ( n2945 & n3227 ) | ( n2945 & n3228 ) | ( n3227 & n3228 ) ;
  assign n3230 = ( ~n222 & n3225 ) | ( ~n222 & n3229 ) | ( n3225 & n3229 ) ;
  assign n3231 = n222 & ~n3229 ;
  assign n3232 = ( ~n3226 & n3230 ) | ( ~n3226 & n3231 ) | ( n3230 & n3231 ) ;
  assign n3233 = ( n3157 & n3224 ) | ( n3157 & n3232 ) | ( n3224 & n3232 ) ;
  assign n3234 = ( n3157 & ~n3224 ) | ( n3157 & n3232 ) | ( ~n3224 & n3232 ) ;
  assign n3235 = ( n3224 & ~n3233 ) | ( n3224 & n3234 ) | ( ~n3233 & n3234 ) ;
  assign n3236 = ( n3160 & ~n3163 ) | ( n3160 & n3235 ) | ( ~n3163 & n3235 ) ;
  assign n3237 = ( n3160 & n3163 ) | ( n3160 & n3235 ) | ( n3163 & n3235 ) ;
  assign n3238 = ( n3163 & n3236 ) | ( n3163 & ~n3237 ) | ( n3236 & ~n3237 ) ;
  assign n3239 = n150 | n947 ;
  assign n3240 = n612 | n3239 ;
  assign n3241 = n497 | n529 ;
  assign n3242 = n3240 | n3241 ;
  assign n3243 = n164 | n1778 ;
  assign n3244 = n1875 | n2928 ;
  assign n3245 = n3243 | n3244 ;
  assign n3246 = n3242 | n3245 ;
  assign n3247 = n2351 | n2851 ;
  assign n3248 = n3246 | n3247 ;
  assign n3249 = ( ~n3176 & n3238 ) | ( ~n3176 & n3248 ) | ( n3238 & n3248 ) ;
  assign n3250 = ( n3176 & n3238 ) | ( n3176 & n3248 ) | ( n3238 & n3248 ) ;
  assign n3251 = ( n3176 & n3249 ) | ( n3176 & ~n3250 ) | ( n3249 & ~n3250 ) ;
  assign n3252 = n3103 & n3106 ;
  assign n3253 = n3177 & n3252 ;
  assign n3254 = n3177 | n3179 ;
  assign n3255 = n2842 | n3253 ;
  assign n3256 = ( n3253 & n3254 ) | ( n3253 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3257 = n3251 & ~n3256 ;
  assign n3258 = ~n3251 & n3256 ;
  assign n3259 = n3257 | n3258 ;
  assign n3260 = n3251 & n3253 ;
  assign n3261 = n2842 | n3260 ;
  assign n3262 = n238 & ~n3077 ;
  assign n3263 = n1941 & ~n2857 ;
  assign n3264 = ( ~n222 & n3262 ) | ( ~n222 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3265 = ( n222 & n3262 ) | ( n222 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3266 = ( n222 & n3264 ) | ( n222 & ~n3265 ) | ( n3264 & ~n3265 ) ;
  assign n3267 = n1994 & n2661 ;
  assign n3268 = ~n553 & n1997 ;
  assign n3269 = n3267 | n3268 ;
  assign n3270 = n1991 & n2635 ;
  assign n3271 = n3269 | n3270 ;
  assign n3272 = ( n1985 & ~n2768 ) | ( n1985 & n3271 ) | ( ~n2768 & n3271 ) ;
  assign n3273 = n902 & ~n3271 ;
  assign n3274 = n3272 | n3273 ;
  assign n3275 = ( n3271 & ~n3272 ) | ( n3271 & n3273 ) | ( ~n3272 & n3273 ) ;
  assign n3276 = ( ~n902 & n3274 ) | ( ~n902 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3277 = n584 & n1895 ;
  assign n3278 = ( n231 & n3187 ) | ( n231 & ~n3277 ) | ( n3187 & ~n3277 ) ;
  assign n3279 = ( n231 & ~n3187 ) | ( n231 & n3277 ) | ( ~n3187 & n3277 ) ;
  assign n3280 = ( ~n231 & n3278 ) | ( ~n231 & n3279 ) | ( n3278 & n3279 ) ;
  assign n3281 = n2023 & n2369 ;
  assign n3282 = n2026 & n2367 ;
  assign n3283 = n3281 | n3282 ;
  assign n3284 = n2012 & ~n2365 ;
  assign n3285 = n3283 | n3284 ;
  assign n3286 = ( n2011 & ~n2379 ) | ( n2011 & n3285 ) | ( ~n2379 & n3285 ) ;
  assign n3287 = n646 & ~n3285 ;
  assign n3288 = n3286 | n3287 ;
  assign n3289 = ( n3285 & ~n3286 ) | ( n3285 & n3287 ) | ( ~n3286 & n3287 ) ;
  assign n3290 = ( ~n646 & n3288 ) | ( ~n646 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = n1918 & n2282 ;
  assign n3292 = n1921 & n2236 ;
  assign n3293 = n3291 | n3292 ;
  assign n3294 = ~n1893 & n2241 ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = ( ~n1938 & n2238 ) | ( ~n1938 & n3295 ) | ( n2238 & n3295 ) ;
  assign n3297 = n584 & ~n3295 ;
  assign n3298 = n3296 | n3297 ;
  assign n3299 = ( n3295 & ~n3296 ) | ( n3295 & n3297 ) | ( ~n3296 & n3297 ) ;
  assign n3300 = ( ~n584 & n3298 ) | ( ~n584 & n3299 ) | ( n3298 & n3299 ) ;
  assign n3301 = ( n3280 & n3290 ) | ( n3280 & n3300 ) | ( n3290 & n3300 ) ;
  assign n3302 = ( ~n3280 & n3290 ) | ( ~n3280 & n3300 ) | ( n3290 & n3300 ) ;
  assign n3303 = ( n3280 & ~n3301 ) | ( n3280 & n3302 ) | ( ~n3301 & n3302 ) ;
  assign n3304 = ( n3209 & ~n3276 ) | ( n3209 & n3303 ) | ( ~n3276 & n3303 ) ;
  assign n3305 = ( n3209 & n3276 ) | ( n3209 & n3303 ) | ( n3276 & n3303 ) ;
  assign n3306 = ( n3276 & n3304 ) | ( n3276 & ~n3305 ) | ( n3304 & ~n3305 ) ;
  assign n3307 = ( ~n3223 & n3266 ) | ( ~n3223 & n3306 ) | ( n3266 & n3306 ) ;
  assign n3308 = ( n3223 & n3266 ) | ( n3223 & n3306 ) | ( n3266 & n3306 ) ;
  assign n3309 = ( n3223 & n3307 ) | ( n3223 & ~n3308 ) | ( n3307 & ~n3308 ) ;
  assign n3310 = ( n3233 & n3237 ) | ( n3233 & n3309 ) | ( n3237 & n3309 ) ;
  assign n3311 = ( n3233 & ~n3237 ) | ( n3233 & n3309 ) | ( ~n3237 & n3309 ) ;
  assign n3312 = ( n3237 & ~n3310 ) | ( n3237 & n3311 ) | ( ~n3310 & n3311 ) ;
  assign n3313 = n260 | n495 ;
  assign n3314 = n2852 | n3313 ;
  assign n3315 = n1777 | n3314 ;
  assign n3316 = n213 | n594 ;
  assign n3317 = n1858 | n3316 ;
  assign n3318 = n2560 | n3317 ;
  assign n3319 = n1826 | n3318 ;
  assign n3320 = n3315 | n3319 ;
  assign n3321 = n180 | n287 ;
  assign n3322 = n320 | n3321 ;
  assign n3323 = n1824 | n3322 ;
  assign n3324 = n344 | n626 ;
  assign n3325 = n889 | n1686 ;
  assign n3326 = n3324 | n3325 ;
  assign n3327 = n3323 | n3326 ;
  assign n3328 = n3320 | n3327 ;
  assign n3329 = n2747 | n3328 ;
  assign n3330 = ( n3250 & ~n3312 ) | ( n3250 & n3329 ) | ( ~n3312 & n3329 ) ;
  assign n3331 = ( n3250 & n3312 ) | ( n3250 & n3329 ) | ( n3312 & n3329 ) ;
  assign n3332 = ( n3312 & n3330 ) | ( n3312 & ~n3331 ) | ( n3330 & ~n3331 ) ;
  assign n3333 = n3261 | n3332 ;
  assign n3334 = n3251 | n3254 ;
  assign n3335 = ( n3261 & ~n3332 ) | ( n3261 & n3334 ) | ( ~n3332 & n3334 ) ;
  assign n3336 = ~n3332 & n3334 ;
  assign n3337 = ( n3333 & ~n3335 ) | ( n3333 & n3336 ) | ( ~n3335 & n3336 ) ;
  assign n3338 = n3260 & n3332 ;
  assign n3339 = n3332 | n3334 ;
  assign n3340 = n2842 | n3338 ;
  assign n3341 = ( n3338 & n3339 ) | ( n3338 & n3340 ) | ( n3339 & n3340 ) ;
  assign n3342 = n1997 & ~n2857 ;
  assign n3343 = ~n553 & n1994 ;
  assign n3344 = n3342 | n3343 ;
  assign n3345 = n1991 & n2661 ;
  assign n3346 = n3344 | n3345 ;
  assign n3347 = ( n1985 & n2861 ) | ( n1985 & n3346 ) | ( n2861 & n3346 ) ;
  assign n3348 = n902 | n3346 ;
  assign n3349 = ~n3347 & n3348 ;
  assign n3350 = ( ~n3346 & n3347 ) | ( ~n3346 & n3348 ) | ( n3347 & n3348 ) ;
  assign n3351 = ( ~n902 & n3349 ) | ( ~n902 & n3350 ) | ( n3349 & n3350 ) ;
  assign n3352 = n2011 & ~n2640 ;
  assign n3353 = n646 & n3352 ;
  assign n3354 = n2026 & ~n2365 ;
  assign n3355 = n2023 & n2367 ;
  assign n3356 = n3354 | n3355 ;
  assign n3357 = n2012 & n2635 ;
  assign n3358 = n3356 | n3357 ;
  assign n3359 = ( ~n646 & n3352 ) | ( ~n646 & n3358 ) | ( n3352 & n3358 ) ;
  assign n3360 = n646 & ~n3358 ;
  assign n3361 = ( ~n3353 & n3359 ) | ( ~n3353 & n3360 ) | ( n3359 & n3360 ) ;
  assign n3362 = ( n231 & n3187 ) | ( n231 & n3277 ) | ( n3187 & n3277 ) ;
  assign n3363 = n1921 & n2282 ;
  assign n3364 = ~n1893 & n2236 ;
  assign n3365 = n3363 | n3364 ;
  assign n3366 = n2241 & n2369 ;
  assign n3367 = n3365 | n3366 ;
  assign n3368 = ( n2238 & ~n2410 ) | ( n2238 & n3367 ) | ( ~n2410 & n3367 ) ;
  assign n3369 = n584 | n3367 ;
  assign n3370 = ~n3368 & n3369 ;
  assign n3371 = ( ~n3367 & n3368 ) | ( ~n3367 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3372 = ( ~n584 & n3370 ) | ( ~n584 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3373 = n584 & n1918 ;
  assign n3374 = ( n222 & ~n231 ) | ( n222 & n3373 ) | ( ~n231 & n3373 ) ;
  assign n3375 = ( n222 & n231 ) | ( n222 & ~n3373 ) | ( n231 & ~n3373 ) ;
  assign n3376 = ( ~n222 & n3374 ) | ( ~n222 & n3375 ) | ( n3374 & n3375 ) ;
  assign n3377 = ( n3362 & n3372 ) | ( n3362 & n3376 ) | ( n3372 & n3376 ) ;
  assign n3378 = ( ~n3362 & n3372 ) | ( ~n3362 & n3376 ) | ( n3372 & n3376 ) ;
  assign n3379 = ( n3362 & ~n3377 ) | ( n3362 & n3378 ) | ( ~n3377 & n3378 ) ;
  assign n3380 = ( n3301 & n3361 ) | ( n3301 & n3379 ) | ( n3361 & n3379 ) ;
  assign n3381 = ( ~n3301 & n3361 ) | ( ~n3301 & n3379 ) | ( n3361 & n3379 ) ;
  assign n3382 = ( n3301 & ~n3380 ) | ( n3301 & n3381 ) | ( ~n3380 & n3381 ) ;
  assign n3383 = ( n3305 & n3351 ) | ( n3305 & n3382 ) | ( n3351 & n3382 ) ;
  assign n3384 = ( ~n3305 & n3351 ) | ( ~n3305 & n3382 ) | ( n3351 & n3382 ) ;
  assign n3385 = ( n3305 & ~n3383 ) | ( n3305 & n3384 ) | ( ~n3383 & n3384 ) ;
  assign n3386 = ( n3308 & n3310 ) | ( n3308 & n3385 ) | ( n3310 & n3385 ) ;
  assign n3387 = ( n3308 & ~n3310 ) | ( n3308 & n3385 ) | ( ~n3310 & n3385 ) ;
  assign n3388 = ( n3310 & ~n3386 ) | ( n3310 & n3387 ) | ( ~n3386 & n3387 ) ;
  assign n3389 = n845 | n2546 ;
  assign n3390 = n504 | n3389 ;
  assign n3391 = n200 | n689 ;
  assign n3392 = n159 | n328 ;
  assign n3393 = n3243 | n3392 ;
  assign n3394 = n3391 | n3393 ;
  assign n3395 = n3390 | n3394 ;
  assign n3396 = n3320 | n3395 ;
  assign n3397 = n1704 | n3396 ;
  assign n3398 = ( n3331 & ~n3388 ) | ( n3331 & n3397 ) | ( ~n3388 & n3397 ) ;
  assign n3399 = ( n3331 & n3388 ) | ( n3331 & n3397 ) | ( n3388 & n3397 ) ;
  assign n3400 = ( n3388 & n3398 ) | ( n3388 & ~n3399 ) | ( n3398 & ~n3399 ) ;
  assign n3401 = ~n3341 & n3400 ;
  assign n3402 = n3341 & ~n3400 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = n3338 & n3400 ;
  assign n3405 = ~n553 & n1991 ;
  assign n3406 = n1985 | n3405 ;
  assign n3407 = ( n2945 & n3405 ) | ( n2945 & n3406 ) | ( n3405 & n3406 ) ;
  assign n3408 = n1994 & ~n2857 ;
  assign n3409 = ( ~n902 & n3407 ) | ( ~n902 & n3408 ) | ( n3407 & n3408 ) ;
  assign n3410 = n902 & ~n3407 ;
  assign n3411 = ( n902 & n3407 ) | ( n902 & n3408 ) | ( n3407 & n3408 ) ;
  assign n3412 = ( n3409 & n3410 ) | ( n3409 & ~n3411 ) | ( n3410 & ~n3411 ) ;
  assign n3413 = n2011 & n2667 ;
  assign n3414 = n646 & n3413 ;
  assign n3415 = n2023 & ~n2365 ;
  assign n3416 = n2026 & n2635 ;
  assign n3417 = n3415 | n3416 ;
  assign n3418 = n2012 & n2661 ;
  assign n3419 = n3417 | n3418 ;
  assign n3420 = ( ~n646 & n3413 ) | ( ~n646 & n3419 ) | ( n3413 & n3419 ) ;
  assign n3421 = n646 & ~n3419 ;
  assign n3422 = ( ~n3414 & n3420 ) | ( ~n3414 & n3421 ) | ( n3420 & n3421 ) ;
  assign n3423 = n584 & ~n1921 ;
  assign n3424 = ~n1893 & n2282 ;
  assign n3425 = n2236 & n2369 ;
  assign n3426 = n3424 | n3425 ;
  assign n3427 = n2241 & n2367 ;
  assign n3428 = n3426 | n3427 ;
  assign n3429 = n2238 & n2394 ;
  assign n3430 = n3428 | n3429 ;
  assign n3431 = ( n3375 & n3423 ) | ( n3375 & n3430 ) | ( n3423 & n3430 ) ;
  assign n3432 = ( n3375 & ~n3423 ) | ( n3375 & n3430 ) | ( ~n3423 & n3430 ) ;
  assign n3433 = ( n3423 & ~n3431 ) | ( n3423 & n3432 ) | ( ~n3431 & n3432 ) ;
  assign n3434 = ( n3377 & ~n3422 ) | ( n3377 & n3433 ) | ( ~n3422 & n3433 ) ;
  assign n3435 = ( n3377 & n3422 ) | ( n3377 & n3433 ) | ( n3422 & n3433 ) ;
  assign n3436 = ( n3422 & n3434 ) | ( n3422 & ~n3435 ) | ( n3434 & ~n3435 ) ;
  assign n3437 = ( n3380 & n3412 ) | ( n3380 & n3436 ) | ( n3412 & n3436 ) ;
  assign n3438 = ( ~n3380 & n3412 ) | ( ~n3380 & n3436 ) | ( n3412 & n3436 ) ;
  assign n3439 = ( n3380 & ~n3437 ) | ( n3380 & n3438 ) | ( ~n3437 & n3438 ) ;
  assign n3440 = ( n3383 & n3386 ) | ( n3383 & n3439 ) | ( n3386 & n3439 ) ;
  assign n3441 = ( n3383 & ~n3386 ) | ( n3383 & n3439 ) | ( ~n3386 & n3439 ) ;
  assign n3442 = ( n3386 & ~n3440 ) | ( n3386 & n3441 ) | ( ~n3440 & n3441 ) ;
  assign n3443 = n877 | n882 ;
  assign n3444 = n112 | n146 ;
  assign n3445 = n1613 | n3444 ;
  assign n3446 = n354 | n360 ;
  assign n3447 = n298 | n3446 ;
  assign n3448 = n3445 | n3447 ;
  assign n3449 = n1850 | n3448 ;
  assign n3450 = n3443 | n3449 ;
  assign n3451 = n491 | n3450 ;
  assign n3452 = n2555 | n3451 ;
  assign n3453 = ( n3399 & ~n3442 ) | ( n3399 & n3452 ) | ( ~n3442 & n3452 ) ;
  assign n3454 = ( n3399 & n3442 ) | ( n3399 & n3452 ) | ( n3442 & n3452 ) ;
  assign n3455 = ( n3442 & n3453 ) | ( n3442 & ~n3454 ) | ( n3453 & ~n3454 ) ;
  assign n3456 = n3404 & ~n3455 ;
  assign n3457 = n3339 | n3400 ;
  assign n3458 = n2842 & n3457 ;
  assign n3459 = ( n3404 & n3455 ) | ( n3404 & n3458 ) | ( n3455 & n3458 ) ;
  assign n3460 = n3455 | n3458 ;
  assign n3461 = ( n3456 & ~n3459 ) | ( n3456 & n3460 ) | ( ~n3459 & n3460 ) ;
  assign n3462 = ( n2842 & n3340 ) | ( n2842 & n3400 ) | ( n3340 & n3400 ) ;
  assign n3463 = ( n3455 & n3458 ) | ( n3455 & n3462 ) | ( n3458 & n3462 ) ;
  assign n3464 = n2023 & n2635 ;
  assign n3465 = n2026 & n2661 ;
  assign n3466 = n3464 | n3465 ;
  assign n3467 = ~n553 & n2012 ;
  assign n3468 = n3466 | n3467 ;
  assign n3469 = ( n2011 & ~n2768 ) | ( n2011 & n3468 ) | ( ~n2768 & n3468 ) ;
  assign n3470 = n646 & ~n3468 ;
  assign n3471 = n3469 | n3470 ;
  assign n3472 = ( n3468 & ~n3469 ) | ( n3468 & n3470 ) | ( ~n3469 & n3470 ) ;
  assign n3473 = ( ~n646 & n3471 ) | ( ~n646 & n3472 ) | ( n3471 & n3472 ) ;
  assign n3474 = ( n584 & n1893 ) | ( n584 & n1921 ) | ( n1893 & n1921 ) ;
  assign n3475 = n2282 & n2369 ;
  assign n3476 = n2236 & n2367 ;
  assign n3477 = n3475 | n3476 ;
  assign n3478 = n2241 & ~n2365 ;
  assign n3479 = n3477 | n3478 ;
  assign n3480 = n2238 & ~n2379 ;
  assign n3481 = n3479 | n3480 ;
  assign n3482 = n1893 & n1921 ;
  assign n3483 = ( ~n3474 & n3481 ) | ( ~n3474 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3484 = ( n3474 & n3481 ) | ( n3474 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3485 = ( n3474 & n3483 ) | ( n3474 & ~n3484 ) | ( n3483 & ~n3484 ) ;
  assign n3486 = ~n584 & n3430 ;
  assign n3487 = n3432 & ~n3486 ;
  assign n3488 = ( n3473 & n3485 ) | ( n3473 & n3487 ) | ( n3485 & n3487 ) ;
  assign n3489 = ( ~n3473 & n3485 ) | ( ~n3473 & n3487 ) | ( n3485 & n3487 ) ;
  assign n3490 = ( n3473 & ~n3488 ) | ( n3473 & n3489 ) | ( ~n3488 & n3489 ) ;
  assign n3491 = ( n1985 & ~n2857 ) | ( n1985 & n2858 ) | ( ~n2857 & n2858 ) ;
  assign n3492 = ( n1991 & ~n3077 ) | ( n1991 & n3491 ) | ( ~n3077 & n3491 ) ;
  assign n3493 = n902 & ~n3492 ;
  assign n3494 = ~n902 & n3492 ;
  assign n3495 = n3493 | n3494 ;
  assign n3496 = ( n3435 & ~n3490 ) | ( n3435 & n3495 ) | ( ~n3490 & n3495 ) ;
  assign n3497 = ( n3435 & n3490 ) | ( n3435 & n3495 ) | ( n3490 & n3495 ) ;
  assign n3498 = ( n3490 & n3496 ) | ( n3490 & ~n3497 ) | ( n3496 & ~n3497 ) ;
  assign n3499 = ( n3437 & n3440 ) | ( n3437 & n3498 ) | ( n3440 & n3498 ) ;
  assign n3500 = ( n3437 & ~n3440 ) | ( n3437 & n3498 ) | ( ~n3440 & n3498 ) ;
  assign n3501 = ( n3440 & ~n3499 ) | ( n3440 & n3500 ) | ( ~n3499 & n3500 ) ;
  assign n3502 = n129 | n252 ;
  assign n3503 = n114 | n3502 ;
  assign n3504 = n2339 | n3503 ;
  assign n3505 = n1677 | n1810 ;
  assign n3506 = n200 | n3324 ;
  assign n3507 = n3505 | n3506 ;
  assign n3508 = n3504 | n3507 ;
  assign n3509 = n718 | n3508 ;
  assign n3510 = n2758 | n3509 ;
  assign n3511 = n1781 | n3510 ;
  assign n3512 = ( n3454 & ~n3501 ) | ( n3454 & n3511 ) | ( ~n3501 & n3511 ) ;
  assign n3513 = ( n3454 & n3501 ) | ( n3454 & n3511 ) | ( n3501 & n3511 ) ;
  assign n3514 = ( n3501 & n3512 ) | ( n3501 & ~n3513 ) | ( n3512 & ~n3513 ) ;
  assign n3515 = n3463 | n3514 ;
  assign n3516 = n3463 & n3514 ;
  assign n3517 = n3515 & ~n3516 ;
  assign n3518 = n3404 & n3455 ;
  assign n3519 = n3514 & n3518 ;
  assign n3520 = ~n1893 & n3423 ;
  assign n3521 = n2238 & ~n2640 ;
  assign n3522 = n2241 & n2635 ;
  assign n3523 = n2282 & n2367 ;
  assign n3524 = n3522 | n3523 ;
  assign n3525 = n2236 & ~n2365 ;
  assign n3526 = n3524 | n3525 ;
  assign n3527 = n3521 | n3526 ;
  assign n3528 = n3520 & n3527 ;
  assign n3529 = n584 & n1921 ;
  assign n3530 = n1893 & n3529 ;
  assign n3531 = n3481 | n3530 ;
  assign n3532 = ( ~n3520 & n3527 ) | ( ~n3520 & n3531 ) | ( n3527 & n3531 ) ;
  assign n3533 = n3527 & n3531 ;
  assign n3534 = ( n3528 & n3532 ) | ( n3528 & ~n3533 ) | ( n3532 & ~n3533 ) ;
  assign n3535 = ( n1891 & n2325 ) | ( n1891 & n3423 ) | ( n2325 & n3423 ) ;
  assign n3536 = ( n1891 & n2325 ) | ( n1891 & ~n3423 ) | ( n2325 & ~n3423 ) ;
  assign n3537 = ( n3529 & n3535 ) | ( n3529 & ~n3536 ) | ( n3535 & ~n3536 ) ;
  assign n3538 = ( n902 & ~n3534 ) | ( n902 & n3537 ) | ( ~n3534 & n3537 ) ;
  assign n3539 = ( n902 & n3534 ) | ( n902 & ~n3537 ) | ( n3534 & ~n3537 ) ;
  assign n3540 = ( ~n902 & n3538 ) | ( ~n902 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3541 = n2012 & ~n2857 ;
  assign n3542 = ~n553 & n2026 ;
  assign n3543 = n3541 | n3542 ;
  assign n3544 = n2023 & n2661 ;
  assign n3545 = n3543 | n3544 ;
  assign n3546 = ( n2011 & n2861 ) | ( n2011 & n3545 ) | ( n2861 & n3545 ) ;
  assign n3547 = n646 | n3545 ;
  assign n3548 = ~n3546 & n3547 ;
  assign n3549 = ( ~n3545 & n3546 ) | ( ~n3545 & n3547 ) | ( n3546 & n3547 ) ;
  assign n3550 = ( ~n646 & n3548 ) | ( ~n646 & n3549 ) | ( n3548 & n3549 ) ;
  assign n3551 = ( n3489 & n3540 ) | ( n3489 & ~n3550 ) | ( n3540 & ~n3550 ) ;
  assign n3552 = ( ~n3489 & n3540 ) | ( ~n3489 & n3550 ) | ( n3540 & n3550 ) ;
  assign n3553 = ( ~n3540 & n3551 ) | ( ~n3540 & n3552 ) | ( n3551 & n3552 ) ;
  assign n3554 = ( n3497 & n3499 ) | ( n3497 & n3553 ) | ( n3499 & n3553 ) ;
  assign n3555 = ( n3497 & ~n3499 ) | ( n3497 & n3553 ) | ( ~n3499 & n3553 ) ;
  assign n3556 = ( n3499 & ~n3554 ) | ( n3499 & n3555 ) | ( ~n3554 & n3555 ) ;
  assign n3557 = n597 | n669 ;
  assign n3558 = n3324 | n3557 ;
  assign n3559 = n2748 | n3558 ;
  assign n3560 = n140 | n173 ;
  assign n3561 = n291 | n3560 ;
  assign n3562 = n744 | n3561 ;
  assign n3563 = n2852 | n3562 ;
  assign n3564 = n3559 | n3563 ;
  assign n3565 = n432 | n2562 ;
  assign n3566 = n968 | n3565 ;
  assign n3567 = n3564 | n3566 ;
  assign n3568 = ( n3513 & ~n3556 ) | ( n3513 & n3567 ) | ( ~n3556 & n3567 ) ;
  assign n3569 = ( n3513 & n3556 ) | ( n3513 & n3567 ) | ( n3556 & n3567 ) ;
  assign n3570 = ( n3556 & n3568 ) | ( n3556 & ~n3569 ) | ( n3568 & ~n3569 ) ;
  assign n3571 = n3519 & ~n3570 ;
  assign n3572 = n2842 & n3515 ;
  assign n3573 = ( n3519 & n3570 ) | ( n3519 & n3572 ) | ( n3570 & n3572 ) ;
  assign n3574 = n3570 | n3572 ;
  assign n3575 = ( n3571 & ~n3573 ) | ( n3571 & n3574 ) | ( ~n3573 & n3574 ) ;
  assign n3576 = n2842 | n3519 ;
  assign n3577 = n3485 & ~n3530 ;
  assign n3578 = n3520 | n3577 ;
  assign n3579 = n3534 | n3578 ;
  assign n3580 = n902 | n3537 ;
  assign n3581 = ( n3538 & n3579 ) | ( n3538 & ~n3580 ) | ( n3579 & ~n3580 ) ;
  assign n3582 = ~n553 & n2023 ;
  assign n3583 = n2011 | n3582 ;
  assign n3584 = ( n2945 & n3582 ) | ( n2945 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3585 = n2026 & ~n2857 ;
  assign n3586 = ( ~n646 & n3584 ) | ( ~n646 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = n646 & ~n3584 ;
  assign n3588 = ( n646 & n3584 ) | ( n646 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3589 = ( n3586 & n3587 ) | ( n3586 & ~n3588 ) | ( n3587 & ~n3588 ) ;
  assign n3590 = n2238 & n2667 ;
  assign n3591 = n2282 & ~n2365 ;
  assign n3592 = n2241 & n2661 ;
  assign n3593 = n3591 | n3592 ;
  assign n3594 = n2236 & n2635 ;
  assign n3595 = n3593 | n3594 ;
  assign n3596 = n3590 | n3595 ;
  assign n3597 = ( ~n902 & n1921 ) | ( ~n902 & n2369 ) | ( n1921 & n2369 ) ;
  assign n3598 = n2367 | n3597 ;
  assign n3599 = n2367 & n3597 ;
  assign n3600 = n3598 & ~n3599 ;
  assign n3601 = n584 & ~n3600 ;
  assign n3602 = ~n3596 & n3601 ;
  assign n3603 = n3596 & ~n3601 ;
  assign n3604 = n3602 | n3603 ;
  assign n3605 = ( n3581 & n3589 ) | ( n3581 & ~n3604 ) | ( n3589 & ~n3604 ) ;
  assign n3606 = ( n3581 & ~n3589 ) | ( n3581 & n3604 ) | ( ~n3589 & n3604 ) ;
  assign n3607 = ( ~n3581 & n3605 ) | ( ~n3581 & n3606 ) | ( n3605 & n3606 ) ;
  assign n3608 = ( n3551 & ~n3554 ) | ( n3551 & n3607 ) | ( ~n3554 & n3607 ) ;
  assign n3609 = ( n3551 & n3554 ) | ( n3551 & n3607 ) | ( n3554 & n3607 ) ;
  assign n3610 = ( n3554 & n3608 ) | ( n3554 & ~n3609 ) | ( n3608 & ~n3609 ) ;
  assign n3611 = n507 | n574 ;
  assign n3612 = n520 | n3611 ;
  assign n3613 = n468 | n3612 ;
  assign n3614 = n537 | n3613 ;
  assign n3615 = n396 | n3614 ;
  assign n3616 = ( n3569 & ~n3610 ) | ( n3569 & n3615 ) | ( ~n3610 & n3615 ) ;
  assign n3617 = ( n3569 & n3610 ) | ( n3569 & n3615 ) | ( n3610 & n3615 ) ;
  assign n3618 = ( n3610 & n3616 ) | ( n3610 & ~n3617 ) | ( n3616 & ~n3617 ) ;
  assign n3619 = ~n3576 & n3618 ;
  assign n3620 = ( n3574 & n3576 ) | ( n3574 & n3618 ) | ( n3576 & n3618 ) ;
  assign n3621 = n3574 & n3618 ;
  assign n3622 = ( n3619 & n3620 ) | ( n3619 & ~n3621 ) | ( n3620 & ~n3621 ) ;
  assign n3623 = ( n2011 & ~n2857 ) | ( n2011 & n2858 ) | ( ~n2857 & n2858 ) ;
  assign n3624 = ( n2023 & ~n3077 ) | ( n2023 & n3623 ) | ( ~n3077 & n3623 ) ;
  assign n3625 = n646 & ~n3624 ;
  assign n3626 = ~n646 & n3624 ;
  assign n3627 = n3625 | n3626 ;
  assign n3628 = ( ~n584 & n2365 ) | ( ~n584 & n3599 ) | ( n2365 & n3599 ) ;
  assign n3629 = n2365 | n3599 ;
  assign n3630 = ( n3596 & ~n3628 ) | ( n3596 & n3629 ) | ( ~n3628 & n3629 ) ;
  assign n3631 = n584 & n3596 ;
  assign n3632 = ( n2365 & n3598 ) | ( n2365 & ~n3631 ) | ( n3598 & ~n3631 ) ;
  assign n3633 = n2365 | n3598 ;
  assign n3634 = ( n3630 & n3632 ) | ( n3630 & ~n3633 ) | ( n3632 & ~n3633 ) ;
  assign n3635 = n2236 & n2661 ;
  assign n3636 = ~n553 & n2241 ;
  assign n3637 = n3635 | n3636 ;
  assign n3638 = n2282 & n2635 ;
  assign n3639 = n3637 | n3638 ;
  assign n3640 = n2238 | n3639 ;
  assign n3641 = ( ~n2768 & n3639 ) | ( ~n2768 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3642 = n584 | n3641 ;
  assign n3643 = n584 & n3641 ;
  assign n3644 = n3642 & ~n3643 ;
  assign n3645 = ( n3627 & n3634 ) | ( n3627 & ~n3644 ) | ( n3634 & ~n3644 ) ;
  assign n3646 = ( n3627 & ~n3634 ) | ( n3627 & n3644 ) | ( ~n3634 & n3644 ) ;
  assign n3647 = ( ~n3627 & n3645 ) | ( ~n3627 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = ( ~n3605 & n3608 ) | ( ~n3605 & n3647 ) | ( n3608 & n3647 ) ;
  assign n3649 = ( n3605 & n3608 ) | ( n3605 & ~n3647 ) | ( n3608 & ~n3647 ) ;
  assign n3650 = ( ~n3608 & n3648 ) | ( ~n3608 & n3649 ) | ( n3648 & n3649 ) ;
  assign n3651 = n1723 | n3011 ;
  assign n3652 = n195 | n247 ;
  assign n3653 = n854 | n3652 ;
  assign n3654 = n130 | n203 ;
  assign n3655 = n112 | n3654 ;
  assign n3656 = n257 | n322 ;
  assign n3657 = n3655 | n3656 ;
  assign n3658 = n3653 | n3657 ;
  assign n3659 = n3651 | n3658 ;
  assign n3660 = n1691 | n3659 ;
  assign n3661 = n1588 | n3660 ;
  assign n3662 = ( ~n3617 & n3650 ) | ( ~n3617 & n3661 ) | ( n3650 & n3661 ) ;
  assign n3663 = ( n3617 & n3650 ) | ( n3617 & n3661 ) | ( n3650 & n3661 ) ;
  assign n3664 = ( n3617 & n3662 ) | ( n3617 & ~n3663 ) | ( n3662 & ~n3663 ) ;
  assign n3665 = n3519 & n3570 ;
  assign n3666 = n3618 & n3665 ;
  assign n3667 = ( n2842 & n3576 ) | ( n2842 & n3666 ) | ( n3576 & n3666 ) ;
  assign n3668 = ( n3572 & n3620 ) | ( n3572 & n3667 ) | ( n3620 & n3667 ) ;
  assign n3669 = n3664 | n3668 ;
  assign n3670 = n3664 & n3668 ;
  assign n3671 = n3669 & ~n3670 ;
  assign n3672 = n240 | n949 ;
  assign n3673 = n1675 | n3168 ;
  assign n3674 = n154 | n711 ;
  assign n3675 = n988 | n3674 ;
  assign n3676 = n3673 | n3675 ;
  assign n3677 = n1649 | n3676 ;
  assign n3678 = n3672 | n3677 ;
  assign n3679 = n2567 | n2928 ;
  assign n3680 = n135 | n3679 ;
  assign n3681 = n3678 | n3680 ;
  assign n3682 = ( n2365 & n3604 ) | ( n2365 & n3634 ) | ( n3604 & n3634 ) ;
  assign n3683 = n2241 & ~n2857 ;
  assign n3684 = ~n553 & n2236 ;
  assign n3685 = n3683 | n3684 ;
  assign n3686 = n2282 & n2661 ;
  assign n3687 = n3685 | n3686 ;
  assign n3688 = ( n2238 & n2861 ) | ( n2238 & n3687 ) | ( n2861 & n3687 ) ;
  assign n3689 = n584 & ~n3687 ;
  assign n3690 = n3688 | n3689 ;
  assign n3691 = ( n3687 & ~n3688 ) | ( n3687 & n3689 ) | ( ~n3688 & n3689 ) ;
  assign n3692 = ( ~n584 & n3690 ) | ( ~n584 & n3691 ) | ( n3690 & n3691 ) ;
  assign n3693 = ( n584 & ~n2365 ) | ( n584 & n2635 ) | ( ~n2365 & n2635 ) ;
  assign n3694 = ~n2365 & n2635 ;
  assign n3695 = ( n646 & ~n3693 ) | ( n646 & n3694 ) | ( ~n3693 & n3694 ) ;
  assign n3696 = ( n646 & n3693 ) | ( n646 & n3694 ) | ( n3693 & n3694 ) ;
  assign n3697 = ( n3693 & n3695 ) | ( n3693 & ~n3696 ) | ( n3695 & ~n3696 ) ;
  assign n3698 = ( n3682 & ~n3692 ) | ( n3682 & n3697 ) | ( ~n3692 & n3697 ) ;
  assign n3699 = ( n3682 & n3692 ) | ( n3682 & ~n3697 ) | ( n3692 & ~n3697 ) ;
  assign n3700 = ( ~n3682 & n3698 ) | ( ~n3682 & n3699 ) | ( n3698 & n3699 ) ;
  assign n3701 = ( ~n3646 & n3648 ) | ( ~n3646 & n3700 ) | ( n3648 & n3700 ) ;
  assign n3702 = ( n3646 & n3648 ) | ( n3646 & ~n3700 ) | ( n3648 & ~n3700 ) ;
  assign n3703 = ( ~n3648 & n3701 ) | ( ~n3648 & n3702 ) | ( n3701 & n3702 ) ;
  assign n3704 = ( n3663 & n3681 ) | ( n3663 & n3703 ) | ( n3681 & n3703 ) ;
  assign n3705 = ( ~n3663 & n3681 ) | ( ~n3663 & n3703 ) | ( n3681 & n3703 ) ;
  assign n3706 = ( n3663 & ~n3704 ) | ( n3663 & n3705 ) | ( ~n3704 & n3705 ) ;
  assign n3707 = ( n2842 & n3664 ) | ( n2842 & n3668 ) | ( n3664 & n3668 ) ;
  assign n3708 = n3706 & ~n3707 ;
  assign n3709 = ~n3706 & n3707 ;
  assign n3710 = n3708 | n3709 ;
  assign n3711 = n2236 & ~n2857 ;
  assign n3712 = ~n553 & n2282 ;
  assign n3713 = n3711 | n3712 ;
  assign n3714 = n2238 | n3713 ;
  assign n3715 = ( n2945 & n3713 ) | ( n2945 & n3714 ) | ( n3713 & n3714 ) ;
  assign n3716 = ( n646 & n2365 ) | ( n646 & ~n2635 ) | ( n2365 & ~n2635 ) ;
  assign n3717 = n584 & ~n3716 ;
  assign n3718 = n584 & ~n2661 ;
  assign n3719 = ( n3715 & n3717 ) | ( n3715 & n3718 ) | ( n3717 & n3718 ) ;
  assign n3720 = ( ~n3715 & n3717 ) | ( ~n3715 & n3718 ) | ( n3717 & n3718 ) ;
  assign n3721 = ( n3715 & ~n3719 ) | ( n3715 & n3720 ) | ( ~n3719 & n3720 ) ;
  assign n3722 = ( n3699 & n3701 ) | ( n3699 & ~n3721 ) | ( n3701 & ~n3721 ) ;
  assign n3723 = ( ~n3699 & n3701 ) | ( ~n3699 & n3721 ) | ( n3701 & n3721 ) ;
  assign n3724 = ( ~n3701 & n3722 ) | ( ~n3701 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = n165 | n397 ;
  assign n3726 = n323 | n3725 ;
  assign n3727 = n209 | n269 ;
  assign n3728 = n3726 | n3727 ;
  assign n3729 = n1723 | n3728 ;
  assign n3730 = n879 | n3729 ;
  assign n3731 = n1194 | n3730 ;
  assign n3732 = n368 | n428 ;
  assign n3733 = n177 | n3324 ;
  assign n3734 = n3732 | n3733 ;
  assign n3735 = n453 | n3734 ;
  assign n3736 = n1621 | n3735 ;
  assign n3737 = n3731 | n3736 ;
  assign n3738 = ( ~n3704 & n3724 ) | ( ~n3704 & n3737 ) | ( n3724 & n3737 ) ;
  assign n3739 = ( n3704 & n3724 ) | ( n3704 & n3737 ) | ( n3724 & n3737 ) ;
  assign n3740 = ( n3704 & n3738 ) | ( n3704 & ~n3739 ) | ( n3738 & ~n3739 ) ;
  assign n3741 = n3664 & n3666 ;
  assign n3742 = n3706 & n3741 ;
  assign n3743 = n2842 | n3742 ;
  assign n3744 = n3740 & ~n3743 ;
  assign n3745 = n3669 | n3706 ;
  assign n3746 = ( n3740 & n3743 ) | ( n3740 & n3745 ) | ( n3743 & n3745 ) ;
  assign n3747 = n3740 & n3745 ;
  assign n3748 = ( n3744 & n3746 ) | ( n3744 & ~n3747 ) | ( n3746 & ~n3747 ) ;
  assign n3749 = ( n553 & ~n584 ) | ( n553 & n2661 ) | ( ~n584 & n2661 ) ;
  assign n3750 = n553 | n2661 ;
  assign n3751 = ( n2238 & ~n2857 ) | ( n2238 & n2858 ) | ( ~n2857 & n2858 ) ;
  assign n3752 = ( n2282 & ~n3077 ) | ( n2282 & n3751 ) | ( ~n3077 & n3751 ) ;
  assign n3753 = ( n3749 & ~n3750 ) | ( n3749 & n3752 ) | ( ~n3750 & n3752 ) ;
  assign n3754 = ( n3749 & n3750 ) | ( n3749 & ~n3752 ) | ( n3750 & ~n3752 ) ;
  assign n3755 = ( ~n3749 & n3753 ) | ( ~n3749 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3756 = n584 | n3721 ;
  assign n3757 = ( ~n584 & n3720 ) | ( ~n584 & n3756 ) | ( n3720 & n3756 ) ;
  assign n3758 = ( n3723 & n3755 ) | ( n3723 & ~n3757 ) | ( n3755 & ~n3757 ) ;
  assign n3759 = ( n3723 & ~n3755 ) | ( n3723 & n3757 ) | ( ~n3755 & n3757 ) ;
  assign n3760 = ( ~n3723 & n3758 ) | ( ~n3723 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3761 = n421 | n1785 ;
  assign n3762 = n999 | n3761 ;
  assign n3763 = n96 | n889 ;
  assign n3764 = n1640 | n3732 ;
  assign n3765 = n3763 | n3764 ;
  assign n3766 = n1854 | n3657 ;
  assign n3767 = n3765 | n3766 ;
  assign n3768 = n940 | n3767 ;
  assign n3769 = n1732 | n3768 ;
  assign n3770 = n3762 | n3769 ;
  assign n3771 = ( ~n3739 & n3760 ) | ( ~n3739 & n3770 ) | ( n3760 & n3770 ) ;
  assign n3772 = ( n3739 & n3760 ) | ( n3739 & n3770 ) | ( n3760 & n3770 ) ;
  assign n3773 = ( n3739 & n3771 ) | ( n3739 & ~n3772 ) | ( n3771 & ~n3772 ) ;
  assign n3774 = ( n2842 & n3707 ) | ( n2842 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3775 = ( n3740 & n3743 ) | ( n3740 & n3774 ) | ( n3743 & n3774 ) ;
  assign n3776 = n3773 & n3775 ;
  assign n3777 = n3773 | n3775 ;
  assign n3778 = ~n3776 & n3777 ;
  assign n3779 = n584 & n2234 ;
  assign n3780 = ~n2857 & n3779 ;
  assign n3781 = ~n3758 & n3780 ;
  assign n3782 = n102 | n1196 ;
  assign n3783 = n668 | n3782 ;
  assign n3784 = n876 | n1694 ;
  assign n3785 = n3783 | n3784 ;
  assign n3786 = n2741 | n3785 ;
  assign n3787 = n416 | n3673 ;
  assign n3788 = n218 | n3787 ;
  assign n3789 = n3786 | n3788 ;
  assign n3790 = n1868 | n3789 ;
  assign n3791 = ( n3772 & n3781 ) | ( n3772 & ~n3790 ) | ( n3781 & ~n3790 ) ;
  assign n3792 = ( n3772 & ~n3781 ) | ( n3772 & n3790 ) | ( ~n3781 & n3790 ) ;
  assign n3793 = ( ~n3772 & n3791 ) | ( ~n3772 & n3792 ) | ( n3791 & n3792 ) ;
  assign n3794 = ( n2842 & n3773 ) | ( n2842 & n3775 ) | ( n3773 & n3775 ) ;
  assign n3795 = ~n3793 & n3794 ;
  assign n3796 = n3793 & ~n3794 ;
  assign n3797 = n3795 | n3796 ;
  assign n3798 = n3740 & n3742 ;
  assign n3799 = n3773 & n3798 ;
  assign n3800 = n3793 & ~n3799 ;
  assign n3801 = ( n3781 & n3790 ) | ( n3781 & ~n3800 ) | ( n3790 & ~n3800 ) ;
  assign n3802 = n750 | n830 ;
  assign n3803 = n695 | n3802 ;
  assign n3804 = n137 | n371 ;
  assign n3805 = n112 | n3804 ;
  assign n3806 = n450 | n1594 ;
  assign n3807 = n3805 | n3806 ;
  assign n3808 = n244 | n3807 ;
  assign n3809 = n3803 | n3808 ;
  assign n3810 = n342 | n3809 ;
  assign n3811 = n2351 | n3810 ;
  assign n3812 = n3801 & n3811 ;
  assign n3813 = n3801 | n3811 ;
  assign n3814 = ~n3812 & n3813 ;
  assign n3815 = ( n2842 & n3795 ) | ( n2842 & n3800 ) | ( n3795 & n3800 ) ;
  assign n3816 = n3814 | n3815 ;
  assign n3817 = n3814 & n3815 ;
  assign n3818 = n3816 & ~n3817 ;
  assign n3819 = n2842 & n3816 ;
  assign n3820 = n528 | n1010 ;
  assign n3821 = n1647 | n3820 ;
  assign n3822 = n513 | n3821 ;
  assign n3823 = n256 | n3822 ;
  assign n3824 = n261 | n390 ;
  assign n3825 = n2327 | n3824 ;
  assign n3826 = n456 | n3825 ;
  assign n3827 = n953 | n3826 ;
  assign n3828 = n2552 | n3827 ;
  assign n3829 = n3823 | n3828 ;
  assign n3830 = n3812 & n3829 ;
  assign n3831 = n3812 | n3829 ;
  assign n3832 = ~n3830 & n3831 ;
  assign n3833 = n3819 | n3832 ;
  assign n3834 = n3819 & n3832 ;
  assign n3835 = n3833 & ~n3834 ;
  assign n3836 = n2842 & n3833 ;
  assign n3837 = n136 | n385 ;
  assign n3838 = n259 | n3837 ;
  assign n3839 = n3243 | n3838 ;
  assign n3840 = n108 | n241 ;
  assign n3841 = n1169 | n3840 ;
  assign n3842 = n373 | n3841 ;
  assign n3843 = n3839 | n3842 ;
  assign n3844 = n2322 | n3843 ;
  assign n3845 = n851 | n3844 ;
  assign n3846 = n3762 | n3845 ;
  assign n3847 = n3830 & n3846 ;
  assign n3848 = n3830 | n3846 ;
  assign n3849 = ~n3847 & n3848 ;
  assign n3850 = n3836 | n3849 ;
  assign n3851 = n3836 & n3849 ;
  assign n3852 = n3850 & ~n3851 ;
  assign n3853 = n503 & n3847 ;
  assign n3854 = n2842 & ~n3853 ;
  assign n3855 = n3850 & n3854 ;
  assign n3856 = n503 | n3847 ;
  assign n3857 = ~n3836 & n3853 ;
  assign n3858 = ( n3855 & n3856 ) | ( n3855 & ~n3857 ) | ( n3856 & ~n3857 ) ;
  assign n3859 = n3855 & n3856 ;
  assign n3860 = n3858 & ~n3859 ;
  assign n3861 = n154 | n593 ;
  assign n3862 = n640 | n3861 ;
  assign n3863 = n559 | n3862 ;
  assign n3864 = n3857 & ~n3863 ;
  assign n3865 = n3854 & n3863 ;
  assign n3866 = ( n3855 & ~n3857 ) | ( n3855 & n3863 ) | ( ~n3857 & n3863 ) ;
  assign n3867 = ( n3864 & ~n3865 ) | ( n3864 & n3866 ) | ( ~n3865 & n3866 ) ;
  assign n3868 = n3853 & n3863 ;
  assign n3869 = n664 & ~n3868 ;
  assign n3870 = ( n600 & ~n664 ) | ( n600 & n3868 ) | ( ~n664 & n3868 ) ;
  assign n3871 = ( n34 & n2842 ) | ( n34 & n3836 ) | ( n2842 & n3836 ) ;
  assign n3872 = ( n3869 & ~n3870 ) | ( n3869 & n3871 ) | ( ~n3870 & n3871 ) ;
  assign n3873 = ( n3869 & n3870 ) | ( n3869 & ~n3871 ) | ( n3870 & ~n3871 ) ;
  assign n3874 = ( ~n664 & n3872 ) | ( ~n664 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = n55 & ~n3871 ;
  assign n3876 = ( ~n3871 & n3874 ) | ( ~n3871 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3877 = n2840 | n3871 ;
  assign y0 = n2839 ;
  assign y1 = n2943 ;
  assign y2 = n3027 ;
  assign y3 = n3110 ;
  assign y4 = n3182 ;
  assign y5 = n3259 ;
  assign y6 = n3337 ;
  assign y7 = n3403 ;
  assign y8 = n3461 ;
  assign y9 = n3517 ;
  assign y10 = n3575 ;
  assign y11 = n3622 ;
  assign y12 = n3671 ;
  assign y13 = n3710 ;
  assign y14 = n3748 ;
  assign y15 = n3778 ;
  assign y16 = n3797 ;
  assign y17 = n3818 ;
  assign y18 = n3835 ;
  assign y19 = n3852 ;
  assign y20 = n3860 ;
  assign y21 = n3867 ;
  assign y22 = n3874 ;
  assign y23 = ~n3876 ;
  assign y24 = n3877 ;
endmodule
