module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 ;
  assign n1205 = x105 & x228 ;
  assign n1206 = x39 | x87 ;
  assign n1207 = x56 | x62 ;
  assign n1208 = n1206 | n1207 ;
  assign n1209 = x100 | n1208 ;
  assign n1210 = x63 | x64 ;
  assign n1211 = x107 | n1210 ;
  assign n1212 = x36 | n1211 ;
  assign n1213 = x69 | x83 ;
  assign n1214 = x82 | x103 ;
  assign n1215 = n1213 | n1214 ;
  assign n1216 = ( ~x67 & n1212 ) | ( ~x67 & n1215 ) | ( n1212 & n1215 ) ;
  assign n1217 = x48 & x49 ;
  assign n1218 = x68 | x71 ;
  assign n1219 = ~x73 & x85 ;
  assign n1220 = x84 | n1219 ;
  assign n1221 = ( x73 & n1218 ) | ( x73 & n1220 ) | ( n1218 & n1220 ) ;
  assign n1222 = n1217 | n1221 ;
  assign n1223 = ( ~x67 & n1216 ) | ( ~x67 & n1222 ) | ( n1216 & n1222 ) ;
  assign n1224 = x67 | n1223 ;
  assign n1225 = x66 | x76 ;
  assign n1226 = x61 | n1225 ;
  assign n1227 = x48 | x49 ;
  assign n1228 = x104 | x106 ;
  assign n1229 = x89 | n1228 ;
  assign n1230 = ( ~n1226 & n1227 ) | ( ~n1226 & n1229 ) | ( n1227 & n1229 ) ;
  assign n1231 = n1226 | n1230 ;
  assign n1232 = n1224 | n1231 ;
  assign n1233 = x73 | x84 ;
  assign n1234 = ( x85 & n1218 ) | ( x85 & ~n1233 ) | ( n1218 & ~n1233 ) ;
  assign n1235 = n1233 | n1234 ;
  assign n1236 = x45 | x111 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = n1232 | n1237 ;
  assign n1239 = x53 | x60 ;
  assign n1240 = x50 | n1239 ;
  assign n1241 = x88 | x98 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = x77 | x86 ;
  assign n1244 = x81 | n1243 ;
  assign n1245 = n1242 | n1244 ;
  assign n1246 = n1238 | n1245 ;
  assign n1247 = x97 | x108 ;
  assign n1248 = x110 | n1247 ;
  assign n1249 = x47 | x58 ;
  assign n1250 = x109 | n1249 ;
  assign n1251 = n1248 | n1250 ;
  assign n1252 = x46 | x91 ;
  assign n1253 = n1251 | n1252 ;
  assign n1254 = x65 | x102 ;
  assign n1255 = x94 | n1254 ;
  assign n1256 = n1253 | n1255 ;
  assign n1257 = n1246 | n1256 ;
  assign n1258 = x90 | x93 ;
  assign n1259 = ( x35 & x90 ) | ( x35 & n1258 ) | ( x90 & n1258 ) ;
  assign n1260 = x35 | x93 ;
  assign n1261 = x90 | n1260 ;
  assign n1262 = x51 | x70 ;
  assign n1263 = n1261 | n1262 ;
  assign n1264 = x72 | n1263 ;
  assign n1265 = ( x32 & x95 ) | ( x32 & ~x96 ) | ( x95 & ~x96 ) ;
  assign n1266 = ( x32 & x40 ) | ( x32 & x95 ) | ( x40 & x95 ) ;
  assign n1267 = ( x32 & x40 ) | ( x32 & x96 ) | ( x40 & x96 ) ;
  assign n1268 = ( x40 & ~x95 ) | ( x40 & x96 ) | ( ~x95 & x96 ) ;
  assign n1269 = ~n1267 & n1268 ;
  assign n1270 = ( n1265 & ~n1266 ) | ( n1265 & n1269 ) | ( ~n1266 & n1269 ) ;
  assign n1271 = n1264 & n1270 ;
  assign n1272 = x40 | x96 ;
  assign n1273 = x32 | n1272 ;
  assign n1274 = x51 & x70 ;
  assign n1275 = x72 | n1274 ;
  assign n1276 = ( n1261 & n1262 ) | ( n1261 & n1275 ) | ( n1262 & n1275 ) ;
  assign n1277 = n1273 | n1276 ;
  assign n1278 = n1264 & ~n1277 ;
  assign n1279 = ~n1264 & n1270 ;
  assign n1280 = ( ~n1271 & n1278 ) | ( ~n1271 & n1279 ) | ( n1278 & n1279 ) ;
  assign n1281 = ~n1259 & n1280 ;
  assign n1282 = ~n1257 & n1281 ;
  assign n1283 = x95 | n1253 ;
  assign n1284 = n1264 | n1283 ;
  assign n1285 = n1277 | n1284 ;
  assign n1286 = n1255 | n1277 ;
  assign n1287 = x47 | n1247 ;
  assign n1288 = x58 | x110 ;
  assign n1289 = n1287 & n1288 ;
  assign n1290 = n1264 | n1289 ;
  assign n1291 = ( x46 & x91 ) | ( x46 & n1251 ) | ( x91 & n1251 ) ;
  assign n1292 = ( n1253 & n1290 ) | ( n1253 & n1291 ) | ( n1290 & n1291 ) ;
  assign n1293 = ( x109 & n1248 ) | ( x109 & n1249 ) | ( n1248 & n1249 ) ;
  assign n1294 = x95 | n1260 ;
  assign n1295 = x97 & x108 ;
  assign n1296 = ( ~n1293 & n1294 ) | ( ~n1293 & n1295 ) | ( n1294 & n1295 ) ;
  assign n1297 = n1293 | n1296 ;
  assign n1298 = ( ~n1286 & n1292 ) | ( ~n1286 & n1297 ) | ( n1292 & n1297 ) ;
  assign n1299 = n1286 | n1298 ;
  assign n1300 = n1285 & n1299 ;
  assign n1301 = ( n1246 & n1285 ) | ( n1246 & n1300 ) | ( n1285 & n1300 ) ;
  assign n1302 = ( x50 & x53 ) | ( x50 & x60 ) | ( x53 & x60 ) ;
  assign n1303 = ( x50 & ~x53 ) | ( x50 & x60 ) | ( ~x53 & x60 ) ;
  assign n1304 = n1238 | n1255 ;
  assign n1305 = n1244 | n1304 ;
  assign n1306 = n1241 | n1305 ;
  assign n1307 = ( x53 & n1303 ) | ( x53 & ~n1306 ) | ( n1303 & ~n1306 ) ;
  assign n1308 = ~n1302 & n1307 ;
  assign n1309 = x90 | x91 ;
  assign n1310 = n1242 | n1304 ;
  assign n1311 = ( x77 & x86 ) | ( x77 & ~n1310 ) | ( x86 & ~n1310 ) ;
  assign n1312 = ( x77 & x81 ) | ( x77 & x86 ) | ( x81 & x86 ) ;
  assign n1313 = n1311 & ~n1312 ;
  assign n1314 = n1309 | n1313 ;
  assign n1315 = n1308 | n1314 ;
  assign n1316 = ( x88 & x98 ) | ( x88 & ~n1240 ) | ( x98 & ~n1240 ) ;
  assign n1317 = ( x88 & x98 ) | ( x88 & n1305 ) | ( x98 & n1305 ) ;
  assign n1318 = n1316 & ~n1317 ;
  assign n1319 = n1251 | n1318 ;
  assign n1320 = ( x65 & x94 ) | ( x65 & x102 ) | ( x94 & x102 ) ;
  assign n1321 = ( x65 & ~x94 ) | ( x65 & x102 ) | ( ~x94 & x102 ) ;
  assign n1322 = ( x94 & ~n1246 ) | ( x94 & n1321 ) | ( ~n1246 & n1321 ) ;
  assign n1323 = ~n1320 & n1322 ;
  assign n1324 = n1319 | n1323 ;
  assign n1325 = n1315 | n1324 ;
  assign n1326 = x81 & ~n1243 ;
  assign n1327 = ~n1310 & n1326 ;
  assign n1328 = x82 & x83 ;
  assign n1329 = n1236 | n1328 ;
  assign n1330 = n1235 & ~n1329 ;
  assign n1331 = x36 & n1211 ;
  assign n1332 = n1245 | n1331 ;
  assign n1333 = ( x67 & n1212 ) | ( x67 & n1215 ) | ( n1212 & n1215 ) ;
  assign n1334 = x69 & x103 ;
  assign n1335 = x68 & x71 ;
  assign n1336 = x63 & x64 ;
  assign n1337 = ( ~n1334 & n1335 ) | ( ~n1334 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1338 = n1334 | n1337 ;
  assign n1339 = n1255 | n1338 ;
  assign n1340 = ( n1226 & n1227 ) | ( n1226 & n1229 ) | ( n1227 & n1229 ) ;
  assign n1341 = ( ~n1333 & n1339 ) | ( ~n1333 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1342 = n1333 | n1341 ;
  assign n1343 = x82 | x83 ;
  assign n1344 = x69 | x103 ;
  assign n1345 = n1343 & n1344 ;
  assign n1346 = x107 & n1210 ;
  assign n1347 = n1345 | n1346 ;
  assign n1348 = ( x89 & x104 ) | ( x89 & x106 ) | ( x104 & x106 ) ;
  assign n1349 = x85 & n1233 ;
  assign n1350 = ( ~n1347 & n1348 ) | ( ~n1347 & n1349 ) | ( n1348 & n1349 ) ;
  assign n1351 = n1347 | n1350 ;
  assign n1352 = ( x61 & x66 ) | ( x61 & x76 ) | ( x66 & x76 ) ;
  assign n1353 = ( ~n1339 & n1351 ) | ( ~n1339 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1354 = ( ~n1332 & n1342 ) | ( ~n1332 & n1353 ) | ( n1342 & n1353 ) ;
  assign n1355 = n1332 | n1354 ;
  assign n1356 = n1235 | n1329 ;
  assign n1357 = n1232 & n1356 ;
  assign n1358 = n1355 | n1357 ;
  assign n1359 = n1224 & n1231 ;
  assign n1360 = n1232 & ~n1359 ;
  assign n1361 = ( ~n1235 & n1329 ) | ( ~n1235 & n1360 ) | ( n1329 & n1360 ) ;
  assign n1362 = ( n1330 & ~n1358 ) | ( n1330 & n1361 ) | ( ~n1358 & n1361 ) ;
  assign n1363 = x45 & x111 ;
  assign n1364 = n1362 & ~n1363 ;
  assign n1365 = n1327 | n1364 ;
  assign n1366 = ~n1301 & n1365 ;
  assign n1367 = ( ~n1301 & n1325 ) | ( ~n1301 & n1366 ) | ( n1325 & n1366 ) ;
  assign n1368 = n1282 | n1367 ;
  assign n1369 = x55 | x92 ;
  assign n1370 = ( ~n1209 & n1368 ) | ( ~n1209 & n1369 ) | ( n1368 & n1369 ) ;
  assign n1371 = n1209 | n1370 ;
  assign n1372 = x74 | x92 ;
  assign n1373 = x75 | x100 ;
  assign n1374 = x38 | x54 ;
  assign n1375 = x57 | x59 ;
  assign n1376 = n1374 | n1375 ;
  assign n1377 = n1373 | n1376 ;
  assign n1378 = x55 | x57 ;
  assign n1379 = n1207 | n1378 ;
  assign n1380 = x59 | n1379 ;
  assign n1381 = ( ~n1372 & n1377 ) | ( ~n1372 & n1380 ) | ( n1377 & n1380 ) ;
  assign n1382 = n1372 | n1381 ;
  assign n1383 = n1206 | n1382 ;
  assign n1384 = x38 | x100 ;
  assign n1385 = n1206 | n1384 ;
  assign n1386 = x75 | n1385 ;
  assign n1387 = x95 | n1273 ;
  assign n1388 = ( n1257 & n1263 ) | ( n1257 & ~n1387 ) | ( n1263 & ~n1387 ) ;
  assign n1389 = n1387 | n1388 ;
  assign n1390 = x72 | n1389 ;
  assign n1391 = n1372 | n1390 ;
  assign n1392 = x54 | n1391 ;
  assign n1393 = n1386 | n1392 ;
  assign n1394 = x59 | n1393 ;
  assign n1395 = x55 | n1394 ;
  assign n1396 = n1380 | n1392 ;
  assign n1397 = x75 | n1206 ;
  assign n1398 = x38 | x39 ;
  assign n1399 = ( x38 & x87 ) | ( x38 & n1398 ) | ( x87 & n1398 ) ;
  assign n1400 = ( n1373 & n1397 ) | ( n1373 & n1399 ) | ( n1397 & n1399 ) ;
  assign n1401 = n1396 | n1400 ;
  assign n1402 = x62 | n1401 ;
  assign n1403 = ( x62 & n1395 ) | ( x62 & n1402 ) | ( n1395 & n1402 ) ;
  assign n1404 = n1378 | n1394 ;
  assign n1405 = ( x56 & n1403 ) | ( x56 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1406 = n1380 | n1386 ;
  assign n1407 = n1390 | n1406 ;
  assign n1408 = ( x54 & x74 ) | ( x54 & x92 ) | ( x74 & x92 ) ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = ( n1385 & n1396 ) | ( n1385 & n1401 ) | ( n1396 & n1401 ) ;
  assign n1411 = n1409 & n1410 ;
  assign n1412 = ( x55 & n1208 ) | ( x55 & n1377 ) | ( n1208 & n1377 ) ;
  assign n1413 = ( x55 & n1391 ) | ( x55 & n1412 ) | ( n1391 & n1412 ) ;
  assign n1414 = x55 & ~n1413 ;
  assign n1415 = n1411 & ~n1414 ;
  assign n1416 = n1405 & n1415 ;
  assign n1417 = n1383 & n1416 ;
  assign n1418 = n1371 & ~n1417 ;
  assign n1419 = x228 & ~n1205 ;
  assign n1420 = ( n1205 & n1418 ) | ( n1205 & ~n1419 ) | ( n1418 & ~n1419 ) ;
  assign n1421 = x299 | n1380 ;
  assign n1422 = ~x215 & n1421 ;
  assign n1423 = ~x221 & n1422 ;
  assign n1424 = ~x216 & n1423 ;
  assign n1425 = n1420 & n1424 ;
  assign n1426 = x223 | x299 ;
  assign n1427 = ( x222 & n1380 ) | ( x222 & ~n1426 ) | ( n1380 & ~n1426 ) ;
  assign n1428 = n1426 | n1427 ;
  assign n1429 = x224 & ~n1428 ;
  assign n1430 = ( ~n1425 & n1428 ) | ( ~n1425 & n1429 ) | ( n1428 & n1429 ) ;
  assign n1431 = x95 & ~x479 ;
  assign n1432 = x96 & ~n1383 ;
  assign n1433 = n1282 & n1432 ;
  assign n1434 = n1431 | n1433 ;
  assign n1435 = ~x161 & x299 ;
  assign n1436 = x152 | x166 ;
  assign n1437 = n1435 & ~n1436 ;
  assign n1438 = x146 & x299 ;
  assign n1439 = n1437 | n1438 ;
  assign n1440 = ~x228 & x252 ;
  assign n1441 = x100 & n1440 ;
  assign n1442 = n1439 & n1441 ;
  assign n1443 = n1434 | n1442 ;
  assign n1444 = n1430 | n1443 ;
  assign n1445 = x198 & ~x299 ;
  assign n1446 = x210 & x299 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = x32 & ~x841 ;
  assign n1449 = ~n1447 & n1448 ;
  assign n1450 = x70 | n1449 ;
  assign n1451 = x32 | x35 ;
  assign n1452 = ~x225 & n1451 ;
  assign n1453 = n1450 | n1452 ;
  assign n1454 = x142 & ~x299 ;
  assign n1455 = n1438 | n1454 ;
  assign n1456 = x174 & ~x299 ;
  assign n1457 = x144 | x299 ;
  assign n1458 = x189 & ~x299 ;
  assign n1459 = ( ~n1437 & n1457 ) | ( ~n1437 & n1458 ) | ( n1457 & n1458 ) ;
  assign n1460 = n1456 | n1459 ;
  assign n1461 = ~n1455 & n1460 ;
  assign n1462 = n1447 | n1461 ;
  assign n1463 = ~x1091 & x1093 ;
  assign n1464 = x829 & x1092 ;
  assign n1465 = ~n1463 & n1464 ;
  assign n1466 = ~x833 & x957 ;
  assign n1467 = x1091 & n1466 ;
  assign n1468 = x950 & ~x1093 ;
  assign n1469 = ( x950 & ~n1467 ) | ( x950 & n1468 ) | ( ~n1467 & n1468 ) ;
  assign n1470 = n1465 & n1469 ;
  assign n1471 = x97 & x1093 ;
  assign n1472 = x96 & ~x841 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1470 & n1473 ;
  assign n1475 = ~n1462 & n1474 ;
  assign n1476 = x137 | n1239 ;
  assign n1477 = n1451 | n1476 ;
  assign n1478 = ~n1453 & n1477 ;
  assign n1479 = ( ~n1453 & n1475 ) | ( ~n1453 & n1478 ) | ( n1475 & n1478 ) ;
  assign n1480 = x70 & x332 ;
  assign n1481 = n1479 | n1480 ;
  assign n1482 = n1301 | n1383 ;
  assign n1483 = x46 & ~n1482 ;
  assign n1484 = ( n1315 & ~n1482 ) | ( n1315 & n1483 ) | ( ~n1482 & n1483 ) ;
  assign n1485 = n1368 & ~n1383 ;
  assign n1486 = ~n1484 & n1485 ;
  assign n1487 = ( n1481 & n1484 ) | ( n1481 & n1486 ) | ( n1484 & n1486 ) ;
  assign n1488 = n1379 | n1393 ;
  assign n1489 = n1416 | n1488 ;
  assign n1490 = n1416 & n1488 ;
  assign n1491 = n1489 & ~n1490 ;
  assign n1492 = x137 | n1373 ;
  assign n1493 = ( x137 & ~n1462 ) | ( x137 & n1492 ) | ( ~n1462 & n1492 ) ;
  assign n1494 = ( n1414 & n1487 ) | ( n1414 & ~n1493 ) | ( n1487 & ~n1493 ) ;
  assign n1495 = n1493 | n1494 ;
  assign n1496 = ( n1487 & n1491 ) | ( n1487 & n1495 ) | ( n1491 & n1495 ) ;
  assign n1497 = n1444 | n1496 ;
  assign n1498 = ~x216 & n1422 ;
  assign n1499 = x223 | x224 ;
  assign n1500 = x833 & ~n1421 ;
  assign n1501 = ~n1499 & n1500 ;
  assign n1502 = ( x833 & n1498 ) | ( x833 & n1501 ) | ( n1498 & n1501 ) ;
  assign n1503 = ~x929 & n1502 ;
  assign n1504 = x265 & ~n1428 ;
  assign n1505 = ~x1144 & n1428 ;
  assign n1506 = ( ~n1502 & n1504 ) | ( ~n1502 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1507 = ( ~n1423 & n1503 ) | ( ~n1423 & n1506 ) | ( n1503 & n1506 ) ;
  assign n1508 = x153 & ~x216 ;
  assign n1509 = x216 & x265 ;
  assign n1510 = ( n1423 & n1508 ) | ( n1423 & n1509 ) | ( n1508 & n1509 ) ;
  assign n1511 = n1507 | n1510 ;
  assign n1512 = ~n1430 & n1434 ;
  assign n1513 = ~x234 & n1512 ;
  assign n1514 = ( ~n1444 & n1511 ) | ( ~n1444 & n1512 ) | ( n1511 & n1512 ) ;
  assign n1515 = ( n1511 & n1513 ) | ( n1511 & ~n1514 ) | ( n1513 & ~n1514 ) ;
  assign n1516 = ( x332 & n1497 ) | ( x332 & ~n1515 ) | ( n1497 & ~n1515 ) ;
  assign n1517 = ~n1423 & n1428 ;
  assign n1518 = n1502 & n1517 ;
  assign n1519 = x939 & n1518 ;
  assign n1520 = ( n1423 & ~n1424 ) | ( n1423 & n1429 ) | ( ~n1424 & n1429 ) ;
  assign n1521 = x276 & n1520 ;
  assign n1522 = n1519 | n1521 ;
  assign n1523 = ~n1502 & n1517 ;
  assign n1524 = x1146 & n1523 ;
  assign n1525 = n1424 & n1442 ;
  assign n1526 = ( ~n1420 & n1424 ) | ( ~n1420 & n1525 ) | ( n1424 & n1525 ) ;
  assign n1527 = x154 & ~n1524 ;
  assign n1528 = ( n1524 & n1526 ) | ( n1524 & ~n1527 ) | ( n1526 & ~n1527 ) ;
  assign n1529 = n1522 | n1528 ;
  assign n1530 = x239 & n1512 ;
  assign n1531 = n1529 | n1530 ;
  assign n1532 = x1145 & n1523 ;
  assign n1533 = ~x274 & n1520 ;
  assign n1534 = x927 & n1518 ;
  assign n1535 = ( ~n1532 & n1533 ) | ( ~n1532 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = n1532 | n1535 ;
  assign n1537 = x151 & ~n1536 ;
  assign n1538 = ( n1526 & n1536 ) | ( n1526 & ~n1537 ) | ( n1536 & ~n1537 ) ;
  assign n1539 = x235 | n1538 ;
  assign n1540 = ( n1512 & n1538 ) | ( n1512 & n1539 ) | ( n1538 & n1539 ) ;
  assign n1541 = x284 & ~n1444 ;
  assign n1542 = ~x238 & n1512 ;
  assign n1543 = ~x944 & n1518 ;
  assign n1544 = x146 & ~n1543 ;
  assign n1545 = ( n1526 & n1543 ) | ( n1526 & ~n1544 ) | ( n1543 & ~n1544 ) ;
  assign n1546 = ~x1143 & n1523 ;
  assign n1547 = x264 & n1520 ;
  assign n1548 = ( ~n1545 & n1546 ) | ( ~n1545 & n1547 ) | ( n1546 & n1547 ) ;
  assign n1549 = n1545 | n1548 ;
  assign n1550 = ( ~n1541 & n1542 ) | ( ~n1541 & n1549 ) | ( n1542 & n1549 ) ;
  assign n1551 = n1541 | n1550 ;
  assign n1552 = ~x277 & n1520 ;
  assign n1553 = x249 | n1552 ;
  assign n1554 = ( n1512 & n1552 ) | ( n1512 & n1553 ) | ( n1552 & n1553 ) ;
  assign n1555 = x932 & n1502 ;
  assign n1556 = x1142 & ~n1502 ;
  assign n1557 = ( n1517 & n1555 ) | ( n1517 & n1556 ) | ( n1555 & n1556 ) ;
  assign n1558 = x172 & ~n1557 ;
  assign n1559 = ( n1526 & n1557 ) | ( n1526 & ~n1558 ) | ( n1557 & ~n1558 ) ;
  assign n1560 = x262 & ~n1559 ;
  assign n1561 = ( n1444 & ~n1559 ) | ( n1444 & n1560 ) | ( ~n1559 & n1560 ) ;
  assign n1562 = ~n1554 & n1561 ;
  assign n1563 = x861 & ~n1444 ;
  assign n1564 = x241 & n1512 ;
  assign n1565 = ~x270 & n1520 ;
  assign n1566 = x171 & ~n1565 ;
  assign n1567 = ( n1526 & n1565 ) | ( n1526 & ~n1566 ) | ( n1565 & ~n1566 ) ;
  assign n1568 = x935 & n1502 ;
  assign n1569 = x1141 & ~n1502 ;
  assign n1570 = ( n1517 & n1568 ) | ( n1517 & n1569 ) | ( n1568 & n1569 ) ;
  assign n1571 = n1567 | n1570 ;
  assign n1572 = ( ~n1563 & n1564 ) | ( ~n1563 & n1571 ) | ( n1564 & n1571 ) ;
  assign n1573 = n1563 | n1572 ;
  assign n1574 = x869 & ~n1444 ;
  assign n1575 = x248 & n1512 ;
  assign n1576 = x921 & n1518 ;
  assign n1577 = x170 & ~n1576 ;
  assign n1578 = ( n1526 & n1576 ) | ( n1526 & ~n1577 ) | ( n1576 & ~n1577 ) ;
  assign n1579 = x1140 & n1523 ;
  assign n1580 = ~x282 & n1520 ;
  assign n1581 = ( ~n1578 & n1579 ) | ( ~n1578 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = n1578 | n1581 ;
  assign n1583 = ( ~n1574 & n1575 ) | ( ~n1574 & n1582 ) | ( n1575 & n1582 ) ;
  assign n1584 = n1574 | n1583 ;
  assign n1585 = x920 & n1518 ;
  assign n1586 = ~x281 & n1520 ;
  assign n1587 = x1139 & n1523 ;
  assign n1588 = ( ~n1585 & n1586 ) | ( ~n1585 & n1587 ) | ( n1586 & n1587 ) ;
  assign n1589 = n1585 | n1588 ;
  assign n1590 = x148 & ~n1589 ;
  assign n1591 = ( n1526 & n1589 ) | ( n1526 & ~n1590 ) | ( n1589 & ~n1590 ) ;
  assign n1592 = x862 | n1591 ;
  assign n1593 = ( ~n1444 & n1591 ) | ( ~n1444 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = x247 & n1512 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = ~x269 & n1520 ;
  assign n1597 = x246 | n1596 ;
  assign n1598 = ( n1512 & n1596 ) | ( n1512 & n1597 ) | ( n1596 & n1597 ) ;
  assign n1599 = x940 & n1502 ;
  assign n1600 = x1138 & ~n1502 ;
  assign n1601 = ( n1517 & n1599 ) | ( n1517 & n1600 ) | ( n1599 & n1600 ) ;
  assign n1602 = x169 & ~n1601 ;
  assign n1603 = ( n1526 & n1601 ) | ( n1526 & ~n1602 ) | ( n1601 & ~n1602 ) ;
  assign n1604 = x877 | n1603 ;
  assign n1605 = ( ~n1444 & n1603 ) | ( ~n1444 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = n1598 | n1605 ;
  assign n1607 = x878 & ~n1444 ;
  assign n1608 = x240 & n1512 ;
  assign n1609 = x933 & n1518 ;
  assign n1610 = x168 & ~n1609 ;
  assign n1611 = ( n1526 & n1609 ) | ( n1526 & ~n1610 ) | ( n1609 & ~n1610 ) ;
  assign n1612 = x1137 & n1523 ;
  assign n1613 = ~x280 & n1520 ;
  assign n1614 = ( ~n1611 & n1612 ) | ( ~n1611 & n1613 ) | ( n1612 & n1613 ) ;
  assign n1615 = n1611 | n1614 ;
  assign n1616 = ( ~n1607 & n1608 ) | ( ~n1607 & n1615 ) | ( n1608 & n1615 ) ;
  assign n1617 = n1607 | n1616 ;
  assign n1618 = x875 & ~n1444 ;
  assign n1619 = x245 & n1512 ;
  assign n1620 = x266 & n1520 ;
  assign n1621 = x166 | n1620 ;
  assign n1622 = ( n1526 & n1620 ) | ( n1526 & n1621 ) | ( n1620 & n1621 ) ;
  assign n1623 = x928 & n1502 ;
  assign n1624 = x1136 & ~n1502 ;
  assign n1625 = ( n1517 & n1623 ) | ( n1517 & n1624 ) | ( n1623 & n1624 ) ;
  assign n1626 = n1622 | n1625 ;
  assign n1627 = ( ~n1618 & n1619 ) | ( ~n1618 & n1626 ) | ( n1619 & n1626 ) ;
  assign n1628 = n1618 | n1627 ;
  assign n1629 = ~x938 & n1518 ;
  assign n1630 = ~x279 & n1520 ;
  assign n1631 = ~x1135 & n1523 ;
  assign n1632 = ( ~n1629 & n1630 ) | ( ~n1629 & n1631 ) | ( n1630 & n1631 ) ;
  assign n1633 = n1629 | n1632 ;
  assign n1634 = x879 & ~n1633 ;
  assign n1635 = ( n1444 & ~n1633 ) | ( n1444 & n1634 ) | ( ~n1633 & n1634 ) ;
  assign n1636 = ~x161 & n1526 ;
  assign n1637 = x244 & ~n1636 ;
  assign n1638 = ( n1512 & n1636 ) | ( n1512 & ~n1637 ) | ( n1636 & ~n1637 ) ;
  assign n1639 = n1635 & ~n1638 ;
  assign n1640 = x278 & n1520 ;
  assign n1641 = x242 | n1640 ;
  assign n1642 = ( n1512 & n1640 ) | ( n1512 & n1641 ) | ( n1640 & n1641 ) ;
  assign n1643 = x930 & n1502 ;
  assign n1644 = x1134 & ~n1502 ;
  assign n1645 = ( n1517 & n1643 ) | ( n1517 & n1644 ) | ( n1643 & n1644 ) ;
  assign n1646 = x152 | n1645 ;
  assign n1647 = ( n1526 & n1645 ) | ( n1526 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = x846 | n1647 ;
  assign n1649 = ( ~n1444 & n1647 ) | ( ~n1444 & n1648 ) | ( n1647 & n1648 ) ;
  assign n1650 = n1642 | n1649 ;
  assign n1651 = ~x215 & x299 ;
  assign n1652 = ( x39 & ~n1426 ) | ( x39 & n1651 ) | ( ~n1426 & n1651 ) ;
  assign n1653 = x74 | n1652 ;
  assign n1654 = x661 | x662 ;
  assign n1655 = x681 | n1654 ;
  assign n1656 = x680 & ~n1655 ;
  assign n1657 = x614 | x616 ;
  assign n1658 = x642 | n1657 ;
  assign n1659 = x603 & ~n1658 ;
  assign n1660 = n1656 | n1659 ;
  assign n1661 = x332 | x468 ;
  assign n1662 = n1660 & n1661 ;
  assign n1663 = x975 | x978 ;
  assign n1664 = x907 | x947 ;
  assign n1665 = ( ~x960 & n1663 ) | ( ~x960 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1666 = x970 | x972 ;
  assign n1667 = x960 | n1666 ;
  assign n1668 = n1665 | n1667 ;
  assign n1669 = x963 | n1668 ;
  assign n1670 = x969 | x971 ;
  assign n1671 = x587 | x602 ;
  assign n1672 = x961 | x967 ;
  assign n1673 = ( ~n1670 & n1671 ) | ( ~n1670 & n1672 ) | ( n1671 & n1672 ) ;
  assign n1674 = x974 | x977 ;
  assign n1675 = n1670 | n1674 ;
  assign n1676 = n1673 | n1675 ;
  assign n1677 = x299 | n1676 ;
  assign n1678 = ~x299 & n1676 ;
  assign n1679 = ( n1669 & n1677 ) | ( n1669 & n1678 ) | ( n1677 & n1678 ) ;
  assign n1680 = ~n1660 & n1661 ;
  assign n1681 = ( n1662 & n1679 ) | ( n1662 & ~n1680 ) | ( n1679 & ~n1680 ) ;
  assign n1682 = x252 | x1001 ;
  assign n1683 = x979 | x984 ;
  assign n1684 = ( x835 & x979 ) | ( x835 & n1683 ) | ( x979 & n1683 ) ;
  assign n1685 = n1682 & ~n1684 ;
  assign n1686 = x835 & n1685 ;
  assign n1687 = ~x287 & n1686 ;
  assign n1688 = n1681 & n1687 ;
  assign n1689 = x824 & x1092 ;
  assign n1690 = n1469 & n1689 ;
  assign n1691 = n1470 | n1690 ;
  assign n1692 = n1688 & n1691 ;
  assign n1693 = x39 & ~n1692 ;
  assign n1694 = n1653 | n1693 ;
  assign n1695 = ~n1416 & n1694 ;
  assign n1696 = x93 & x841 ;
  assign n1697 = n1450 | n1696 ;
  assign n1698 = n1280 & n1485 ;
  assign n1699 = ( n1484 & ~n1485 ) | ( n1484 & n1698 ) | ( ~n1485 & n1698 ) ;
  assign n1700 = ( n1486 & ~n1697 ) | ( n1486 & n1699 ) | ( ~n1697 & n1699 ) ;
  assign n1701 = x87 | n1382 ;
  assign n1702 = ~n1405 & n1701 ;
  assign n1703 = n1700 | n1702 ;
  assign n1704 = n1695 | n1703 ;
  assign n1705 = x222 & ~n1426 ;
  assign n1706 = x221 & n1651 ;
  assign n1707 = n1705 | n1706 ;
  assign n1708 = x39 & n1707 ;
  assign n1709 = x216 & x299 ;
  assign n1710 = x224 & ~x299 ;
  assign n1711 = n1709 | n1710 ;
  assign n1712 = n1708 & n1711 ;
  assign n1713 = ~n1416 & n1712 ;
  assign n1714 = x1093 & n1470 ;
  assign n1715 = n1688 & n1714 ;
  assign n1716 = n1713 & n1715 ;
  assign n1717 = x44 | x114 ;
  assign n1718 = x101 | x113 ;
  assign n1719 = x41 | x42 ;
  assign n1720 = ( ~x43 & n1718 ) | ( ~x43 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1721 = x52 | x99 ;
  assign n1722 = x43 | n1721 ;
  assign n1723 = n1720 | n1722 ;
  assign n1724 = x115 | x116 ;
  assign n1725 = ( ~n1717 & n1723 ) | ( ~n1717 & n1724 ) | ( n1723 & n1724 ) ;
  assign n1726 = n1717 | n1725 ;
  assign n1727 = x232 & ~n1661 ;
  assign n1728 = ~n1460 & n1727 ;
  assign n1729 = n1726 & ~n1728 ;
  assign n1730 = n1468 & n1689 ;
  assign n1731 = n1464 & n1468 ;
  assign n1732 = n1730 | n1731 ;
  assign n1733 = x250 | n1732 ;
  assign n1734 = x129 & x250 ;
  assign n1735 = ( n1461 & ~n1733 ) | ( n1461 & n1734 ) | ( ~n1733 & n1734 ) ;
  assign n1736 = x683 & n1735 ;
  assign n1737 = n1729 & n1736 ;
  assign n1738 = x100 & ~x252 ;
  assign n1739 = ( x100 & n1461 ) | ( x100 & n1738 ) | ( n1461 & n1738 ) ;
  assign n1740 = ~n1737 & n1739 ;
  assign n1741 = x1093 & n1691 ;
  assign n1742 = n1687 & n1741 ;
  assign n1743 = x829 & x1091 ;
  assign n1744 = ( n1708 & n1712 ) | ( n1708 & ~n1743 ) | ( n1712 & ~n1743 ) ;
  assign n1745 = n1208 & ~n1744 ;
  assign n1746 = ( n1208 & ~n1742 ) | ( n1208 & n1745 ) | ( ~n1742 & n1745 ) ;
  assign n1747 = n1740 | n1746 ;
  assign n1748 = x100 & ~n1747 ;
  assign n1749 = ( n1716 & ~n1747 ) | ( n1716 & n1748 ) | ( ~n1747 & n1748 ) ;
  assign n1750 = n1704 & ~n1749 ;
  assign n1751 = x82 | n1431 ;
  assign n1752 = x66 | x67 ;
  assign n1753 = ( x81 & n1213 ) | ( x81 & ~n1752 ) | ( n1213 & ~n1752 ) ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1235 | n1754 ;
  assign n1756 = x103 & ~x314 ;
  assign n1757 = ( ~n1751 & n1755 ) | ( ~n1751 & n1756 ) | ( n1755 & n1756 ) ;
  assign n1758 = n1751 | n1757 ;
  assign n1759 = x72 & ~n1389 ;
  assign n1760 = x197 & x299 ;
  assign n1761 = x145 & ~x299 ;
  assign n1762 = ( n1727 & n1760 ) | ( n1727 & n1761 ) | ( n1760 & n1761 ) ;
  assign n1763 = x109 & ~n1762 ;
  assign n1764 = x158 & x299 ;
  assign n1765 = x180 & ~x299 ;
  assign n1766 = n1764 | n1765 ;
  assign n1767 = x182 & ~x299 ;
  assign n1768 = x160 & x299 ;
  assign n1769 = n1767 | n1768 ;
  assign n1770 = n1766 & n1769 ;
  assign n1771 = x159 & x299 ;
  assign n1772 = x181 & ~x299 ;
  assign n1773 = n1771 | n1772 ;
  assign n1774 = n1770 & n1773 ;
  assign n1775 = ( x109 & n1763 ) | ( x109 & ~n1774 ) | ( n1763 & ~n1774 ) ;
  assign n1776 = n1697 | n1775 ;
  assign n1777 = ( ~n1758 & n1759 ) | ( ~n1758 & n1776 ) | ( n1759 & n1776 ) ;
  assign n1778 = ( ~n1484 & n1758 ) | ( ~n1484 & n1777 ) | ( n1758 & n1777 ) ;
  assign n1779 = n1484 | n1778 ;
  assign n1780 = ( n1484 & n1485 ) | ( n1484 & n1779 ) | ( n1485 & n1779 ) ;
  assign n1781 = n1491 & ~n1747 ;
  assign n1782 = n1780 | n1781 ;
  assign n1783 = ~x30 & x228 ;
  assign n1784 = x30 & x228 ;
  assign n1785 = ( n1782 & ~n1783 ) | ( n1782 & n1784 ) | ( ~n1783 & n1784 ) ;
  assign n1786 = n1656 & n1661 ;
  assign n1787 = ~n1656 & n1661 ;
  assign n1788 = x602 & ~n1421 ;
  assign n1789 = x907 & n1421 ;
  assign n1790 = n1788 | n1789 ;
  assign n1791 = ( n1786 & ~n1787 ) | ( n1786 & n1790 ) | ( ~n1787 & n1790 ) ;
  assign n1792 = n1785 & n1791 ;
  assign n1793 = x587 | n1421 ;
  assign n1794 = n1659 & n1661 ;
  assign n1795 = ~x947 & n1421 ;
  assign n1796 = ( n1661 & ~n1794 ) | ( n1661 & n1795 ) | ( ~n1794 & n1795 ) ;
  assign n1797 = ( n1793 & n1794 ) | ( n1793 & ~n1796 ) | ( n1794 & ~n1796 ) ;
  assign n1798 = n1785 & n1797 ;
  assign n1799 = ~n1661 & n1785 ;
  assign n1800 = x967 & ~n1421 ;
  assign n1801 = x970 & n1421 ;
  assign n1802 = ( n1799 & n1800 ) | ( n1799 & n1801 ) | ( n1800 & n1801 ) ;
  assign n1803 = x961 & ~n1421 ;
  assign n1804 = x972 & n1421 ;
  assign n1805 = ( n1799 & n1803 ) | ( n1799 & n1804 ) | ( n1803 & n1804 ) ;
  assign n1806 = x977 & ~n1421 ;
  assign n1807 = x960 & n1421 ;
  assign n1808 = ( n1799 & n1806 ) | ( n1799 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = x969 & ~n1421 ;
  assign n1810 = x963 & n1421 ;
  assign n1811 = ( n1799 & n1809 ) | ( n1799 & n1810 ) | ( n1809 & n1810 ) ;
  assign n1812 = x971 & ~n1421 ;
  assign n1813 = x975 & n1421 ;
  assign n1814 = ( n1799 & n1812 ) | ( n1799 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = x974 & ~n1421 ;
  assign n1816 = x978 & n1421 ;
  assign n1817 = ( n1799 & n1815 ) | ( n1799 & n1816 ) | ( n1815 & n1816 ) ;
  assign n1818 = ~n1693 & n1782 ;
  assign n1819 = ~x24 & x954 ;
  assign n1820 = x24 & x954 ;
  assign n1821 = ( n1818 & n1819 ) | ( n1818 & ~n1820 ) | ( n1819 & ~n1820 ) ;
  assign n1822 = ~n1407 & n1418 ;
  assign n1823 = n1414 | n1822 ;
  assign n1824 = n1208 | n1739 ;
  assign n1825 = ( n1485 & n1489 ) | ( n1485 & ~n1490 ) | ( n1489 & ~n1490 ) ;
  assign n1826 = ( n1485 & n1824 ) | ( n1485 & n1825 ) | ( n1824 & n1825 ) ;
  assign n1827 = n1823 | n1826 ;
  assign n1828 = ( n1205 & ~n1419 ) | ( n1205 & n1827 ) | ( ~n1419 & n1827 ) ;
  assign n1829 = x119 | x468 ;
  assign n1830 = n1440 & ~n1829 ;
  assign n1831 = x119 & ~x468 ;
  assign n1832 = ~x1056 & n1831 ;
  assign n1833 = n1830 | n1832 ;
  assign n1834 = ~x1077 & n1831 ;
  assign n1835 = n1830 | n1834 ;
  assign n1836 = ~x1073 & n1831 ;
  assign n1837 = n1830 | n1836 ;
  assign n1838 = ~x1041 & n1831 ;
  assign n1839 = n1830 | n1838 ;
  assign n1840 = x1161 & x1162 ;
  assign n1841 = x1092 & x1093 ;
  assign n1842 = ( x1163 & n1840 ) | ( x1163 & ~n1841 ) | ( n1840 & ~n1841 ) ;
  assign n1843 = n1840 & ~n1842 ;
  assign n1844 = ~x31 & n1843 ;
  assign n1845 = ~x24 & x91 ;
  assign n1846 = n1714 & n1845 ;
  assign n1847 = ~x122 & n1474 ;
  assign n1848 = ( ~x122 & n1846 ) | ( ~x122 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1849 = ~x841 & n1258 ;
  assign n1850 = x51 | x98 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = n1848 | n1851 ;
  assign n1853 = n1368 & n1852 ;
  assign n1854 = n1707 & ~n1711 ;
  assign n1855 = x39 & ~n1854 ;
  assign n1856 = ( x39 & ~n1715 ) | ( x39 & n1855 ) | ( ~n1715 & n1855 ) ;
  assign n1857 = n1691 & ~n1856 ;
  assign n1858 = x122 | n1732 ;
  assign n1859 = ~x24 & x75 ;
  assign n1860 = x100 | x252 ;
  assign n1861 = ( x100 & n1859 ) | ( x100 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1862 = ( n1470 & n1858 ) | ( n1470 & n1861 ) | ( n1858 & n1861 ) ;
  assign n1863 = ~n1858 & n1862 ;
  assign n1864 = n1729 & n1863 ;
  assign n1865 = x228 | n1397 ;
  assign n1866 = ( n1206 & n1864 ) | ( n1206 & n1865 ) | ( n1864 & n1865 ) ;
  assign n1867 = n1857 & n1866 ;
  assign n1868 = ( n1853 & n1857 ) | ( n1853 & n1867 ) | ( n1857 & n1867 ) ;
  assign n1869 = ~n1417 & n1868 ;
  assign n1870 = x824 & x950 ;
  assign n1871 = ~x1091 & n1841 ;
  assign n1872 = n1870 & n1871 ;
  assign n1873 = x286 | x288 ;
  assign n1874 = x285 | x289 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = ~x122 & n1875 ;
  assign n1877 = n1872 & n1876 ;
  assign n1878 = n1869 | n1877 ;
  assign n1879 = ~x98 & x567 ;
  assign n1880 = n1841 & ~n1879 ;
  assign n1881 = x590 | x592 ;
  assign n1882 = x588 & ~x591 ;
  assign n1883 = ( ~x426 & x428 ) | ( ~x426 & x430 ) | ( x428 & x430 ) ;
  assign n1884 = ( x426 & x428 ) | ( x426 & x430 ) | ( x428 & x430 ) ;
  assign n1885 = ( x426 & n1883 ) | ( x426 & ~n1884 ) | ( n1883 & ~n1884 ) ;
  assign n1886 = ( x427 & ~x451 ) | ( x427 & n1885 ) | ( ~x451 & n1885 ) ;
  assign n1887 = ( x427 & x451 ) | ( x427 & ~n1885 ) | ( x451 & ~n1885 ) ;
  assign n1888 = ( ~x427 & n1886 ) | ( ~x427 & n1887 ) | ( n1886 & n1887 ) ;
  assign n1889 = x433 & x445 ;
  assign n1890 = x433 | x445 ;
  assign n1891 = ~n1889 & n1890 ;
  assign n1892 = ( x448 & ~x449 ) | ( x448 & n1891 ) | ( ~x449 & n1891 ) ;
  assign n1893 = ( x448 & x449 ) | ( x448 & ~n1891 ) | ( x449 & ~n1891 ) ;
  assign n1894 = ( ~x448 & n1892 ) | ( ~x448 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1895 = ( x1199 & n1888 ) | ( x1199 & n1894 ) | ( n1888 & n1894 ) ;
  assign n1896 = ( ~x1199 & n1888 ) | ( ~x1199 & n1894 ) | ( n1888 & n1894 ) ;
  assign n1897 = n1895 & ~n1896 ;
  assign n1898 = x419 & x432 ;
  assign n1899 = x419 | x432 ;
  assign n1900 = ~n1898 & n1899 ;
  assign n1901 = ( x454 & ~x459 ) | ( x454 & n1900 ) | ( ~x459 & n1900 ) ;
  assign n1902 = ( x454 & x459 ) | ( x454 & ~n1900 ) | ( x459 & ~n1900 ) ;
  assign n1903 = ( ~x454 & n1901 ) | ( ~x454 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = ( x423 & ~x425 ) | ( x423 & n1903 ) | ( ~x425 & n1903 ) ;
  assign n1905 = ( x423 & x425 ) | ( x423 & ~n1903 ) | ( x425 & ~n1903 ) ;
  assign n1906 = ( ~x423 & n1904 ) | ( ~x423 & n1905 ) | ( n1904 & n1905 ) ;
  assign n1907 = ( ~x420 & x421 ) | ( ~x420 & x424 ) | ( x421 & x424 ) ;
  assign n1908 = ( x420 & x421 ) | ( x420 & x424 ) | ( x421 & x424 ) ;
  assign n1909 = ( x420 & n1907 ) | ( x420 & ~n1908 ) | ( n1907 & ~n1908 ) ;
  assign n1910 = ( x1198 & n1906 ) | ( x1198 & n1909 ) | ( n1906 & n1909 ) ;
  assign n1911 = n1906 & n1909 ;
  assign n1912 = ( n1897 & n1910 ) | ( n1897 & ~n1911 ) | ( n1910 & ~n1911 ) ;
  assign n1913 = ( ~x414 & x429 ) | ( ~x414 & x446 ) | ( x429 & x446 ) ;
  assign n1914 = ( x414 & x429 ) | ( x414 & x446 ) | ( x429 & x446 ) ;
  assign n1915 = ( x414 & n1913 ) | ( x414 & ~n1914 ) | ( n1913 & ~n1914 ) ;
  assign n1916 = ( x422 & ~x434 ) | ( x422 & n1915 ) | ( ~x434 & n1915 ) ;
  assign n1917 = ( x422 & x434 ) | ( x422 & ~n1915 ) | ( x434 & ~n1915 ) ;
  assign n1918 = ( ~x422 & n1916 ) | ( ~x422 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = x435 & x436 ;
  assign n1920 = x435 | x436 ;
  assign n1921 = ~n1919 & n1920 ;
  assign n1922 = ( x443 & ~x444 ) | ( x443 & n1921 ) | ( ~x444 & n1921 ) ;
  assign n1923 = ( x443 & x444 ) | ( x443 & ~n1921 ) | ( x444 & ~n1921 ) ;
  assign n1924 = ( ~x443 & n1922 ) | ( ~x443 & n1923 ) | ( n1922 & n1923 ) ;
  assign n1925 = ( x1196 & n1918 ) | ( x1196 & n1924 ) | ( n1918 & n1924 ) ;
  assign n1926 = ( ~x1196 & n1918 ) | ( ~x1196 & n1924 ) | ( n1918 & n1924 ) ;
  assign n1927 = n1925 & ~n1926 ;
  assign n1928 = x431 & x437 ;
  assign n1929 = x431 | x437 ;
  assign n1930 = ~n1928 & n1929 ;
  assign n1931 = ( x438 & ~x464 ) | ( x438 & n1930 ) | ( ~x464 & n1930 ) ;
  assign n1932 = ( x438 & x464 ) | ( x438 & ~n1930 ) | ( x464 & ~n1930 ) ;
  assign n1933 = ( ~x438 & n1931 ) | ( ~x438 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1934 = ( x415 & ~x416 ) | ( x415 & n1933 ) | ( ~x416 & n1933 ) ;
  assign n1935 = ( x415 & x416 ) | ( x415 & ~n1933 ) | ( x416 & ~n1933 ) ;
  assign n1936 = ( ~x415 & n1934 ) | ( ~x415 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1937 = ( ~x417 & x418 ) | ( ~x417 & x453 ) | ( x418 & x453 ) ;
  assign n1938 = ( x417 & x418 ) | ( x417 & x453 ) | ( x418 & x453 ) ;
  assign n1939 = ( x417 & n1937 ) | ( x417 & ~n1938 ) | ( n1937 & ~n1938 ) ;
  assign n1940 = ( x1197 & n1936 ) | ( x1197 & n1939 ) | ( n1936 & n1939 ) ;
  assign n1941 = n1936 & n1939 ;
  assign n1942 = ( n1927 & n1940 ) | ( n1927 & ~n1941 ) | ( n1940 & ~n1941 ) ;
  assign n1943 = n1912 | n1942 ;
  assign n1944 = n1882 & n1943 ;
  assign n1945 = ~x588 & x591 ;
  assign n1946 = x391 & x407 ;
  assign n1947 = x391 | x407 ;
  assign n1948 = ~n1946 & n1947 ;
  assign n1949 = ( x413 & ~x463 ) | ( x413 & n1948 ) | ( ~x463 & n1948 ) ;
  assign n1950 = ( x413 & x463 ) | ( x413 & ~n1948 ) | ( x463 & ~n1948 ) ;
  assign n1951 = ( ~x413 & n1949 ) | ( ~x413 & n1950 ) | ( n1949 & n1950 ) ;
  assign n1952 = ( x334 & ~x335 ) | ( x334 & n1951 ) | ( ~x335 & n1951 ) ;
  assign n1953 = ( x334 & x335 ) | ( x334 & ~n1951 ) | ( x335 & ~n1951 ) ;
  assign n1954 = ( ~x334 & n1952 ) | ( ~x334 & n1953 ) | ( n1952 & n1953 ) ;
  assign n1955 = ( ~x333 & x392 ) | ( ~x333 & x393 ) | ( x392 & x393 ) ;
  assign n1956 = ( x333 & x392 ) | ( x333 & x393 ) | ( x392 & x393 ) ;
  assign n1957 = ( x333 & n1955 ) | ( x333 & ~n1956 ) | ( n1955 & ~n1956 ) ;
  assign n1958 = ( ~x1197 & n1954 ) | ( ~x1197 & n1957 ) | ( n1954 & n1957 ) ;
  assign n1959 = ( x1197 & n1954 ) | ( x1197 & n1957 ) | ( n1954 & n1957 ) ;
  assign n1960 = ~n1958 & n1959 ;
  assign n1961 = x329 & x395 ;
  assign n1962 = x329 | x395 ;
  assign n1963 = ~n1961 & n1962 ;
  assign n1964 = ( x400 & ~x408 ) | ( x400 & n1963 ) | ( ~x408 & n1963 ) ;
  assign n1965 = ( x400 & x408 ) | ( x400 & ~n1963 ) | ( x408 & ~n1963 ) ;
  assign n1966 = ( ~x400 & n1964 ) | ( ~x400 & n1965 ) | ( n1964 & n1965 ) ;
  assign n1967 = ( x396 & ~x399 ) | ( x396 & n1966 ) | ( ~x399 & n1966 ) ;
  assign n1968 = ( x396 & x399 ) | ( x396 & ~n1966 ) | ( x399 & ~n1966 ) ;
  assign n1969 = ( ~x396 & n1967 ) | ( ~x396 & n1968 ) | ( n1967 & n1968 ) ;
  assign n1970 = ( ~x328 & x394 ) | ( ~x328 & x398 ) | ( x394 & x398 ) ;
  assign n1971 = ( x328 & x394 ) | ( x328 & x398 ) | ( x394 & x398 ) ;
  assign n1972 = ( x328 & n1970 ) | ( x328 & ~n1971 ) | ( n1970 & ~n1971 ) ;
  assign n1973 = ( x1198 & n1969 ) | ( x1198 & n1972 ) | ( n1969 & n1972 ) ;
  assign n1974 = n1969 & n1972 ;
  assign n1975 = ( n1960 & n1973 ) | ( n1960 & ~n1974 ) | ( n1973 & ~n1974 ) ;
  assign n1976 = x402 & x403 ;
  assign n1977 = x402 | x403 ;
  assign n1978 = ~n1976 & n1977 ;
  assign n1979 = x325 & x326 ;
  assign n1980 = x325 | x326 ;
  assign n1981 = ~n1979 & n1980 ;
  assign n1982 = ( ~x318 & x401 ) | ( ~x318 & x405 ) | ( x401 & x405 ) ;
  assign n1983 = ( x318 & x401 ) | ( x318 & x405 ) | ( x401 & x405 ) ;
  assign n1984 = ( x318 & n1982 ) | ( x318 & ~n1983 ) | ( n1982 & ~n1983 ) ;
  assign n1985 = ( n1978 & ~n1981 ) | ( n1978 & n1984 ) | ( ~n1981 & n1984 ) ;
  assign n1986 = ( n1978 & n1981 ) | ( n1978 & ~n1984 ) | ( n1981 & ~n1984 ) ;
  assign n1987 = ( ~n1978 & n1985 ) | ( ~n1978 & n1986 ) | ( n1985 & n1986 ) ;
  assign n1988 = ( x406 & ~x409 ) | ( x406 & n1987 ) | ( ~x409 & n1987 ) ;
  assign n1989 = ( x406 & x409 ) | ( x406 & ~n1987 ) | ( x409 & ~n1987 ) ;
  assign n1990 = ( ~x406 & n1988 ) | ( ~x406 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1991 = x1199 & n1990 ;
  assign n1992 = ( ~x324 & x397 ) | ( ~x324 & x456 ) | ( x397 & x456 ) ;
  assign n1993 = ( x324 & x397 ) | ( x324 & x456 ) | ( x397 & x456 ) ;
  assign n1994 = ( x324 & n1992 ) | ( x324 & ~n1993 ) | ( n1992 & ~n1993 ) ;
  assign n1995 = ( x390 & ~x411 ) | ( x390 & n1994 ) | ( ~x411 & n1994 ) ;
  assign n1996 = ( x390 & x411 ) | ( x390 & ~n1994 ) | ( x411 & ~n1994 ) ;
  assign n1997 = ( ~x390 & n1995 ) | ( ~x390 & n1996 ) | ( n1995 & n1996 ) ;
  assign n1998 = x319 & x404 ;
  assign n1999 = x319 | x404 ;
  assign n2000 = ~n1998 & n1999 ;
  assign n2001 = ( x410 & ~x412 ) | ( x410 & n2000 ) | ( ~x412 & n2000 ) ;
  assign n2002 = ( x410 & x412 ) | ( x410 & ~n2000 ) | ( x412 & ~n2000 ) ;
  assign n2003 = ( ~x410 & n2001 ) | ( ~x410 & n2002 ) | ( n2001 & n2002 ) ;
  assign n2004 = ( x1196 & n1997 ) | ( x1196 & n2003 ) | ( n1997 & n2003 ) ;
  assign n2005 = n1997 & n2003 ;
  assign n2006 = ( n1991 & n2004 ) | ( n1991 & ~n2005 ) | ( n2004 & ~n2005 ) ;
  assign n2007 = n1945 & n2006 ;
  assign n2008 = ( n1945 & n1975 ) | ( n1945 & n2007 ) | ( n1975 & n2007 ) ;
  assign n2009 = n1944 | n2008 ;
  assign n2010 = ~n1881 & n2009 ;
  assign n2011 = x588 | x591 ;
  assign n2012 = x590 & ~x592 ;
  assign n2013 = ~n2011 & n2012 ;
  assign n2014 = ( ~x352 & x357 ) | ( ~x352 & x462 ) | ( x357 & x462 ) ;
  assign n2015 = ( x352 & x357 ) | ( x352 & x462 ) | ( x357 & x462 ) ;
  assign n2016 = ( x352 & n2014 ) | ( x352 & ~n2015 ) | ( n2014 & ~n2015 ) ;
  assign n2017 = ( x351 & ~x461 ) | ( x351 & n2016 ) | ( ~x461 & n2016 ) ;
  assign n2018 = ( x351 & x461 ) | ( x351 & ~n2016 ) | ( x461 & ~n2016 ) ;
  assign n2019 = ( ~x351 & n2017 ) | ( ~x351 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2020 = x353 & x354 ;
  assign n2021 = x353 | x354 ;
  assign n2022 = ~n2020 & n2021 ;
  assign n2023 = ( x356 & ~x360 ) | ( x356 & n2022 ) | ( ~x360 & n2022 ) ;
  assign n2024 = ( x356 & x360 ) | ( x356 & ~n2022 ) | ( x360 & ~n2022 ) ;
  assign n2025 = ( ~x356 & n2023 ) | ( ~x356 & n2024 ) | ( n2023 & n2024 ) ;
  assign n2026 = ( x1199 & n2019 ) | ( x1199 & n2025 ) | ( n2019 & n2025 ) ;
  assign n2027 = ( ~x1199 & n2019 ) | ( ~x1199 & n2025 ) | ( n2019 & n2025 ) ;
  assign n2028 = n2026 & ~n2027 ;
  assign n2029 = ( ~x327 & x344 ) | ( ~x327 & x362 ) | ( x344 & x362 ) ;
  assign n2030 = ( x327 & x344 ) | ( x327 & x362 ) | ( x344 & x362 ) ;
  assign n2031 = ( x327 & n2029 ) | ( x327 & ~n2030 ) | ( n2029 & ~n2030 ) ;
  assign n2032 = ( x343 & ~x345 ) | ( x343 & n2031 ) | ( ~x345 & n2031 ) ;
  assign n2033 = ( x343 & x345 ) | ( x343 & ~n2031 ) | ( x345 & ~n2031 ) ;
  assign n2034 = ( ~x343 & n2032 ) | ( ~x343 & n2033 ) | ( n2032 & n2033 ) ;
  assign n2035 = x323 & x346 ;
  assign n2036 = x323 | x346 ;
  assign n2037 = ~n2035 & n2036 ;
  assign n2038 = ( x358 & ~x450 ) | ( x358 & n2037 ) | ( ~x450 & n2037 ) ;
  assign n2039 = ( x358 & x450 ) | ( x358 & ~n2037 ) | ( x450 & ~n2037 ) ;
  assign n2040 = ( ~x358 & n2038 ) | ( ~x358 & n2039 ) | ( n2038 & n2039 ) ;
  assign n2041 = ( x1197 & n2034 ) | ( x1197 & n2040 ) | ( n2034 & n2040 ) ;
  assign n2042 = n2034 & n2040 ;
  assign n2043 = ( n2028 & n2041 ) | ( n2028 & ~n2042 ) | ( n2041 & ~n2042 ) ;
  assign n2044 = x315 & x316 ;
  assign n2045 = x315 | x316 ;
  assign n2046 = ~n2044 & n2045 ;
  assign n2047 = ( x350 & ~x359 ) | ( x350 & n2046 ) | ( ~x359 & n2046 ) ;
  assign n2048 = ( x350 & x359 ) | ( x350 & ~n2046 ) | ( x359 & ~n2046 ) ;
  assign n2049 = ( ~x350 & n2047 ) | ( ~x350 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2050 = ( x321 & ~x322 ) | ( x321 & n2049 ) | ( ~x322 & n2049 ) ;
  assign n2051 = ( x321 & x322 ) | ( x321 & ~n2049 ) | ( x322 & ~n2049 ) ;
  assign n2052 = ( ~x321 & n2050 ) | ( ~x321 & n2051 ) | ( n2050 & n2051 ) ;
  assign n2053 = ( ~x347 & x348 ) | ( ~x347 & x349 ) | ( x348 & x349 ) ;
  assign n2054 = ( x347 & x348 ) | ( x347 & x349 ) | ( x348 & x349 ) ;
  assign n2055 = ( x347 & n2053 ) | ( x347 & ~n2054 ) | ( n2053 & ~n2054 ) ;
  assign n2056 = ( x1198 & n2052 ) | ( x1198 & n2055 ) | ( n2052 & n2055 ) ;
  assign n2057 = n2052 & n2055 ;
  assign n2058 = ( n2043 & n2056 ) | ( n2043 & ~n2057 ) | ( n2056 & ~n2057 ) ;
  assign n2059 = ( ~x355 & x361 ) | ( ~x355 & x455 ) | ( x361 & x455 ) ;
  assign n2060 = ( x355 & x361 ) | ( x355 & x455 ) | ( x361 & x455 ) ;
  assign n2061 = ( x355 & n2059 ) | ( x355 & ~n2060 ) | ( n2059 & ~n2060 ) ;
  assign n2062 = ( x342 & ~x441 ) | ( x342 & n2061 ) | ( ~x441 & n2061 ) ;
  assign n2063 = ( x342 & x441 ) | ( x342 & ~n2061 ) | ( x441 & ~n2061 ) ;
  assign n2064 = ( ~x342 & n2062 ) | ( ~x342 & n2063 ) | ( n2062 & n2063 ) ;
  assign n2065 = x320 & x452 ;
  assign n2066 = x320 | x452 ;
  assign n2067 = ~n2065 & n2066 ;
  assign n2068 = ( x458 & ~x460 ) | ( x458 & n2067 ) | ( ~x460 & n2067 ) ;
  assign n2069 = ( x458 & x460 ) | ( x458 & ~n2067 ) | ( x460 & ~n2067 ) ;
  assign n2070 = ( ~x458 & n2068 ) | ( ~x458 & n2069 ) | ( n2068 & n2069 ) ;
  assign n2071 = ( x1196 & n2064 ) | ( x1196 & n2070 ) | ( n2064 & n2070 ) ;
  assign n2072 = n2064 & n2070 ;
  assign n2073 = ( n2058 & n2071 ) | ( n2058 & ~n2072 ) | ( n2071 & ~n2072 ) ;
  assign n2074 = n2013 & ~n2073 ;
  assign n2075 = ( ~x317 & x377 ) | ( ~x317 & x385 ) | ( x377 & x385 ) ;
  assign n2076 = ( x317 & x377 ) | ( x317 & x385 ) | ( x377 & x385 ) ;
  assign n2077 = ( x317 & n2075 ) | ( x317 & ~n2076 ) | ( n2075 & ~n2076 ) ;
  assign n2078 = ( x376 & ~x378 ) | ( x376 & n2077 ) | ( ~x378 & n2077 ) ;
  assign n2079 = ( x376 & x378 ) | ( x376 & ~n2077 ) | ( x378 & ~n2077 ) ;
  assign n2080 = ( ~x376 & n2078 ) | ( ~x376 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2081 = x379 & x381 ;
  assign n2082 = x379 | x381 ;
  assign n2083 = ~n2081 & n2082 ;
  assign n2084 = ( x382 & ~x439 ) | ( x382 & n2083 ) | ( ~x439 & n2083 ) ;
  assign n2085 = ( x382 & x439 ) | ( x382 & ~n2083 ) | ( x439 & ~n2083 ) ;
  assign n2086 = ( ~x382 & n2084 ) | ( ~x382 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2087 = ( x1199 & n2080 ) | ( x1199 & n2086 ) | ( n2080 & n2086 ) ;
  assign n2088 = ( ~x1199 & n2080 ) | ( ~x1199 & n2086 ) | ( n2080 & n2086 ) ;
  assign n2089 = n2087 & ~n2088 ;
  assign n2090 = ( ~x364 & x366 ) | ( ~x364 & x368 ) | ( x366 & x368 ) ;
  assign n2091 = ( x364 & x366 ) | ( x364 & x368 ) | ( x366 & x368 ) ;
  assign n2092 = ( x364 & n2090 ) | ( x364 & ~n2091 ) | ( n2090 & ~n2091 ) ;
  assign n2093 = ( x365 & ~x367 ) | ( x365 & n2092 ) | ( ~x367 & n2092 ) ;
  assign n2094 = ( x365 & x367 ) | ( x365 & ~n2092 ) | ( x367 & ~n2092 ) ;
  assign n2095 = ( ~x365 & n2093 ) | ( ~x365 & n2094 ) | ( n2093 & n2094 ) ;
  assign n2096 = x336 & x383 ;
  assign n2097 = x336 | x383 ;
  assign n2098 = ~n2096 & n2097 ;
  assign n2099 = ( x389 & ~x447 ) | ( x389 & n2098 ) | ( ~x447 & n2098 ) ;
  assign n2100 = ( x389 & x447 ) | ( x389 & ~n2098 ) | ( x447 & ~n2098 ) ;
  assign n2101 = ( ~x389 & n2099 ) | ( ~x389 & n2100 ) | ( n2099 & n2100 ) ;
  assign n2102 = ( x1197 & n2095 ) | ( x1197 & n2101 ) | ( n2095 & n2101 ) ;
  assign n2103 = n2095 & n2101 ;
  assign n2104 = ( n2089 & n2102 ) | ( n2089 & ~n2103 ) | ( n2102 & ~n2103 ) ;
  assign n2105 = ( ~x373 & x384 ) | ( ~x373 & x440 ) | ( x384 & x440 ) ;
  assign n2106 = ( x373 & x384 ) | ( x373 & x440 ) | ( x384 & x440 ) ;
  assign n2107 = ( x373 & n2105 ) | ( x373 & ~n2106 ) | ( n2105 & ~n2106 ) ;
  assign n2108 = ( x375 & ~x442 ) | ( x375 & n2107 ) | ( ~x442 & n2107 ) ;
  assign n2109 = ( x375 & x442 ) | ( x375 & ~n2107 ) | ( x442 & ~n2107 ) ;
  assign n2110 = ( ~x375 & n2108 ) | ( ~x375 & n2109 ) | ( n2108 & n2109 ) ;
  assign n2111 = x369 & x370 ;
  assign n2112 = x369 | x370 ;
  assign n2113 = ~n2111 & n2112 ;
  assign n2114 = ( x371 & ~x374 ) | ( x371 & n2113 ) | ( ~x374 & n2113 ) ;
  assign n2115 = ( x371 & x374 ) | ( x371 & ~n2113 ) | ( x374 & ~n2113 ) ;
  assign n2116 = ( ~x371 & n2114 ) | ( ~x371 & n2115 ) | ( n2114 & n2115 ) ;
  assign n2117 = ( x1198 & n2110 ) | ( x1198 & n2116 ) | ( n2110 & n2116 ) ;
  assign n2118 = n2110 & n2116 ;
  assign n2119 = ( n2104 & n2117 ) | ( n2104 & ~n2118 ) | ( n2117 & ~n2118 ) ;
  assign n2120 = ( ~x337 & x339 ) | ( ~x337 & x363 ) | ( x339 & x363 ) ;
  assign n2121 = ( x337 & x339 ) | ( x337 & x363 ) | ( x339 & x363 ) ;
  assign n2122 = ( x337 & n2120 ) | ( x337 & ~n2121 ) | ( n2120 & ~n2121 ) ;
  assign n2123 = ( x338 & ~x387 ) | ( x338 & n2122 ) | ( ~x387 & n2122 ) ;
  assign n2124 = ( x338 & x387 ) | ( x338 & ~n2122 ) | ( x387 & ~n2122 ) ;
  assign n2125 = ( ~x338 & n2123 ) | ( ~x338 & n2124 ) | ( n2123 & n2124 ) ;
  assign n2126 = x372 & x380 ;
  assign n2127 = x372 | x380 ;
  assign n2128 = ~n2126 & n2127 ;
  assign n2129 = ( x386 & ~x388 ) | ( x386 & n2128 ) | ( ~x388 & n2128 ) ;
  assign n2130 = ( x386 & x388 ) | ( x386 & ~n2128 ) | ( x388 & ~n2128 ) ;
  assign n2131 = ( ~x386 & n2129 ) | ( ~x386 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2132 = ( x1196 & n2125 ) | ( x1196 & n2131 ) | ( n2125 & n2131 ) ;
  assign n2133 = n2125 & n2131 ;
  assign n2134 = ( n2119 & n2132 ) | ( n2119 & ~n2133 ) | ( n2132 & ~n2133 ) ;
  assign n2135 = ~x590 & x592 ;
  assign n2136 = ~n2011 & n2135 ;
  assign n2137 = n2013 | n2136 ;
  assign n2138 = ( n2013 & n2134 ) | ( n2013 & n2137 ) | ( n2134 & n2137 ) ;
  assign n2139 = ( n2010 & ~n2074 ) | ( n2010 & n2138 ) | ( ~n2074 & n2138 ) ;
  assign n2140 = n1872 & n2139 ;
  assign n2141 = x217 & ~n1880 ;
  assign n2142 = ( n1880 & n2140 ) | ( n1880 & ~n2141 ) | ( n2140 & ~n2141 ) ;
  assign n2143 = x1161 | x1162 ;
  assign n2144 = x1163 | n2143 ;
  assign n2145 = ~n1844 & n2144 ;
  assign n2146 = ( ~n1844 & n2142 ) | ( ~n1844 & n2145 ) | ( n2142 & n2145 ) ;
  assign n2147 = ( n1844 & n1878 ) | ( n1844 & ~n2146 ) | ( n1878 & ~n2146 ) ;
  assign n2148 = n1206 | n1373 ;
  assign n2149 = ~x24 & x38 ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = ~n1385 & n1859 ;
  assign n2152 = x252 & n2151 ;
  assign n2153 = n1729 & n2152 ;
  assign n2154 = ( n2150 & n2152 ) | ( n2150 & ~n2153 ) | ( n2152 & ~n2153 ) ;
  assign n2155 = x137 | n2154 ;
  assign n2156 = ~x38 & x100 ;
  assign n2157 = ~n1397 & n2156 ;
  assign n2158 = x129 & n2157 ;
  assign n2159 = ~n1461 & n2158 ;
  assign n2160 = x252 & n2159 ;
  assign n2161 = n1735 & n2157 ;
  assign n2162 = n2160 | n2161 ;
  assign n2163 = ~n1729 & n2162 ;
  assign n2164 = ~n1470 & n2151 ;
  assign n2165 = n1461 & n1726 ;
  assign n2166 = ( n2163 & n2164 ) | ( n2163 & ~n2165 ) | ( n2164 & ~n2165 ) ;
  assign n2167 = ~n2155 & n2166 ;
  assign n2168 = n1396 | n2167 ;
  assign n2169 = ~n1470 & n1875 ;
  assign n2170 = n1365 & ~n1482 ;
  assign n2171 = x76 & n2170 ;
  assign n2172 = ~n2169 & n2171 ;
  assign n2173 = x137 | n1447 ;
  assign n2174 = n2172 & ~n2173 ;
  assign n2175 = n1239 | n1383 ;
  assign n2176 = n1306 & ~n2175 ;
  assign n2177 = x24 | x841 ;
  assign n2178 = ( x841 & ~n1447 ) | ( x841 & n2177 ) | ( ~n1447 & n2177 ) ;
  assign n2179 = x50 | n1272 ;
  assign n2180 = n2178 & ~n2179 ;
  assign n2181 = x24 | n1285 ;
  assign n2182 = ( n1284 & ~n2180 ) | ( n1284 & n2181 ) | ( ~n2180 & n2181 ) ;
  assign n2183 = ( n2175 & ~n2176 ) | ( n2175 & n2182 ) | ( ~n2176 & n2182 ) ;
  assign n2184 = ( n1396 & n2176 ) | ( n1396 & n2183 ) | ( n2176 & n2183 ) ;
  assign n2185 = ( n2168 & n2174 ) | ( n2168 & ~n2184 ) | ( n2174 & ~n2184 ) ;
  assign n2186 = ~x33 & x954 ;
  assign n2187 = x34 | x79 ;
  assign n2188 = x118 | x139 ;
  assign n2189 = x195 | x196 ;
  assign n2190 = x138 | n2189 ;
  assign n2191 = n2188 | n2190 ;
  assign n2192 = n2187 | n2191 ;
  assign n2193 = x33 | n2192 ;
  assign n2194 = ( ~x33 & x954 ) | ( ~x33 & n2193 ) | ( x954 & n2193 ) ;
  assign n2195 = n1688 & n1741 ;
  assign n2196 = n1713 & n2195 ;
  assign n2197 = x40 | x74 ;
  assign n2198 = n1377 | n2197 ;
  assign n2199 = x63 | x107 ;
  assign n2200 = n2198 | n2199 ;
  assign n2201 = n1240 | n1450 ;
  assign n2202 = x58 | x90 ;
  assign n2203 = x90 & x841 ;
  assign n2204 = ( x73 & n2202 ) | ( x73 & ~n2203 ) | ( n2202 & ~n2203 ) ;
  assign n2205 = n2201 | n2204 ;
  assign n2206 = n1431 | n2205 ;
  assign n2207 = n2200 | n2206 ;
  assign n2208 = ( n1485 & n2200 ) | ( n1485 & n2207 ) | ( n2200 & n2207 ) ;
  assign n2209 = ( n1823 & ~n2196 ) | ( n1823 & n2208 ) | ( ~n2196 & n2208 ) ;
  assign n2210 = n2196 | n2209 ;
  assign n2211 = ( n2186 & n2194 ) | ( n2186 & ~n2210 ) | ( n2194 & ~n2210 ) ;
  assign n2212 = x95 & ~n1766 ;
  assign n2213 = ~x193 & n2202 ;
  assign n2214 = x183 | n2202 ;
  assign n2215 = ( x73 & ~n2213 ) | ( x73 & n2214 ) | ( ~n2213 & n2214 ) ;
  assign n2216 = ( x73 & x95 ) | ( x73 & ~x174 ) | ( x95 & ~x174 ) ;
  assign n2217 = x73 & ~n2216 ;
  assign n2218 = ( x95 & n2215 ) | ( x95 & ~n2217 ) | ( n2215 & ~n2217 ) ;
  assign n2219 = ~x299 & n2218 ;
  assign n2220 = x73 & x152 ;
  assign n2221 = x299 & ~n2220 ;
  assign n2222 = ~x172 & n2202 ;
  assign n2223 = n2221 & ~n2222 ;
  assign n2224 = x32 | x70 ;
  assign n2225 = ~x149 & n2224 ;
  assign n2226 = ( ~x149 & n1240 ) | ( ~x149 & n2225 ) | ( n1240 & n2225 ) ;
  assign n2227 = ( n2212 & n2223 ) | ( n2212 & n2226 ) | ( n2223 & n2226 ) ;
  assign n2228 = n2223 & ~n2227 ;
  assign n2229 = ( ~n2212 & n2219 ) | ( ~n2212 & n2228 ) | ( n2219 & n2228 ) ;
  assign n2230 = n2206 & ~n2229 ;
  assign n2231 = x154 & x299 ;
  assign n2232 = x176 & ~x299 ;
  assign n2233 = n2231 | n2232 ;
  assign n2234 = n1470 & ~n2233 ;
  assign n2235 = x152 & x299 ;
  assign n2236 = ( n1456 & ~n1470 ) | ( n1456 & n2235 ) | ( ~n1470 & n2235 ) ;
  assign n2237 = ( x39 & n2234 ) | ( x39 & n2236 ) | ( n2234 & n2236 ) ;
  assign n2238 = x38 | n2237 ;
  assign n2239 = n2230 | n2238 ;
  assign n2240 = ~n1417 & n2239 ;
  assign n2241 = x178 & x183 ;
  assign n2242 = ~n1421 & n1727 ;
  assign n2243 = n1373 & n2242 ;
  assign n2244 = ( x178 & x183 ) | ( x178 & n2243 ) | ( x183 & n2243 ) ;
  assign n2245 = ( n2240 & ~n2241 ) | ( n2240 & n2244 ) | ( ~n2241 & n2244 ) ;
  assign n2246 = ~x149 & n1380 ;
  assign n2247 = n1727 & n2233 ;
  assign n2248 = ( ~x92 & n1727 ) | ( ~x92 & n2247 ) | ( n1727 & n2247 ) ;
  assign n2249 = ( n2200 & ~n2246 ) | ( n2200 & n2248 ) | ( ~n2246 & n2248 ) ;
  assign n2250 = ~n2200 & n2249 ;
  assign n2251 = x191 & ~n1421 ;
  assign n2252 = x169 & n1421 ;
  assign n2253 = ( n1727 & n2251 ) | ( n1727 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2254 = x74 | n1373 ;
  assign n2255 = ( n1373 & n2253 ) | ( n1373 & n2254 ) | ( n2253 & n2254 ) ;
  assign n2256 = n2250 | n2255 ;
  assign n2257 = x186 & ~n1421 ;
  assign n2258 = x164 & n1421 ;
  assign n2259 = ( n1727 & n2257 ) | ( n1727 & n2258 ) | ( n2257 & n2258 ) ;
  assign n2260 = ~x74 & n1376 ;
  assign n2261 = n2259 & n2260 ;
  assign n2262 = n2256 | n2261 ;
  assign n2263 = n1421 & n1727 ;
  assign n2264 = n1373 & n2263 ;
  assign n2265 = ( x149 & x157 ) | ( x149 & n2264 ) | ( x157 & n2264 ) ;
  assign n2266 = x149 & x157 ;
  assign n2267 = ( n2262 & ~n2265 ) | ( n2262 & n2266 ) | ( ~n2265 & n2266 ) ;
  assign n2268 = ~n2245 & n2267 ;
  assign n2269 = n2210 & ~n2268 ;
  assign n2270 = ( ~n2186 & n2211 ) | ( ~n2186 & n2269 ) | ( n2211 & n2269 ) ;
  assign n2271 = x33 | x954 ;
  assign n2272 = x34 | n2271 ;
  assign n2273 = ( x34 & n2192 ) | ( x34 & ~n2271 ) | ( n2192 & ~n2271 ) ;
  assign n2274 = ( n2271 & ~n2272 ) | ( n2271 & n2273 ) | ( ~n2272 & n2273 ) ;
  assign n2275 = n2210 | n2274 ;
  assign n2276 = n1679 & n1712 ;
  assign n2277 = n1742 & n2276 ;
  assign n2278 = x155 & x299 ;
  assign n2279 = x177 & ~x299 ;
  assign n2280 = ( n1743 & n2278 ) | ( n1743 & n2279 ) | ( n2278 & n2279 ) ;
  assign n2281 = ( ~n1435 & n1457 ) | ( ~n1435 & n1743 ) | ( n1457 & n1743 ) ;
  assign n2282 = ( n2277 & n2280 ) | ( n2277 & ~n2281 ) | ( n2280 & ~n2281 ) ;
  assign n2283 = ~n1411 & n2282 ;
  assign n2284 = n2202 & ~n2203 ;
  assign n2285 = ~n1455 & n2284 ;
  assign n2286 = ( n1431 & n1771 ) | ( n1431 & n1772 ) | ( n1771 & n1772 ) ;
  assign n2287 = ( x73 & n1435 ) | ( x73 & ~n1457 ) | ( n1435 & ~n1457 ) ;
  assign n2288 = n2286 | n2287 ;
  assign n2289 = n2285 | n2288 ;
  assign n2290 = x140 & ~x299 ;
  assign n2291 = x162 & x299 ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = n2201 & n2292 ;
  assign n2294 = n2289 | n2293 ;
  assign n2295 = n1485 & n2294 ;
  assign n2296 = x38 & ~n1401 ;
  assign n2297 = x188 & ~n1421 ;
  assign n2298 = x167 & n1421 ;
  assign n2299 = ( n2260 & n2297 ) | ( n2260 & n2298 ) | ( n2297 & n2298 ) ;
  assign n2300 = n1373 | n2299 ;
  assign n2301 = x149 | x157 ;
  assign n2302 = ( x162 & x197 ) | ( x162 & n2301 ) | ( x197 & n2301 ) ;
  assign n2303 = ( ~x162 & x197 ) | ( ~x162 & n2301 ) | ( x197 & n2301 ) ;
  assign n2304 = ( x162 & ~n2302 ) | ( x162 & n2303 ) | ( ~n2302 & n2303 ) ;
  assign n2305 = n1421 & ~n2304 ;
  assign n2306 = x178 | x183 ;
  assign n2307 = ( x140 & x145 ) | ( x140 & n2306 ) | ( x145 & n2306 ) ;
  assign n2308 = ( ~x140 & x145 ) | ( ~x140 & n2306 ) | ( x145 & n2306 ) ;
  assign n2309 = ( x140 & ~n2307 ) | ( x140 & n2308 ) | ( ~n2307 & n2308 ) ;
  assign n2310 = n1421 | n2309 ;
  assign n2311 = ( n1373 & n2305 ) | ( n1373 & ~n2310 ) | ( n2305 & ~n2310 ) ;
  assign n2312 = x141 & ~n1421 ;
  assign n2313 = x148 & n1421 ;
  assign n2314 = ( x74 & n2312 ) | ( x74 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2315 = ~n2311 & n2314 ;
  assign n2316 = ( n2300 & ~n2311 ) | ( n2300 & n2315 ) | ( ~n2311 & n2315 ) ;
  assign n2317 = x162 | n2316 ;
  assign n2318 = ( n1414 & n2316 ) | ( n1414 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2319 = n2296 | n2318 ;
  assign n2320 = ( n2295 & ~n2296 ) | ( n2295 & n2319 ) | ( ~n2296 & n2319 ) ;
  assign n2321 = n2283 | n2320 ;
  assign n2322 = ( n1727 & n2278 ) | ( n1727 & n2279 ) | ( n2278 & n2279 ) ;
  assign n2323 = n1822 & n2322 ;
  assign n2324 = ( n1727 & n2321 ) | ( n1727 & n2323 ) | ( n2321 & n2323 ) ;
  assign n2325 = n2275 & ~n2324 ;
  assign n2326 = ~n1858 & n2173 ;
  assign n2327 = n2172 & n2326 ;
  assign n2328 = n2168 & ~n2327 ;
  assign n2329 = x683 & n1690 ;
  assign n2330 = x252 & ~n2329 ;
  assign n2331 = n2159 & ~n2330 ;
  assign n2332 = ( n2154 & n2166 ) | ( n2154 & ~n2331 ) | ( n2166 & ~n2331 ) ;
  assign n2333 = n2331 | n2332 ;
  assign n2334 = n1396 | n2333 ;
  assign n2335 = ~n2328 & n2334 ;
  assign n2336 = x54 & ~n1372 ;
  assign n2337 = ~n1407 & n2336 ;
  assign n2338 = ( n1394 & ~n1488 ) | ( n1394 & n2337 ) | ( ~n1488 & n2337 ) ;
  assign n2339 = x24 & n2338 ;
  assign n2340 = ( n2335 & n2338 ) | ( n2335 & ~n2339 ) | ( n2338 & ~n2339 ) ;
  assign n2341 = ~x24 & n1449 ;
  assign n2342 = x40 & x1082 ;
  assign n2343 = x93 | x841 ;
  assign n2344 = ~x35 & x841 ;
  assign n2345 = ( x58 & n2343 ) | ( x58 & ~n2344 ) | ( n2343 & ~n2344 ) ;
  assign n2346 = n2342 | n2345 ;
  assign n2347 = n2341 | n2346 ;
  assign n2348 = n1485 & n2347 ;
  assign n2349 = n2340 | n2348 ;
  assign n2350 = n1285 | n1383 ;
  assign n2351 = n1364 & ~n2350 ;
  assign n2352 = x36 & n2351 ;
  assign n2353 = x91 & ~n1482 ;
  assign n2354 = ~x24 & n1732 ;
  assign n2355 = n2353 & n2354 ;
  assign n2356 = ( n1732 & n2352 ) | ( n1732 & n2355 ) | ( n2352 & n2355 ) ;
  assign n2357 = x89 & x332 ;
  assign n2358 = x64 & ~x841 ;
  assign n2359 = ( ~x841 & n2357 ) | ( ~x841 & n2358 ) | ( n2357 & n2358 ) ;
  assign n2360 = n2351 & n2359 ;
  assign n2361 = x24 | n2360 ;
  assign n2362 = ( n2296 & n2360 ) | ( n2296 & n2361 ) | ( n2360 & n2361 ) ;
  assign n2363 = x986 | n1732 ;
  assign n2364 = x108 & x314 ;
  assign n2365 = ~x252 & n2364 ;
  assign n2366 = ( ~n2363 & n2364 ) | ( ~n2363 & n2365 ) | ( n2364 & n2365 ) ;
  assign n2367 = ( x35 & n1447 ) | ( x35 & n1451 ) | ( n1447 & n1451 ) ;
  assign n2368 = x48 & ~x841 ;
  assign n2369 = ( ~x841 & n2367 ) | ( ~x841 & n2368 ) | ( n2367 & n2368 ) ;
  assign n2370 = x47 | n2369 ;
  assign n2371 = n2366 | n2370 ;
  assign n2372 = n1485 & n2371 ;
  assign n2373 = n1652 & n1688 ;
  assign n2374 = n1732 & n2373 ;
  assign n2375 = ~x287 & n1685 ;
  assign n2376 = n1693 & n2375 ;
  assign n2377 = x786 & ~x1082 ;
  assign n2378 = ~n2374 & n2377 ;
  assign n2379 = ( n2374 & n2376 ) | ( n2374 & ~n2378 ) | ( n2376 & ~n2378 ) ;
  assign n2380 = ~n1416 & n2379 ;
  assign n2381 = n2372 | n2380 ;
  assign n2382 = x40 | x102 ;
  assign n2383 = ( ~n1485 & n2342 ) | ( ~n1485 & n2382 ) | ( n2342 & n2382 ) ;
  assign n2384 = n2382 & ~n2383 ;
  assign n2385 = x39 & ~x72 ;
  assign n2386 = ( x41 & x72 ) | ( x41 & ~n2385 ) | ( x72 & ~n2385 ) ;
  assign n2387 = x287 & ~n1701 ;
  assign n2388 = ~n1389 & n2387 ;
  assign n2389 = n2385 & ~n2388 ;
  assign n2390 = ( x152 & n1380 ) | ( x152 & n2235 ) | ( n1380 & n2235 ) ;
  assign n2391 = ~n1380 & n1456 ;
  assign n2392 = n2390 | n2391 ;
  assign n2393 = ~x166 & n2263 ;
  assign n2394 = ~x161 & n2393 ;
  assign n2395 = ~x189 & n2242 ;
  assign n2396 = ~x144 & n2395 ;
  assign n2397 = n2394 | n2396 ;
  assign n2398 = n2393 | n2395 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2400 = ~n2392 & n2399 ;
  assign n2401 = n2386 | n2400 ;
  assign n2402 = ( n2386 & n2389 ) | ( n2386 & n2401 ) | ( n2389 & n2401 ) ;
  assign n2403 = x87 | n1864 ;
  assign n2404 = ( x228 & n1852 ) | ( x228 & n2403 ) | ( n1852 & n2403 ) ;
  assign n2405 = x228 & ~n2404 ;
  assign n2406 = ( n1368 & n2403 ) | ( n1368 & ~n2405 ) | ( n2403 & ~n2405 ) ;
  assign n2407 = x252 & x901 ;
  assign n2408 = ( x94 & x250 ) | ( x94 & x959 ) | ( x250 & x959 ) ;
  assign n2409 = ( x94 & ~n2407 ) | ( x94 & n2408 ) | ( ~n2407 & n2408 ) ;
  assign n2410 = x94 & ~n2409 ;
  assign n2411 = x110 & ~x480 ;
  assign n2412 = x949 & n2411 ;
  assign n2413 = n2410 | n2412 ;
  assign n2414 = x228 | n2413 ;
  assign n2415 = ( n1417 & n2406 ) | ( n1417 & n2414 ) | ( n2406 & n2414 ) ;
  assign n2416 = ~n1417 & n2415 ;
  assign n2417 = ~x44 & n2416 ;
  assign n2418 = ~x101 & n2417 ;
  assign n2419 = ~n2402 & n2418 ;
  assign n2420 = n2402 & ~n2418 ;
  assign n2421 = n2419 | n2420 ;
  assign n2422 = ~x99 & n2419 ;
  assign n2423 = ~x113 & n2422 ;
  assign n2424 = ~n1724 & n2423 ;
  assign n2425 = ~x114 & n2424 ;
  assign n2426 = ~n1421 & n2385 ;
  assign n2427 = n1727 & ~n2388 ;
  assign n2428 = x189 & n2426 ;
  assign n2429 = ( n2426 & ~n2427 ) | ( n2426 & n2428 ) | ( ~n2427 & n2428 ) ;
  assign n2430 = x207 & x208 ;
  assign n2431 = x199 | x200 ;
  assign n2432 = ( x199 & n2430 ) | ( x199 & n2431 ) | ( n2430 & n2431 ) ;
  assign n2433 = n2429 & n2432 ;
  assign n2434 = n1421 & n2385 ;
  assign n2435 = x166 & n2434 ;
  assign n2436 = ( ~n2427 & n2434 ) | ( ~n2427 & n2435 ) | ( n2434 & n2435 ) ;
  assign n2437 = x39 | x72 ;
  assign n2438 = x42 & ~n2437 ;
  assign n2439 = x212 & x214 ;
  assign n2440 = x211 & n2439 ;
  assign n2441 = ( x219 & n2438 ) | ( x219 & ~n2440 ) | ( n2438 & ~n2440 ) ;
  assign n2442 = n2440 | n2441 ;
  assign n2443 = ( n2436 & n2438 ) | ( n2436 & n2442 ) | ( n2438 & n2442 ) ;
  assign n2444 = n2433 | n2443 ;
  assign n2445 = n2425 & ~n2444 ;
  assign n2446 = ~n2425 & n2444 ;
  assign n2447 = n2445 | n2446 ;
  assign n2448 = x43 & ~n2437 ;
  assign n2449 = x200 & ~n2430 ;
  assign n2450 = n2437 & ~n2449 ;
  assign n2451 = ( n2429 & n2448 ) | ( n2429 & ~n2450 ) | ( n2448 & ~n2450 ) ;
  assign n2452 = x211 | x219 ;
  assign n2453 = x212 | x214 ;
  assign n2454 = ~n2439 & n2453 ;
  assign n2455 = ~n2452 & n2454 ;
  assign n2456 = ~x219 & n2453 ;
  assign n2457 = ~n2440 & n2456 ;
  assign n2458 = ~n2455 & n2457 ;
  assign n2459 = ( x211 & ~n2440 ) | ( x211 & n2458 ) | ( ~n2440 & n2458 ) ;
  assign n2460 = n2436 & n2459 ;
  assign n2461 = n2430 & ~n2431 ;
  assign n2462 = n2429 & n2461 ;
  assign n2463 = ( ~n2451 & n2460 ) | ( ~n2451 & n2462 ) | ( n2460 & n2462 ) ;
  assign n2464 = n2451 | n2463 ;
  assign n2465 = n2445 & ~n2464 ;
  assign n2466 = ~n2445 & n2464 ;
  assign n2467 = n2465 | n2466 ;
  assign n2468 = ~n2392 & n2397 ;
  assign n2469 = n2389 & n2468 ;
  assign n2470 = ~x44 & n2469 ;
  assign n2471 = ( x44 & ~n2437 ) | ( x44 & n2469 ) | ( ~n2437 & n2469 ) ;
  assign n2472 = ( ~n2416 & n2470 ) | ( ~n2416 & n2471 ) | ( n2470 & n2471 ) ;
  assign n2473 = ( n2416 & n2470 ) | ( n2416 & n2471 ) | ( n2470 & n2471 ) ;
  assign n2474 = ( n2416 & n2472 ) | ( n2416 & ~n2473 ) | ( n2472 & ~n2473 ) ;
  assign n2475 = x39 & ~x287 ;
  assign n2476 = ~n1416 & n2475 ;
  assign n2477 = x979 & n2476 ;
  assign n2478 = x24 & ~n1482 ;
  assign n2479 = x46 & n2478 ;
  assign n2480 = ~x841 & n2170 ;
  assign n2481 = x61 | n2479 ;
  assign n2482 = ( n2479 & n2480 ) | ( n2479 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2483 = n1484 | n2170 ;
  assign n2484 = x94 & ~n1254 ;
  assign n2485 = ( n1246 & n2350 ) | ( n1246 & n2484 ) | ( n2350 & n2484 ) ;
  assign n2486 = n2484 & ~n2485 ;
  assign n2487 = ( n1319 & ~n1482 ) | ( n1319 & n2486 ) | ( ~n1482 & n2486 ) ;
  assign n2488 = n2483 | n2487 ;
  assign n2489 = x88 | x104 ;
  assign n2490 = ~n1690 & n2489 ;
  assign n2491 = n1470 | n1730 ;
  assign n2492 = x36 & ~n2491 ;
  assign n2493 = n2490 | n2492 ;
  assign n2494 = n1845 & ~n2491 ;
  assign n2495 = n2493 | n2494 ;
  assign n2496 = n2488 & n2495 ;
  assign n2497 = x841 & n2351 ;
  assign n2498 = x48 & n2497 ;
  assign n2499 = x49 & x841 ;
  assign n2500 = ~x24 & x74 ;
  assign n2501 = n2499 | n2500 ;
  assign n2502 = n1825 & n2501 ;
  assign n2503 = x252 & n1470 ;
  assign n2504 = ~x252 & n1729 ;
  assign n2505 = ( n2486 & n2503 ) | ( n2486 & n2504 ) | ( n2503 & n2504 ) ;
  assign n2506 = x24 & x50 ;
  assign n2507 = ( n1306 & n2175 ) | ( n1306 & n2506 ) | ( n2175 & n2506 ) ;
  assign n2508 = n2506 & ~n2507 ;
  assign n2509 = ( ~n1285 & n2505 ) | ( ~n1285 & n2508 ) | ( n2505 & n2508 ) ;
  assign n2510 = n1737 & n2157 ;
  assign n2511 = n2164 & n2165 ;
  assign n2512 = ( ~n2509 & n2510 ) | ( ~n2509 & n2511 ) | ( n2510 & n2511 ) ;
  assign n2513 = n2509 | n2512 ;
  assign n2514 = ( ~n1396 & n2509 ) | ( ~n1396 & n2513 ) | ( n2509 & n2513 ) ;
  assign n2515 = x82 & n2351 ;
  assign n2516 = n2429 & n2430 ;
  assign n2517 = n2439 & ~n2448 ;
  assign n2518 = ( n2436 & n2448 ) | ( n2436 & ~n2517 ) | ( n2448 & ~n2517 ) ;
  assign n2519 = n2429 | n2518 ;
  assign n2520 = n1421 & ~n2452 ;
  assign n2521 = n1421 | n2431 ;
  assign n2522 = ( x39 & n2520 ) | ( x39 & ~n2521 ) | ( n2520 & ~n2521 ) ;
  assign n2523 = ~x39 & x52 ;
  assign n2524 = ( n2519 & n2522 ) | ( n2519 & n2523 ) | ( n2522 & n2523 ) ;
  assign n2525 = ~n2516 & n2524 ;
  assign n2526 = x52 & ~n2437 ;
  assign n2527 = n2445 & n2526 ;
  assign n2528 = ( n2525 & n2526 ) | ( n2525 & ~n2527 ) | ( n2526 & ~n2527 ) ;
  assign n2529 = ( x43 & n2445 ) | ( x43 & ~n2527 ) | ( n2445 & ~n2527 ) ;
  assign n2530 = ( ~x43 & n2528 ) | ( ~x43 & n2529 ) | ( n2528 & n2529 ) ;
  assign n2531 = x53 & ~x60 ;
  assign n2532 = x50 | n2350 ;
  assign n2533 = n1306 | n2532 ;
  assign n2534 = n2531 & ~n2533 ;
  assign n2535 = ( x979 & n1684 ) | ( x979 & ~n2475 ) | ( n1684 & ~n2475 ) ;
  assign n2536 = ( n1684 & n2534 ) | ( n1684 & ~n2535 ) | ( n2534 & ~n2535 ) ;
  assign n2537 = x24 & ~n1383 ;
  assign n2538 = n2536 & n2537 ;
  assign n2539 = ( ~n1416 & n2536 ) | ( ~n1416 & n2538 ) | ( n2536 & n2538 ) ;
  assign n2540 = x106 & n2170 ;
  assign n2541 = ~x841 & n2540 ;
  assign n2542 = x24 & n2337 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = x45 & n2351 ;
  assign n2545 = x24 | n2544 ;
  assign n2546 = ( n1414 & n2544 ) | ( n1414 & n2545 ) | ( n2544 & n2545 ) ;
  assign n2547 = ~x24 & n1414 ;
  assign n2548 = x841 & ~n1404 ;
  assign n2549 = x56 & ~x62 ;
  assign n2550 = n2547 | n2549 ;
  assign n2551 = ( n2547 & n2548 ) | ( n2547 & n2550 ) | ( n2548 & n2550 ) ;
  assign n2552 = x57 & ~n1207 ;
  assign n2553 = x24 & n2552 ;
  assign n2554 = x57 | x841 ;
  assign n2555 = ~x56 & x62 ;
  assign n2556 = ~x924 & n2555 ;
  assign n2557 = ( n2549 & ~n2554 ) | ( n2549 & n2556 ) | ( ~n2554 & n2556 ) ;
  assign n2558 = n2553 | n2557 ;
  assign n2559 = ~n1395 & n2558 ;
  assign n2560 = x90 & ~x841 ;
  assign n2561 = ~n1482 & n2560 ;
  assign n2562 = x924 & ~n2554 ;
  assign n2563 = ( n1395 & ~n2555 ) | ( n1395 & n2562 ) | ( ~n2555 & n2562 ) ;
  assign n2564 = x24 & x59 ;
  assign n2565 = ~n1488 & n2564 ;
  assign n2566 = n2562 | n2565 ;
  assign n2567 = ( ~n2563 & n2565 ) | ( ~n2563 & n2566 ) | ( n2565 & n2566 ) ;
  assign n2568 = n1682 | n1684 ;
  assign n2569 = n2476 & ~n2568 ;
  assign n2570 = x53 | n2533 ;
  assign n2571 = n1416 & ~n2570 ;
  assign n2572 = x24 & n2571 ;
  assign n2573 = n2569 | n2572 ;
  assign n2574 = x61 & n2497 ;
  assign n2575 = x24 & ~n2574 ;
  assign n2576 = ( n2571 & n2574 ) | ( n2571 & ~n2575 ) | ( n2574 & ~n2575 ) ;
  assign n2577 = n2548 & n2555 ;
  assign n2578 = ~x24 & n2552 ;
  assign n2579 = ( ~n1395 & n2577 ) | ( ~n1395 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = x63 & n2351 ;
  assign n2581 = x999 & n2580 ;
  assign n2582 = x24 | n1482 ;
  assign n2583 = x46 & ~n2582 ;
  assign n2584 = n2581 | n2583 ;
  assign n2585 = ( x64 & x107 ) | ( x64 & ~n2358 ) | ( x107 & ~n2358 ) ;
  assign n2586 = n2170 & n2585 ;
  assign n2587 = n2376 & n2377 ;
  assign n2588 = ~n1416 & n2587 ;
  assign n2589 = x314 & ~n2350 ;
  assign n2590 = n1327 & n2589 ;
  assign n2591 = x199 & ~n1421 ;
  assign n2592 = x219 & n1421 ;
  assign n2593 = n2591 | n2592 ;
  assign n2594 = n2590 & n2593 ;
  assign n2595 = x314 & n2351 ;
  assign n2596 = x83 & n2595 ;
  assign n2597 = x39 & ~n1411 ;
  assign n2598 = n1692 & n2597 ;
  assign n2599 = ~n2491 & n2598 ;
  assign n2600 = n1520 & n2599 ;
  assign n2601 = x69 & x314 ;
  assign n2602 = ( x69 & x71 ) | ( x69 & ~n2601 ) | ( x71 & ~n2601 ) ;
  assign n2603 = n2170 & n2602 ;
  assign n2604 = x287 & n2597 ;
  assign n2605 = x70 & n2478 ;
  assign n2606 = n2604 | n2605 ;
  assign n2607 = ~x221 & x299 ;
  assign n2608 = x222 | x299 ;
  assign n2609 = ( n1711 & ~n2607 ) | ( n1711 & n2608 ) | ( ~n2607 & n2608 ) ;
  assign n2610 = n1652 & n1686 ;
  assign n2611 = ~n2609 & n2610 ;
  assign n2612 = n1681 & n1741 ;
  assign n2613 = n2611 & n2612 ;
  assign n2614 = ~n1416 & n2613 ;
  assign n2615 = ( x589 & n1445 ) | ( x589 & n1446 ) | ( n1445 & n1446 ) ;
  assign n2616 = ~x593 & n2615 ;
  assign n2617 = n2614 & n2616 ;
  assign n2618 = n2606 | n2617 ;
  assign n2619 = x211 & ~x219 ;
  assign n2620 = n1421 & ~n2619 ;
  assign n2621 = ~x199 & x200 ;
  assign n2622 = n1421 | n2621 ;
  assign n2623 = ~n2620 & n2622 ;
  assign n2624 = n2590 & n2623 ;
  assign n2625 = ~x85 & n2595 ;
  assign n2626 = ( n2595 & n2624 ) | ( n2595 & ~n2625 ) | ( n2624 & ~n2625 ) ;
  assign n2627 = x24 & n1759 ;
  assign n2628 = x88 & x1093 ;
  assign n2629 = n1690 & n2628 ;
  assign n2630 = ( ~n1318 & n1482 ) | ( ~n1318 & n2629 ) | ( n1482 & n2629 ) ;
  assign n2631 = n2629 & ~n2630 ;
  assign n2632 = ( ~n1482 & n2627 ) | ( ~n1482 & n2631 ) | ( n2627 & n2631 ) ;
  assign n2633 = n1854 | n2632 ;
  assign n2634 = ( n2599 & n2632 ) | ( n2599 & n2633 ) | ( n2632 & n2633 ) ;
  assign n2635 = ~n1743 & n2196 ;
  assign n2636 = x73 & ~n1301 ;
  assign n2637 = ( ~n1362 & n1417 ) | ( ~n1362 & n2636 ) | ( n1417 & n2636 ) ;
  assign n2638 = n2636 & ~n2637 ;
  assign n2639 = n2635 | n2638 ;
  assign n2640 = ~x314 & x1050 ;
  assign n2641 = x39 | n2640 ;
  assign n2642 = n2639 & n2641 ;
  assign n2643 = x24 & x74 ;
  assign n2644 = n1491 & n2643 ;
  assign n2645 = ( x479 & n1445 ) | ( x479 & n1446 ) | ( n1445 & n1446 ) ;
  assign n2646 = x97 & ~n1732 ;
  assign n2647 = ~x479 & n1473 ;
  assign n2648 = ( ~n2645 & n2646 ) | ( ~n2645 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2649 = ~n1470 & n2648 ;
  assign n2650 = n1485 & n2649 ;
  assign n2651 = n2644 | n2650 ;
  assign n2652 = x55 | n1376 ;
  assign n2653 = n1825 & ~n2652 ;
  assign n2654 = ( x75 & n1474 ) | ( x75 & ~n1859 ) | ( n1474 & ~n1859 ) ;
  assign n2655 = n2653 & n2654 ;
  assign n2656 = ( n2172 & ~n2173 ) | ( n2172 & n2326 ) | ( ~n2173 & n2326 ) ;
  assign n2657 = n1729 | n2503 ;
  assign n2658 = n2486 | n2657 ;
  assign n2659 = ( n2171 & ~n2657 ) | ( n2171 & n2658 ) | ( ~n2657 & n2658 ) ;
  assign n2660 = ~n2656 & n2659 ;
  assign n2661 = n1313 & ~n2350 ;
  assign n2662 = x314 & n2661 ;
  assign n2663 = ~x86 & n2662 ;
  assign n2664 = n2661 & ~n2663 ;
  assign n2665 = x232 & n1831 ;
  assign n2666 = x163 | n2302 ;
  assign n2667 = ( x163 & ~n2264 ) | ( x163 & n2302 ) | ( ~n2264 & n2302 ) ;
  assign n2668 = ( n2198 & ~n2666 ) | ( n2198 & n2667 ) | ( ~n2666 & n2667 ) ;
  assign n2669 = n1376 & ~n2254 ;
  assign n2670 = ~x147 & n2669 ;
  assign n2671 = ( ~n2263 & n2669 ) | ( ~n2263 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2672 = ( x184 & n2243 ) | ( x184 & n2307 ) | ( n2243 & n2307 ) ;
  assign n2673 = x184 & n2307 ;
  assign n2674 = ( n2671 & n2672 ) | ( n2671 & ~n2673 ) | ( n2672 & ~n2673 ) ;
  assign n2675 = x187 & n2242 ;
  assign n2676 = n2671 & n2675 ;
  assign n2677 = ( n2668 & ~n2674 ) | ( n2668 & n2676 ) | ( ~n2674 & n2676 ) ;
  assign n2678 = ~n2296 & n2677 ;
  assign n2679 = x153 & x299 ;
  assign n2680 = x175 & ~x299 ;
  assign n2681 = ( n2284 & n2679 ) | ( n2284 & n2680 ) | ( n2679 & n2680 ) ;
  assign n2682 = ( n1431 & n1767 ) | ( n1431 & n1768 ) | ( n1767 & n1768 ) ;
  assign n2683 = n2681 | n2682 ;
  assign n2684 = x166 & x299 ;
  assign n2685 = n1458 | n2684 ;
  assign n2686 = x73 & ~n2685 ;
  assign n2687 = n2683 | n2686 ;
  assign n2688 = x163 & x299 ;
  assign n2689 = x184 & ~x299 ;
  assign n2690 = n2688 | n2689 ;
  assign n2691 = n2201 & n2690 ;
  assign n2692 = n2687 | n2691 ;
  assign n2693 = n1368 & n2692 ;
  assign n2694 = x156 & x299 ;
  assign n2695 = x179 & ~x299 ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = x92 & ~n2696 ;
  assign n2698 = n1727 & ~n2697 ;
  assign n2699 = n1743 | n2685 ;
  assign n2700 = ( n1743 & n2694 ) | ( n1743 & n2695 ) | ( n2694 & n2695 ) ;
  assign n2701 = ( n2277 & ~n2699 ) | ( n2277 & n2700 ) | ( ~n2699 & n2700 ) ;
  assign n2702 = ( x92 & x163 ) | ( x92 & n1369 ) | ( x163 & n1369 ) ;
  assign n2703 = n2698 & n2702 ;
  assign n2704 = ( n2698 & n2701 ) | ( n2698 & n2703 ) | ( n2701 & n2703 ) ;
  assign n2705 = ( n2693 & n2698 ) | ( n2693 & n2704 ) | ( n2698 & n2704 ) ;
  assign n2706 = n2678 | n2705 ;
  assign n2707 = ( ~n1417 & n2678 ) | ( ~n1417 & n2706 ) | ( n2678 & n2706 ) ;
  assign n2708 = n2187 | n2271 ;
  assign n2709 = n2191 & ~n2708 ;
  assign n2710 = ~n2707 & n2709 ;
  assign n2711 = x79 & n2272 ;
  assign n2712 = n2210 | n2711 ;
  assign n2713 = ( ~n2707 & n2710 ) | ( ~n2707 & n2712 ) | ( n2710 & n2712 ) ;
  assign n2714 = ~n1876 & n1879 ;
  assign n2715 = x51 | x87 ;
  assign n2716 = ( n1849 & n2714 ) | ( n1849 & ~n2715 ) | ( n2714 & ~n2715 ) ;
  assign n2717 = ~n1849 & n2716 ;
  assign n2718 = ( ~n2653 & n2714 ) | ( ~n2653 & n2717 ) | ( n2714 & n2717 ) ;
  assign n2719 = x80 | n2144 ;
  assign n2720 = n2142 & ~n2719 ;
  assign n2721 = ~n2718 & n2720 ;
  assign n2722 = x314 | n1238 ;
  assign n2723 = ~x68 & n2722 ;
  assign n2724 = n2170 & ~n2723 ;
  assign n2725 = x66 | n2601 ;
  assign n2726 = n2170 & n2725 ;
  assign n2727 = x83 & ~x314 ;
  assign n2728 = x84 | n2727 ;
  assign n2729 = n2170 & n2728 ;
  assign n2730 = ~n2520 & n2521 ;
  assign n2731 = n2590 & ~n2730 ;
  assign n2732 = x85 & ~x314 ;
  assign n2733 = x67 | n2732 ;
  assign n2734 = n2170 & n2733 ;
  assign n2735 = n1520 & n1715 ;
  assign n2736 = n2597 & n2735 ;
  assign n2737 = x103 & n2595 ;
  assign n2738 = x104 & n1690 ;
  assign n2739 = x88 & n1730 ;
  assign n2740 = n1875 & ~n2739 ;
  assign n2741 = ( n2738 & n2739 ) | ( n2738 & ~n2740 ) | ( n2739 & ~n2740 ) ;
  assign n2742 = n2488 & n2741 ;
  assign n2743 = x70 & ~n2582 ;
  assign n2744 = x89 & n2497 ;
  assign n2745 = n2743 | n2744 ;
  assign n2746 = x73 & ~x1050 ;
  assign n2747 = n2203 | n2746 ;
  assign n2748 = n2488 & n2747 ;
  assign n2749 = x24 | n1714 ;
  assign n2750 = n1714 | n2353 ;
  assign n2751 = ( n2352 & n2353 ) | ( n2352 & n2750 ) | ( n2353 & n2750 ) ;
  assign n2752 = n2749 & n2751 ;
  assign n2753 = ( n2597 & n2749 ) | ( n2597 & n2752 ) | ( n2749 & n2752 ) ;
  assign n2754 = ~n1856 & n2753 ;
  assign n2755 = n1716 | n2640 ;
  assign n2756 = ( n1716 & n1822 ) | ( n1716 & n2755 ) | ( n1822 & n2755 ) ;
  assign n2757 = n1485 & n1696 ;
  assign n2758 = x1050 & ~n2757 ;
  assign n2759 = ( n1822 & n2757 ) | ( n1822 & ~n2758 ) | ( n2757 & ~n2758 ) ;
  assign n2760 = x252 & n1729 ;
  assign n2761 = ( n1470 & ~n2486 ) | ( n1470 & n2760 ) | ( ~n2486 & n2760 ) ;
  assign n2762 = n2760 & ~n2761 ;
  assign n2763 = x49 | n2762 ;
  assign n2764 = ( n2480 & n2762 ) | ( n2480 & n2763 ) | ( n2762 & n2763 ) ;
  assign n2765 = x24 & x95 ;
  assign n2766 = ( x89 & ~x841 ) | ( x89 & n2357 ) | ( ~x841 & n2357 ) ;
  assign n2767 = ( ~n2357 & n2765 ) | ( ~n2357 & n2766 ) | ( n2765 & n2766 ) ;
  assign n2768 = n1485 & n2767 ;
  assign n2769 = ~x287 & n2614 ;
  assign n2770 = n2615 & ~n2768 ;
  assign n2771 = ( n2768 & n2769 ) | ( n2768 & ~n2770 ) | ( n2769 & ~n2770 ) ;
  assign n2772 = ~x24 & x95 ;
  assign n2773 = ~x479 & n1472 ;
  assign n2774 = ( n1470 & n1472 ) | ( n1470 & n2773 ) | ( n1472 & n2773 ) ;
  assign n2775 = ( x96 & n2772 ) | ( x96 & ~n2774 ) | ( n2772 & ~n2774 ) ;
  assign n2776 = n1485 & n2775 ;
  assign n2777 = ~n1470 & n2645 ;
  assign n2778 = x97 & n1732 ;
  assign n2779 = ( x97 & n2777 ) | ( x97 & n2778 ) | ( n2777 & n2778 ) ;
  assign n2780 = ~n1482 & n2779 ;
  assign n2781 = x593 & n2615 ;
  assign n2782 = n2769 & n2781 ;
  assign n2783 = n2780 | n2782 ;
  assign n2784 = x314 & x1050 ;
  assign n2785 = n1822 | n2638 ;
  assign n2786 = n2784 & n2785 ;
  assign n2787 = x99 & ~n2437 ;
  assign n2788 = n2389 & n2392 ;
  assign n2789 = n2399 | n2787 ;
  assign n2790 = ( n2787 & n2788 ) | ( n2787 & n2789 ) | ( n2788 & n2789 ) ;
  assign n2791 = n2419 & ~n2790 ;
  assign n2792 = ~n2419 & n2790 ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = ~n1736 & n2157 ;
  assign n2795 = n1470 & n2151 ;
  assign n2796 = n2794 | n2795 ;
  assign n2797 = ~n2334 & n2796 ;
  assign n2798 = x101 & ~n2437 ;
  assign n2799 = n2397 | n2798 ;
  assign n2800 = ( n2788 & n2798 ) | ( n2788 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = n2417 & ~n2800 ;
  assign n2802 = ~n2417 & n2800 ;
  assign n2803 = n2801 | n2802 ;
  assign n2804 = n1324 & ~n1482 ;
  assign n2805 = x65 & n2804 ;
  assign n2806 = x109 | n1756 ;
  assign n2807 = n2488 & n2806 ;
  assign n2808 = n1875 & n2738 ;
  assign n2809 = n2351 & n2808 ;
  assign n2810 = x110 & ~n1482 ;
  assign n2811 = n1690 & n1729 ;
  assign n2812 = n2810 & ~n2811 ;
  assign n2813 = n2809 | n2812 ;
  assign n2814 = ~x24 & n2534 ;
  assign n2815 = x841 & n2540 ;
  assign n2816 = n2814 | n2815 ;
  assign n2817 = ~x999 & n2580 ;
  assign n2818 = ~x108 & n1850 ;
  assign n2819 = x108 & ~n2366 ;
  assign n2820 = ( n1485 & n2818 ) | ( n1485 & n2819 ) | ( n2818 & n2819 ) ;
  assign n2821 = x87 & ~n1411 ;
  assign n2822 = n2820 | n2821 ;
  assign n2823 = ~x39 & x110 ;
  assign n2824 = n1690 & n1726 ;
  assign n2825 = n2823 & n2824 ;
  assign n2826 = ~n2468 & n2825 ;
  assign n2827 = x111 & n2351 ;
  assign n2828 = x314 & n2827 ;
  assign n2829 = ( ~n1482 & n2826 ) | ( ~n1482 & n2828 ) | ( n2826 & n2828 ) ;
  assign n2830 = ~n1383 & n1759 ;
  assign n2831 = ~x24 & n2830 ;
  assign n2832 = ~x314 & n2827 ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = x124 & ~x468 ;
  assign n2835 = x113 & n2422 ;
  assign n2836 = x113 & ~n2437 ;
  assign n2837 = ~n2422 & n2836 ;
  assign n2838 = ( n2422 & ~n2835 ) | ( n2422 & n2837 ) | ( ~n2835 & n2837 ) ;
  assign n2839 = ( x114 & n2424 ) | ( x114 & n2437 ) | ( n2424 & n2437 ) ;
  assign n2840 = x114 | n2424 ;
  assign n2841 = ~n2839 & n2840 ;
  assign n2842 = x115 & ~n2437 ;
  assign n2843 = ~x116 & n2423 ;
  assign n2844 = n2842 & ~n2843 ;
  assign n2845 = n2424 | n2844 ;
  assign n2846 = x116 & n2423 ;
  assign n2847 = x116 & ~n2437 ;
  assign n2848 = ( n2843 & ~n2846 ) | ( n2843 & n2847 ) | ( ~n2846 & n2847 ) ;
  assign n2849 = x185 & ~n1421 ;
  assign n2850 = x150 & n1421 ;
  assign n2851 = ( n1727 & n2849 ) | ( n1727 & n2850 ) | ( n2849 & n2850 ) ;
  assign n2852 = n1414 & ~n2851 ;
  assign n2853 = n2296 | n2852 ;
  assign n2854 = ( x150 & ~n2264 ) | ( x150 & n2666 ) | ( ~n2264 & n2666 ) ;
  assign n2855 = x150 | n2666 ;
  assign n2856 = ~x185 & n2672 ;
  assign n2857 = x185 & ~n2672 ;
  assign n2858 = ( n2243 & n2856 ) | ( n2243 & n2857 ) | ( n2856 & n2857 ) ;
  assign n2859 = ( ~n2854 & n2855 ) | ( ~n2854 & n2858 ) | ( n2855 & n2858 ) ;
  assign n2860 = ( x143 & n1727 ) | ( x143 & n2263 ) | ( n1727 & n2263 ) ;
  assign n2861 = ~x165 & n2263 ;
  assign n2862 = ( n2669 & ~n2860 ) | ( n2669 & n2861 ) | ( ~n2860 & n2861 ) ;
  assign n2863 = n2859 | n2862 ;
  assign n2864 = x73 & ~x190 ;
  assign n2865 = x185 & ~n2864 ;
  assign n2866 = ( n2201 & n2864 ) | ( n2201 & ~n2865 ) | ( n2864 & ~n2865 ) ;
  assign n2867 = x173 | x299 ;
  assign n2868 = n2284 & ~n2867 ;
  assign n2869 = ( ~x299 & n2866 ) | ( ~x299 & n2868 ) | ( n2866 & n2868 ) ;
  assign n2870 = x73 & ~x168 ;
  assign n2871 = x73 | x150 ;
  assign n2872 = ( n2202 & ~n2870 ) | ( n2202 & n2871 ) | ( ~n2870 & n2871 ) ;
  assign n2873 = ~x151 & n2202 ;
  assign n2874 = ( x299 & ~n2872 ) | ( x299 & n2873 ) | ( ~n2872 & n2873 ) ;
  assign n2875 = n1727 & ~n2874 ;
  assign n2876 = n2205 & n2875 ;
  assign n2877 = ( n2205 & n2869 ) | ( n2205 & ~n2876 ) | ( n2869 & ~n2876 ) ;
  assign n2878 = n2863 | n2877 ;
  assign n2879 = ( n1485 & n2863 ) | ( n1485 & n2878 ) | ( n2863 & n2878 ) ;
  assign n2880 = n2853 | n2879 ;
  assign n2881 = x157 & x299 ;
  assign n2882 = x178 & ~x299 ;
  assign n2883 = ( n1727 & n2881 ) | ( n1727 & n2882 ) | ( n2881 & n2882 ) ;
  assign n2884 = n1716 & ~n2883 ;
  assign n2885 = ( n1822 & ~n2883 ) | ( n1822 & n2884 ) | ( ~n2883 & n2884 ) ;
  assign n2886 = n2880 | n2885 ;
  assign n2887 = ( x118 & n2210 ) | ( x118 & n2709 ) | ( n2210 & n2709 ) ;
  assign n2888 = x118 | n2709 ;
  assign n2889 = ( n2886 & ~n2887 ) | ( n2886 & n2888 ) | ( ~n2887 & n2888 ) ;
  assign n2890 = ( x190 & n1727 ) | ( x190 & n2263 ) | ( n1727 & n2263 ) ;
  assign n2891 = ~x168 & n2263 ;
  assign n2892 = ( n2715 & n2890 ) | ( n2715 & ~n2891 ) | ( n2890 & ~n2891 ) ;
  assign n2893 = n2635 & ~n2892 ;
  assign n2894 = n2889 | n2893 ;
  assign n2895 = n1243 | n1373 ;
  assign n2896 = x91 | x92 ;
  assign n2897 = ( ~x93 & n2895 ) | ( ~x93 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2898 = ( ~x93 & n1775 ) | ( ~x93 & n2897 ) | ( n1775 & n2897 ) ;
  assign n2899 = x93 | n2898 ;
  assign n2900 = x36 | x97 ;
  assign n2901 = n2373 & n2609 ;
  assign n2902 = n2900 | n2901 ;
  assign n2903 = n1714 | n2899 ;
  assign n2904 = ( n2899 & n2902 ) | ( n2899 & n2903 ) | ( n2902 & n2903 ) ;
  assign n2905 = n2653 & n2904 ;
  assign n2906 = x128 & x228 ;
  assign n2907 = ~x128 & x228 ;
  assign n2908 = ( n2905 & n2906 ) | ( n2905 & ~n2907 ) | ( n2906 & ~n2907 ) ;
  assign n2909 = x951 & x982 ;
  assign n2910 = ( ~n1841 & n2144 ) | ( ~n1841 & n2909 ) | ( n2144 & n2909 ) ;
  assign n2911 = x31 | x80 ;
  assign n2912 = x818 & ~n2911 ;
  assign n2913 = n2909 | n2912 ;
  assign n2914 = ( ~n2910 & n2912 ) | ( ~n2910 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = x1093 & n2914 ;
  assign n2916 = x120 | n2915 ;
  assign n2917 = ~n1878 & n2916 ;
  assign n2918 = ~x24 & x77 ;
  assign n2919 = n2661 & ~n2918 ;
  assign n2920 = n1766 & n2662 ;
  assign n2921 = x51 & ~x87 ;
  assign n2922 = ~x146 & n2921 ;
  assign n2923 = ~x87 & x163 ;
  assign n2924 = ( x163 & n2922 ) | ( x163 & ~n2923 ) | ( n2922 & ~n2923 ) ;
  assign n2925 = x67 | x84 ;
  assign n2926 = n1218 | n2925 ;
  assign n2927 = ~n2715 & n2926 ;
  assign n2928 = ~x161 & n2927 ;
  assign n2929 = ( n1421 & n2924 ) | ( n1421 & n2928 ) | ( n2924 & n2928 ) ;
  assign n2930 = n1421 & ~n2929 ;
  assign n2931 = x87 & x184 ;
  assign n2932 = x144 & ~n2931 ;
  assign n2933 = ( n2927 & n2931 ) | ( n2927 & ~n2932 ) | ( n2931 & ~n2932 ) ;
  assign n2934 = ~x142 & n2921 ;
  assign n2935 = ( n1421 & ~n2933 ) | ( n1421 & n2934 ) | ( ~n2933 & n2934 ) ;
  assign n2936 = n2933 | n2935 ;
  assign n2937 = ( n2920 & ~n2930 ) | ( n2920 & n2936 ) | ( ~n2930 & n2936 ) ;
  assign n2938 = ~n2919 & n2937 ;
  assign n2939 = n2696 & n2919 ;
  assign n2940 = ( n1727 & n2938 ) | ( n1727 & n2939 ) | ( n2938 & n2939 ) ;
  assign n2941 = n2715 | n2926 ;
  assign n2942 = x39 | n1382 ;
  assign n2943 = ( n1382 & n1390 ) | ( n1382 & n2942 ) | ( n1390 & n2942 ) ;
  assign n2944 = x24 | x86 ;
  assign n2945 = x314 | n2944 ;
  assign n2946 = ~n1285 & n2945 ;
  assign n2947 = n1313 & n2946 ;
  assign n2948 = n2941 | n2947 ;
  assign n2949 = ( n2941 & ~n2943 ) | ( n2941 & n2948 ) | ( ~n2943 & n2948 ) ;
  assign n2950 = n1708 | n1759 ;
  assign n2951 = ~n2943 & n2950 ;
  assign n2952 = n2949 | n2951 ;
  assign n2953 = x125 | x133 ;
  assign n2954 = ~x121 & n2953 ;
  assign n2955 = x121 | n2953 ;
  assign n2956 = x126 | n2955 ;
  assign n2957 = x132 | n2956 ;
  assign n2958 = x130 | n2957 ;
  assign n2959 = x136 | n2958 ;
  assign n2960 = x135 | n2959 ;
  assign n2961 = x134 | n2960 ;
  assign n2962 = ( ~x121 & n2953 ) | ( ~x121 & n2961 ) | ( n2953 & n2961 ) ;
  assign n2963 = ( n2952 & ~n2954 ) | ( n2952 & n2962 ) | ( ~n2954 & n2962 ) ;
  assign n2964 = ~n2940 & n2963 ;
  assign n2965 = ~x287 & n1727 ;
  assign n2966 = n1773 & n2965 ;
  assign n2967 = n1713 & n2966 ;
  assign n2968 = n2964 & ~n2967 ;
  assign n2969 = ~n1380 & n1707 ;
  assign n2970 = n1681 & n2969 ;
  assign n2971 = ~x215 & x221 ;
  assign n2972 = n1380 & n2971 ;
  assign n2973 = ~n1661 & n1669 ;
  assign n2974 = ( n1662 & n2972 ) | ( n1662 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = x39 & ~x110 ;
  assign n2976 = ( ~n1742 & n1743 ) | ( ~n1742 & n2975 ) | ( n1743 & n2975 ) ;
  assign n2977 = n2975 & ~n2976 ;
  assign n2978 = ( n2970 & n2974 ) | ( n2970 & n2977 ) | ( n2974 & n2977 ) ;
  assign n2979 = n2826 | n2978 ;
  assign n2980 = n2830 | n2979 ;
  assign n2981 = x90 | x111 ;
  assign n2982 = ( n1755 & n2980 ) | ( n1755 & ~n2981 ) | ( n2980 & ~n2981 ) ;
  assign n2983 = n2981 | n2982 ;
  assign n2984 = ( n2488 & n2980 ) | ( n2488 & n2983 ) | ( n2980 & n2983 ) ;
  assign n2985 = x125 & ~x133 ;
  assign n2986 = ~n1762 & n2662 ;
  assign n2987 = x193 | n1421 ;
  assign n2988 = ~x172 & n1421 ;
  assign n2989 = ( n2921 & ~n2987 ) | ( n2921 & n2988 ) | ( ~n2987 & n2988 ) ;
  assign n2990 = ~x162 & n1421 ;
  assign n2991 = x140 | n1421 ;
  assign n2992 = ( x87 & n2990 ) | ( x87 & ~n2991 ) | ( n2990 & ~n2991 ) ;
  assign n2993 = n2989 | n2992 ;
  assign n2994 = n2392 & n2927 ;
  assign n2995 = ~n1727 & n2941 ;
  assign n2996 = ( ~n2993 & n2994 ) | ( ~n2993 & n2995 ) | ( n2994 & n2995 ) ;
  assign n2997 = n2993 | n2996 ;
  assign n2998 = n2919 | n2997 ;
  assign n2999 = n2986 | n2998 ;
  assign n3000 = ~n2952 & n2961 ;
  assign n3001 = ( x125 & ~x133 ) | ( x125 & n3000 ) | ( ~x133 & n3000 ) ;
  assign n3002 = ( ~n2985 & n2999 ) | ( ~n2985 & n3001 ) | ( n2999 & n3001 ) ;
  assign n3003 = n1766 & n2965 ;
  assign n3004 = ~n3002 & n3003 ;
  assign n3005 = ( n1713 & n3002 ) | ( n1713 & ~n3004 ) | ( n3002 & ~n3004 ) ;
  assign n3006 = n2322 & n2919 ;
  assign n3007 = n3005 & ~n3006 ;
  assign n3008 = ( n1243 & ~n2883 ) | ( n1243 & n2918 ) | ( ~n2883 & n2918 ) ;
  assign n3009 = n1727 & n2918 ;
  assign n3010 = n1773 & n3009 ;
  assign n3011 = n3008 & ~n3010 ;
  assign n3012 = n1727 & n1769 ;
  assign n3013 = ~x287 & n3012 ;
  assign n3014 = ( x39 & n1709 ) | ( x39 & n1710 ) | ( n1709 & n1710 ) ;
  assign n3015 = n2941 | n3014 ;
  assign n3016 = ( n2941 & ~n3013 ) | ( n2941 & n3015 ) | ( ~n3013 & n3015 ) ;
  assign n3017 = n3011 | n3016 ;
  assign n3018 = x87 & n2851 ;
  assign n3019 = n3017 & ~n3018 ;
  assign n3020 = n2398 & n2927 ;
  assign n3021 = ~n1380 & n2680 ;
  assign n3022 = ( x153 & n1380 ) | ( x153 & n2679 ) | ( n1380 & n2679 ) ;
  assign n3023 = ( n1727 & n3021 ) | ( n1727 & n3022 ) | ( n3021 & n3022 ) ;
  assign n3024 = n2921 & n3023 ;
  assign n3025 = ( n3019 & n3020 ) | ( n3019 & n3024 ) | ( n3020 & n3024 ) ;
  assign n3026 = n3019 & ~n3025 ;
  assign n3027 = n2952 & n3026 ;
  assign n3028 = x126 & ~n2955 ;
  assign n3029 = ( x126 & ~n2955 ) | ( x126 & n3000 ) | ( ~n2955 & n3000 ) ;
  assign n3030 = ( n3027 & ~n3028 ) | ( n3027 & n3029 ) | ( ~n3028 & n3029 ) ;
  assign n3031 = n1491 | n1698 ;
  assign n3032 = ~x63 & x129 ;
  assign n3033 = x250 & n2760 ;
  assign n3034 = x127 | n3033 ;
  assign n3035 = n1732 & n3033 ;
  assign n3036 = ( n1254 & n3034 ) | ( n1254 & ~n3035 ) | ( n3034 & ~n3035 ) ;
  assign n3037 = ( n1319 & n1324 ) | ( n1319 & n3036 ) | ( n1324 & n3036 ) ;
  assign n3038 = ( ~n1482 & n2483 ) | ( ~n1482 & n3037 ) | ( n2483 & n3037 ) ;
  assign n3039 = n3032 & n3038 ;
  assign n3040 = ( x129 & n3031 ) | ( x129 & n3039 ) | ( n3031 & n3039 ) ;
  assign n3041 = x75 | x250 ;
  assign n3042 = ( x250 & ~n2760 ) | ( x250 & n3041 ) | ( ~n2760 & n3041 ) ;
  assign n3043 = ~x129 & n3042 ;
  assign n3044 = n1732 & ~n3042 ;
  assign n3045 = ( n1373 & n3043 ) | ( n1373 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3046 = n1825 & ~n3045 ;
  assign n3047 = ~n2253 & n2927 ;
  assign n3048 = ( x167 & n1727 ) | ( x167 & n2242 ) | ( n1727 & n2242 ) ;
  assign n3049 = ~x188 & n2242 ;
  assign n3050 = ( x87 & ~n3048 ) | ( x87 & n3049 ) | ( ~n3048 & n3049 ) ;
  assign n3051 = n3047 | n3050 ;
  assign n3052 = ~x130 & n2957 ;
  assign n3053 = ( ~x130 & n2957 ) | ( ~x130 & n3000 ) | ( n2957 & n3000 ) ;
  assign n3054 = ( n3051 & ~n3052 ) | ( n3051 & n3053 ) | ( ~n3052 & n3053 ) ;
  assign n3055 = n2292 & n2965 ;
  assign n3056 = ~n3054 & n3055 ;
  assign n3057 = ( n1713 & n3054 ) | ( n1713 & ~n3056 ) | ( n3054 & ~n3056 ) ;
  assign n3058 = ~x132 & n2956 ;
  assign n3059 = ( ~x132 & n2956 ) | ( ~x132 & n2961 ) | ( n2956 & n2961 ) ;
  assign n3060 = ( n2952 & ~n3058 ) | ( n2952 & n3059 ) | ( ~n3058 & n3059 ) ;
  assign n3061 = n2892 & n2941 ;
  assign n3062 = ( x151 & n1727 ) | ( x151 & n2242 ) | ( n1727 & n2242 ) ;
  assign n3063 = ~x173 & n2242 ;
  assign n3064 = ( n2921 & ~n3062 ) | ( n2921 & n3063 ) | ( ~n3062 & n3063 ) ;
  assign n3065 = n3061 & ~n3064 ;
  assign n3066 = ( ~x232 & n1709 ) | ( ~x232 & n1710 ) | ( n1709 & n1710 ) ;
  assign n3067 = x39 & ~n3066 ;
  assign n3068 = n1759 | n3067 ;
  assign n3069 = n2944 | n3012 ;
  assign n3070 = n2947 & n3069 ;
  assign n3071 = n3068 | n3070 ;
  assign n3072 = x287 | n1661 ;
  assign n3073 = x183 & n1705 ;
  assign n3074 = x149 & n1706 ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = n3072 | n3075 ;
  assign n3077 = ( n1855 & n3072 ) | ( n1855 & ~n3076 ) | ( n3072 & ~n3076 ) ;
  assign n3078 = ~n3065 & n3077 ;
  assign n3079 = ( n2943 & ~n3065 ) | ( n2943 & n3078 ) | ( ~n3065 & n3078 ) ;
  assign n3080 = ( n3065 & n3071 ) | ( n3065 & ~n3079 ) | ( n3071 & ~n3079 ) ;
  assign n3081 = x87 & ~n2259 ;
  assign n3082 = n3080 & ~n3081 ;
  assign n3083 = n3060 & ~n3082 ;
  assign n3084 = x183 & ~n1421 ;
  assign n3085 = x149 & n1421 ;
  assign n3086 = ( n1727 & n3084 ) | ( n1727 & n3085 ) | ( n3084 & n3085 ) ;
  assign n3087 = ( ~x87 & n2921 ) | ( ~x87 & n2926 ) | ( n2921 & n2926 ) ;
  assign n3088 = ( n2941 & ~n3086 ) | ( n2941 & n3087 ) | ( ~n3086 & n3087 ) ;
  assign n3089 = x133 & ~n3088 ;
  assign n3090 = ( n3000 & n3088 ) | ( n3000 & ~n3089 ) | ( n3088 & ~n3089 ) ;
  assign n3091 = ~x287 & n1762 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3093 = ( n1713 & n3090 ) | ( n1713 & ~n3092 ) | ( n3090 & ~n3092 ) ;
  assign n3094 = ~n2247 & n2919 ;
  assign n3095 = n3093 | n3094 ;
  assign n3096 = x134 & n2960 ;
  assign n3097 = ~n2952 & n3096 ;
  assign n3098 = x192 & ~n1421 ;
  assign n3099 = x171 & n1421 ;
  assign n3100 = ( n1727 & n3098 ) | ( n1727 & n3099 ) | ( n3098 & n3099 ) ;
  assign n3101 = n2927 & ~n3100 ;
  assign n3102 = n3097 | n3101 ;
  assign n3103 = ~x287 & n2259 ;
  assign n3104 = ~n3102 & n3103 ;
  assign n3105 = ( n1713 & n3102 ) | ( n1713 & ~n3104 ) | ( n3102 & ~n3104 ) ;
  assign n3106 = x194 & ~n1421 ;
  assign n3107 = x170 & n1421 ;
  assign n3108 = ( n1727 & n3106 ) | ( n1727 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3109 = n2927 | n3108 ;
  assign n3110 = x135 & n2959 ;
  assign n3111 = ( ~n2960 & n3000 ) | ( ~n2960 & n3110 ) | ( n3000 & n3110 ) ;
  assign n3112 = ( ~n3108 & n3109 ) | ( ~n3108 & n3111 ) | ( n3109 & n3111 ) ;
  assign n3113 = ~x287 & n2851 ;
  assign n3114 = ~n3112 & n3113 ;
  assign n3115 = ( n1713 & n3112 ) | ( n1713 & ~n3114 ) | ( n3112 & ~n3114 ) ;
  assign n3116 = x136 & ~n2958 ;
  assign n3117 = ( n1727 & n2312 ) | ( n1727 & n2313 ) | ( n2312 & n2313 ) ;
  assign n3118 = n2927 & ~n3117 ;
  assign n3119 = ( x136 & ~n2958 ) | ( x136 & n3000 ) | ( ~n2958 & n3000 ) ;
  assign n3120 = ( ~n3116 & n3118 ) | ( ~n3116 & n3119 ) | ( n3118 & n3119 ) ;
  assign n3121 = n2690 & n2965 ;
  assign n3122 = ~n3120 & n3121 ;
  assign n3123 = ( n1713 & n3120 ) | ( n1713 & ~n3122 ) | ( n3120 & ~n3122 ) ;
  assign n3124 = ~x39 & x137 ;
  assign n3125 = ~n1380 & n1445 ;
  assign n3126 = ( x210 & n1380 ) | ( x210 & n1446 ) | ( n1380 & n1446 ) ;
  assign n3127 = n3125 | n3126 ;
  assign n3128 = x39 & n2468 ;
  assign n3129 = ~n3127 & n3128 ;
  assign n3130 = ( ~n2604 & n3124 ) | ( ~n2604 & n3129 ) | ( n3124 & n3129 ) ;
  assign n3131 = n2639 & ~n3117 ;
  assign n3132 = n2188 | n2708 ;
  assign n3133 = ( x138 & n2210 ) | ( x138 & ~n3132 ) | ( n2210 & ~n3132 ) ;
  assign n3134 = ( x138 & n2190 ) | ( x138 & ~n3132 ) | ( n2190 & ~n3132 ) ;
  assign n3135 = n3131 | n3134 ;
  assign n3136 = ( n3131 & ~n3133 ) | ( n3131 & n3135 ) | ( ~n3133 & n3135 ) ;
  assign n3137 = ~n2253 & n2639 ;
  assign n3138 = ~x118 & n2709 ;
  assign n3139 = ( x139 & ~n2210 ) | ( x139 & n3138 ) | ( ~n2210 & n3138 ) ;
  assign n3140 = x139 & n3138 ;
  assign n3141 = ( n3137 & n3139 ) | ( n3137 & ~n3140 ) | ( n3139 & ~n3140 ) ;
  assign n3142 = ( n1448 & n1741 ) | ( n1448 & n2629 ) | ( n1741 & n2629 ) ;
  assign n3143 = ( n1741 & n2901 ) | ( n1741 & n3142 ) | ( n2901 & n3142 ) ;
  assign n3144 = x45 | n2382 ;
  assign n3145 = x35 & ~x841 ;
  assign n3146 = ( x47 & ~n2364 ) | ( x47 & n3145 ) | ( ~n2364 & n3145 ) ;
  assign n3147 = n2364 | n3146 ;
  assign n3148 = ( x47 & ~n1732 ) | ( x47 & n3147 ) | ( ~n1732 & n3147 ) ;
  assign n3149 = ( x38 & x120 ) | ( x38 & n1398 ) | ( x120 & n1398 ) ;
  assign n3150 = x252 | n3149 ;
  assign n3151 = ( n3148 & n3149 ) | ( n3148 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3152 = n3144 | n3151 ;
  assign n3153 = ~n1685 & n2475 ;
  assign n3154 = ( ~n3143 & n3152 ) | ( ~n3143 & n3153 ) | ( n3152 & n3153 ) ;
  assign n3155 = n3143 | n3154 ;
  assign n3156 = n1704 & n3155 ;
  assign n3157 = x832 | n3156 ;
  assign n3158 = n1841 & n3157 ;
  assign n3159 = ( x629 & ~x792 ) | ( x629 & x1156 ) | ( ~x792 & x1156 ) ;
  assign n3160 = ( x629 & x792 ) | ( x629 & x1156 ) | ( x792 & x1156 ) ;
  assign n3161 = ~n3159 & n3160 ;
  assign n3162 = ( x618 & x781 ) | ( x618 & x1154 ) | ( x781 & x1154 ) ;
  assign n3163 = x618 & x1154 ;
  assign n3164 = ( n3161 & n3162 ) | ( n3161 & ~n3163 ) | ( n3162 & ~n3163 ) ;
  assign n3165 = ( x608 & ~x778 ) | ( x608 & x1153 ) | ( ~x778 & x1153 ) ;
  assign n3166 = x608 | x1153 ;
  assign n3167 = ( n3164 & ~n3165 ) | ( n3164 & n3166 ) | ( ~n3165 & n3166 ) ;
  assign n3168 = ( x619 & x789 ) | ( x619 & x1159 ) | ( x789 & x1159 ) ;
  assign n3169 = x619 & x1159 ;
  assign n3170 = ( x603 & ~n3168 ) | ( x603 & n3169 ) | ( ~n3168 & n3169 ) ;
  assign n3171 = ( x644 & ~x790 ) | ( x644 & x1160 ) | ( ~x790 & x1160 ) ;
  assign n3172 = ( x644 & x790 ) | ( x644 & x1160 ) | ( x790 & x1160 ) ;
  assign n3173 = ~n3171 & n3172 ;
  assign n3174 = ( x609 & x785 ) | ( x609 & x1155 ) | ( x785 & x1155 ) ;
  assign n3175 = x609 & x1155 ;
  assign n3176 = ( n3173 & n3174 ) | ( n3173 & ~n3175 ) | ( n3174 & ~n3175 ) ;
  assign n3177 = ( x626 & ~x788 ) | ( x626 & x1158 ) | ( ~x788 & x1158 ) ;
  assign n3178 = ( x626 & x788 ) | ( x626 & x1158 ) | ( x788 & x1158 ) ;
  assign n3179 = ~n3177 & n3178 ;
  assign n3180 = ( x630 & x787 ) | ( x630 & x1157 ) | ( x787 & x1157 ) ;
  assign n3181 = x630 & x1157 ;
  assign n3182 = ( n3179 & n3180 ) | ( n3179 & ~n3181 ) | ( n3180 & ~n3181 ) ;
  assign n3183 = n3176 | n3182 ;
  assign n3184 = n3170 & ~n3183 ;
  assign n3185 = ~n3167 & n3184 ;
  assign n3186 = x621 & x1091 ;
  assign n3187 = n3185 & ~n3186 ;
  assign n3188 = n3158 & n3187 ;
  assign n3189 = ~x761 & n3188 ;
  assign n3190 = x140 & ~n3158 ;
  assign n3191 = ( x628 & ~x792 ) | ( x628 & x1156 ) | ( ~x792 & x1156 ) ;
  assign n3192 = ( x628 & x792 ) | ( x628 & x1156 ) | ( x792 & x1156 ) ;
  assign n3193 = ~n3191 & n3192 ;
  assign n3194 = ( x647 & x787 ) | ( x647 & x1157 ) | ( x787 & x1157 ) ;
  assign n3195 = x647 & x1157 ;
  assign n3196 = ( n3193 & n3194 ) | ( n3193 & ~n3195 ) | ( n3194 & ~n3195 ) ;
  assign n3197 = ( x627 & ~x781 ) | ( x627 & x1154 ) | ( ~x781 & x1154 ) ;
  assign n3198 = x627 | x1154 ;
  assign n3199 = ( n3196 & ~n3197 ) | ( n3196 & n3198 ) | ( ~n3197 & n3198 ) ;
  assign n3200 = ( x660 & ~x785 ) | ( x660 & x1155 ) | ( ~x785 & x1155 ) ;
  assign n3201 = x660 | x1155 ;
  assign n3202 = ( x680 & n3200 ) | ( x680 & ~n3201 ) | ( n3200 & ~n3201 ) ;
  assign n3203 = ( x715 & ~x790 ) | ( x715 & x1160 ) | ( ~x790 & x1160 ) ;
  assign n3204 = ( x715 & x790 ) | ( x715 & x1160 ) | ( x790 & x1160 ) ;
  assign n3205 = ~n3203 & n3204 ;
  assign n3206 = ( x625 & x778 ) | ( x625 & x1153 ) | ( x778 & x1153 ) ;
  assign n3207 = x625 & x1153 ;
  assign n3208 = ( n3205 & n3206 ) | ( n3205 & ~n3207 ) | ( n3206 & ~n3207 ) ;
  assign n3209 = ( x641 & ~x788 ) | ( x641 & x1158 ) | ( ~x788 & x1158 ) ;
  assign n3210 = ( x641 & x788 ) | ( x641 & x1158 ) | ( x788 & x1158 ) ;
  assign n3211 = ~n3209 & n3210 ;
  assign n3212 = ( x648 & x789 ) | ( x648 & x1159 ) | ( x789 & x1159 ) ;
  assign n3213 = x648 & x1159 ;
  assign n3214 = ( n3211 & n3212 ) | ( n3211 & ~n3213 ) | ( n3212 & ~n3213 ) ;
  assign n3215 = n3208 | n3214 ;
  assign n3216 = n3202 & ~n3215 ;
  assign n3217 = ~n3199 & n3216 ;
  assign n3218 = x665 & x1091 ;
  assign n3219 = n3217 & ~n3218 ;
  assign n3220 = n1841 & ~n3187 ;
  assign n3221 = n3219 & n3220 ;
  assign n3222 = ~x738 & n3221 ;
  assign n3223 = n3158 & ~n3222 ;
  assign n3224 = ( ~n3189 & n3190 ) | ( ~n3189 & n3223 ) | ( n3190 & n3223 ) ;
  assign n3225 = n3157 & n3221 ;
  assign n3226 = x706 & n3225 ;
  assign n3227 = x141 | n3158 ;
  assign n3228 = ~n3226 & n3227 ;
  assign n3229 = x749 & n3188 ;
  assign n3230 = n3228 & ~n3229 ;
  assign n3231 = x735 & n3225 ;
  assign n3232 = x142 & ~n3158 ;
  assign n3233 = n3231 | n3232 ;
  assign n3234 = x743 & n3188 ;
  assign n3235 = n3233 | n3234 ;
  assign n3236 = x687 & n3225 ;
  assign n3237 = x143 | n3158 ;
  assign n3238 = ~n3236 & n3237 ;
  assign n3239 = ~x774 & n3188 ;
  assign n3240 = n3238 & ~n3239 ;
  assign n3241 = x736 & n3225 ;
  assign n3242 = x144 & ~n3158 ;
  assign n3243 = n3241 | n3242 ;
  assign n3244 = x758 & n3188 ;
  assign n3245 = n3243 | n3244 ;
  assign n3246 = ~x698 & n3225 ;
  assign n3247 = x145 | n3158 ;
  assign n3248 = ~n3246 & n3247 ;
  assign n3249 = ~x767 & n3188 ;
  assign n3250 = n3248 & ~n3249 ;
  assign n3251 = x907 & ~x947 ;
  assign n3252 = n3158 & n3251 ;
  assign n3253 = x735 & n3252 ;
  assign n3254 = x146 | n3158 ;
  assign n3255 = x947 & n3158 ;
  assign n3256 = x743 & n3255 ;
  assign n3257 = n3158 & ~n3256 ;
  assign n3258 = ( n3253 & n3254 ) | ( n3253 & ~n3257 ) | ( n3254 & ~n3257 ) ;
  assign n3259 = ~x770 & n3255 ;
  assign n3260 = x726 & n3252 ;
  assign n3261 = x147 | n3158 ;
  assign n3262 = ~n3260 & n3261 ;
  assign n3263 = ~n3259 & n3262 ;
  assign n3264 = x749 & n3255 ;
  assign n3265 = x706 & n3252 ;
  assign n3266 = x148 | n3158 ;
  assign n3267 = ~n3265 & n3266 ;
  assign n3268 = ~n3264 & n3267 ;
  assign n3269 = ~x755 & n3255 ;
  assign n3270 = ~x725 & n3252 ;
  assign n3271 = x149 | n3158 ;
  assign n3272 = ~n3270 & n3271 ;
  assign n3273 = ~n3269 & n3272 ;
  assign n3274 = ~x751 & n3255 ;
  assign n3275 = ~x701 & n3252 ;
  assign n3276 = x150 | n3158 ;
  assign n3277 = ~n3275 & n3276 ;
  assign n3278 = ~n3274 & n3277 ;
  assign n3279 = ~x745 & n3255 ;
  assign n3280 = ~x723 & n3252 ;
  assign n3281 = x151 | n3158 ;
  assign n3282 = ~n3280 & n3281 ;
  assign n3283 = ~n3279 & n3282 ;
  assign n3284 = x759 & n3255 ;
  assign n3285 = x152 & ~n3158 ;
  assign n3286 = x696 & n3252 ;
  assign n3287 = ( ~n3284 & n3285 ) | ( ~n3284 & n3286 ) | ( n3285 & n3286 ) ;
  assign n3288 = n3284 | n3287 ;
  assign n3289 = x766 & n3255 ;
  assign n3290 = x700 & n3252 ;
  assign n3291 = x153 | n3158 ;
  assign n3292 = ~n3290 & n3291 ;
  assign n3293 = ~n3289 & n3292 ;
  assign n3294 = ~x742 & n3255 ;
  assign n3295 = ~x704 & n3252 ;
  assign n3296 = x154 | n3158 ;
  assign n3297 = ~n3295 & n3296 ;
  assign n3298 = ~n3294 & n3297 ;
  assign n3299 = ~x757 & n3255 ;
  assign n3300 = ~x686 & n3252 ;
  assign n3301 = x155 | n3158 ;
  assign n3302 = ~n3300 & n3301 ;
  assign n3303 = ~n3299 & n3302 ;
  assign n3304 = ~x741 & n3255 ;
  assign n3305 = ~x724 & n3252 ;
  assign n3306 = x156 | n3158 ;
  assign n3307 = ~n3305 & n3306 ;
  assign n3308 = ~n3304 & n3307 ;
  assign n3309 = ~x760 & n3255 ;
  assign n3310 = ~x688 & n3252 ;
  assign n3311 = x157 | n3158 ;
  assign n3312 = ~n3310 & n3311 ;
  assign n3313 = ~n3309 & n3312 ;
  assign n3314 = ~x753 & n3255 ;
  assign n3315 = ~x702 & n3252 ;
  assign n3316 = x158 | n3158 ;
  assign n3317 = ~n3315 & n3316 ;
  assign n3318 = ~n3314 & n3317 ;
  assign n3319 = ~x754 & n3255 ;
  assign n3320 = ~x709 & n3252 ;
  assign n3321 = x159 | n3158 ;
  assign n3322 = ~n3320 & n3321 ;
  assign n3323 = ~n3319 & n3322 ;
  assign n3324 = ~x756 & n3255 ;
  assign n3325 = ~x734 & n3252 ;
  assign n3326 = x160 | n3158 ;
  assign n3327 = ~n3325 & n3326 ;
  assign n3328 = ~n3324 & n3327 ;
  assign n3329 = x758 & n3255 ;
  assign n3330 = x161 & ~n3158 ;
  assign n3331 = x736 & n3252 ;
  assign n3332 = ( ~n3329 & n3330 ) | ( ~n3329 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3333 = n3329 | n3332 ;
  assign n3334 = ~x761 & n3255 ;
  assign n3335 = ~x738 & n3252 ;
  assign n3336 = x162 | n3158 ;
  assign n3337 = ~n3335 & n3336 ;
  assign n3338 = ~n3334 & n3337 ;
  assign n3339 = ~x777 & n3255 ;
  assign n3340 = ~x737 & n3252 ;
  assign n3341 = x163 | n3158 ;
  assign n3342 = ~n3340 & n3341 ;
  assign n3343 = ~n3339 & n3342 ;
  assign n3344 = ~x752 & n3255 ;
  assign n3345 = x703 & n3252 ;
  assign n3346 = x164 | n3158 ;
  assign n3347 = ~n3345 & n3346 ;
  assign n3348 = ~n3344 & n3347 ;
  assign n3349 = ~x774 & n3255 ;
  assign n3350 = x687 & n3252 ;
  assign n3351 = x165 | n3158 ;
  assign n3352 = ~n3350 & n3351 ;
  assign n3353 = ~n3349 & n3352 ;
  assign n3354 = x772 & n3255 ;
  assign n3355 = x166 & ~n3158 ;
  assign n3356 = x727 & n3252 ;
  assign n3357 = ( ~n3354 & n3355 ) | ( ~n3354 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3358 = n3354 | n3357 ;
  assign n3359 = ~x768 & n3255 ;
  assign n3360 = x705 & n3252 ;
  assign n3361 = x167 | n3158 ;
  assign n3362 = ~n3360 & n3361 ;
  assign n3363 = ~n3359 & n3362 ;
  assign n3364 = x763 & n3255 ;
  assign n3365 = x699 & n3252 ;
  assign n3366 = x168 | n3158 ;
  assign n3367 = ~n3365 & n3366 ;
  assign n3368 = ~n3364 & n3367 ;
  assign n3369 = x746 & n3255 ;
  assign n3370 = x729 & n3252 ;
  assign n3371 = x169 | n3158 ;
  assign n3372 = ~n3370 & n3371 ;
  assign n3373 = ~n3369 & n3372 ;
  assign n3374 = x748 & n3255 ;
  assign n3375 = x730 & n3252 ;
  assign n3376 = x170 | n3158 ;
  assign n3377 = ~n3375 & n3376 ;
  assign n3378 = ~n3374 & n3377 ;
  assign n3379 = x764 & n3255 ;
  assign n3380 = x691 & n3252 ;
  assign n3381 = x171 | n3158 ;
  assign n3382 = ~n3380 & n3381 ;
  assign n3383 = ~n3379 & n3382 ;
  assign n3384 = x739 & n3255 ;
  assign n3385 = x690 & n3252 ;
  assign n3386 = x172 | n3158 ;
  assign n3387 = ~n3385 & n3386 ;
  assign n3388 = ~n3384 & n3387 ;
  assign n3389 = ~x723 & n3225 ;
  assign n3390 = x173 | n3158 ;
  assign n3391 = ~n3389 & n3390 ;
  assign n3392 = ~x745 & n3188 ;
  assign n3393 = n3391 & ~n3392 ;
  assign n3394 = x696 & n3225 ;
  assign n3395 = x174 & ~n3158 ;
  assign n3396 = n3394 | n3395 ;
  assign n3397 = x759 & n3188 ;
  assign n3398 = n3396 | n3397 ;
  assign n3399 = x700 & n3225 ;
  assign n3400 = x175 | n3158 ;
  assign n3401 = ~n3399 & n3400 ;
  assign n3402 = x766 & n3188 ;
  assign n3403 = n3401 & ~n3402 ;
  assign n3404 = ~x704 & n3225 ;
  assign n3405 = x176 | n3158 ;
  assign n3406 = ~n3404 & n3405 ;
  assign n3407 = ~x742 & n3188 ;
  assign n3408 = n3406 & ~n3407 ;
  assign n3409 = ~x686 & n3225 ;
  assign n3410 = x177 | n3158 ;
  assign n3411 = ~n3409 & n3410 ;
  assign n3412 = ~x757 & n3188 ;
  assign n3413 = n3411 & ~n3412 ;
  assign n3414 = ~x688 & n3225 ;
  assign n3415 = x178 | n3158 ;
  assign n3416 = ~n3414 & n3415 ;
  assign n3417 = ~x760 & n3188 ;
  assign n3418 = n3416 & ~n3417 ;
  assign n3419 = ~x724 & n3225 ;
  assign n3420 = x179 | n3158 ;
  assign n3421 = ~n3419 & n3420 ;
  assign n3422 = ~x741 & n3188 ;
  assign n3423 = n3421 & ~n3422 ;
  assign n3424 = ~x702 & n3225 ;
  assign n3425 = x180 | n3158 ;
  assign n3426 = ~n3424 & n3425 ;
  assign n3427 = ~x753 & n3188 ;
  assign n3428 = n3426 & ~n3427 ;
  assign n3429 = ~x709 & n3225 ;
  assign n3430 = x181 | n3158 ;
  assign n3431 = ~n3429 & n3430 ;
  assign n3432 = ~x754 & n3188 ;
  assign n3433 = n3431 & ~n3432 ;
  assign n3434 = ~x734 & n3225 ;
  assign n3435 = x182 | n3158 ;
  assign n3436 = ~n3434 & n3435 ;
  assign n3437 = ~x756 & n3188 ;
  assign n3438 = n3436 & ~n3437 ;
  assign n3439 = ~x725 & n3225 ;
  assign n3440 = x183 | n3158 ;
  assign n3441 = ~n3439 & n3440 ;
  assign n3442 = ~x755 & n3188 ;
  assign n3443 = n3441 & ~n3442 ;
  assign n3444 = ~x737 & n3225 ;
  assign n3445 = x184 | n3158 ;
  assign n3446 = ~n3444 & n3445 ;
  assign n3447 = ~x777 & n3188 ;
  assign n3448 = n3446 & ~n3447 ;
  assign n3449 = ~x701 & n3225 ;
  assign n3450 = x185 | n3158 ;
  assign n3451 = ~n3449 & n3450 ;
  assign n3452 = ~x751 & n3188 ;
  assign n3453 = n3451 & ~n3452 ;
  assign n3454 = x703 & n3225 ;
  assign n3455 = x186 | n3158 ;
  assign n3456 = ~n3454 & n3455 ;
  assign n3457 = ~x752 & n3188 ;
  assign n3458 = n3456 & ~n3457 ;
  assign n3459 = x726 & n3225 ;
  assign n3460 = x187 | n3158 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3462 = ~x770 & n3188 ;
  assign n3463 = n3461 & ~n3462 ;
  assign n3464 = x705 & n3225 ;
  assign n3465 = x188 | n3158 ;
  assign n3466 = ~n3464 & n3465 ;
  assign n3467 = ~x768 & n3188 ;
  assign n3468 = n3466 & ~n3467 ;
  assign n3469 = x727 & n3225 ;
  assign n3470 = x189 & ~n3158 ;
  assign n3471 = n3469 | n3470 ;
  assign n3472 = x772 & n3188 ;
  assign n3473 = n3471 | n3472 ;
  assign n3474 = x699 & n3225 ;
  assign n3475 = x190 | n3158 ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = x763 & n3188 ;
  assign n3478 = n3476 & ~n3477 ;
  assign n3479 = x729 & n3225 ;
  assign n3480 = x191 | n3158 ;
  assign n3481 = ~n3479 & n3480 ;
  assign n3482 = x746 & n3188 ;
  assign n3483 = n3481 & ~n3482 ;
  assign n3484 = x691 & n3225 ;
  assign n3485 = x192 | n3158 ;
  assign n3486 = ~n3484 & n3485 ;
  assign n3487 = x764 & n3188 ;
  assign n3488 = n3486 & ~n3487 ;
  assign n3489 = x690 & n3225 ;
  assign n3490 = x193 | n3158 ;
  assign n3491 = ~n3489 & n3490 ;
  assign n3492 = x739 & n3188 ;
  assign n3493 = n3491 & ~n3492 ;
  assign n3494 = x730 & n3225 ;
  assign n3495 = x194 | n3158 ;
  assign n3496 = ~n3494 & n3495 ;
  assign n3497 = x748 & n3188 ;
  assign n3498 = n3496 & ~n3497 ;
  assign n3499 = n2639 & ~n3100 ;
  assign n3500 = x138 | n3132 ;
  assign n3501 = x196 | n3500 ;
  assign n3502 = ~n2210 & n3501 ;
  assign n3503 = x195 | n3499 ;
  assign n3504 = ( n3499 & n3502 ) | ( n3499 & n3503 ) | ( n3502 & n3503 ) ;
  assign n3505 = n2639 & ~n3108 ;
  assign n3506 = x196 & n3500 ;
  assign n3507 = ( n2189 & ~n3501 ) | ( n2189 & n3506 ) | ( ~n3501 & n3506 ) ;
  assign n3508 = ~n2210 & n3507 ;
  assign n3509 = n3505 | n3508 ;
  assign n3510 = ~x767 & n3255 ;
  assign n3511 = ~x698 & n3252 ;
  assign n3512 = x197 | n3158 ;
  assign n3513 = ~n3511 & n3512 ;
  assign n3514 = ~n3510 & n3513 ;
  assign n3515 = n1841 & n3156 ;
  assign n3516 = n3187 & n3515 ;
  assign n3517 = x633 & n3516 ;
  assign n3518 = n3156 & n3221 ;
  assign n3519 = x634 & n3518 ;
  assign n3520 = x198 | n3515 ;
  assign n3521 = ( ~n3515 & n3519 ) | ( ~n3515 & n3520 ) | ( n3519 & n3520 ) ;
  assign n3522 = n3517 | n3521 ;
  assign n3523 = x637 & n3518 ;
  assign n3524 = x199 & ~n3515 ;
  assign n3525 = n3523 | n3524 ;
  assign n3526 = x617 & n3516 ;
  assign n3527 = n3525 | n3526 ;
  assign n3528 = x643 & n3518 ;
  assign n3529 = x200 & ~n3515 ;
  assign n3530 = n3528 | n3529 ;
  assign n3531 = x606 & n3516 ;
  assign n3532 = n3530 | n3531 ;
  assign n3533 = x96 & n3127 ;
  assign n3534 = n1797 & n3533 ;
  assign n3535 = x233 & x237 ;
  assign n3536 = n3534 & n3535 ;
  assign n3537 = n1325 & n2533 ;
  assign n3538 = ( n1325 & n1414 ) | ( n1325 & ~n3537 ) | ( n1414 & ~n3537 ) ;
  assign n3539 = n2338 | n3538 ;
  assign n3540 = n1797 & n3539 ;
  assign n3541 = x332 | n3540 ;
  assign n3542 = ~x32 & x70 ;
  assign n3543 = ~x70 & n1448 ;
  assign n3544 = n3542 | n3543 ;
  assign n3545 = ( ~n3127 & n3542 ) | ( ~n3127 & n3544 ) | ( n3542 & n3544 ) ;
  assign n3546 = n1797 & n3545 ;
  assign n3547 = n3535 & n3546 ;
  assign n3548 = x201 | n3547 ;
  assign n3549 = ~n3536 & n3548 ;
  assign n3550 = ( ~n3536 & n3541 ) | ( ~n3536 & n3549 ) | ( n3541 & n3549 ) ;
  assign n3551 = ~x233 & x237 ;
  assign n3552 = n3534 & n3551 ;
  assign n3553 = x202 | n3551 ;
  assign n3554 = ( x202 & n3546 ) | ( x202 & n3553 ) | ( n3546 & n3553 ) ;
  assign n3555 = n3541 | n3554 ;
  assign n3556 = ~n3552 & n3555 ;
  assign n3557 = x233 | x237 ;
  assign n3558 = n3534 & ~n3557 ;
  assign n3559 = ~x203 & n3557 ;
  assign n3560 = ( x203 & n3546 ) | ( x203 & ~n3559 ) | ( n3546 & ~n3559 ) ;
  assign n3561 = n3541 | n3560 ;
  assign n3562 = ~n3558 & n3561 ;
  assign n3563 = n1791 & n3533 ;
  assign n3564 = n3535 & n3563 ;
  assign n3565 = x468 & ~n1656 ;
  assign n3566 = x468 & n1656 ;
  assign n3567 = ( n1790 & ~n3565 ) | ( n1790 & n3566 ) | ( ~n3565 & n3566 ) ;
  assign n3568 = x332 | n3567 ;
  assign n3569 = ( x332 & n3539 ) | ( x332 & n3568 ) | ( n3539 & n3568 ) ;
  assign n3570 = n3545 & n3567 ;
  assign n3571 = x204 | n3535 ;
  assign n3572 = ( x204 & n3570 ) | ( x204 & n3571 ) | ( n3570 & n3571 ) ;
  assign n3573 = ~n3564 & n3572 ;
  assign n3574 = ( ~n3564 & n3569 ) | ( ~n3564 & n3573 ) | ( n3569 & n3573 ) ;
  assign n3575 = n3551 & n3563 ;
  assign n3576 = n3551 & n3570 ;
  assign n3577 = n3569 | n3576 ;
  assign n3578 = x205 & ~n3575 ;
  assign n3579 = ( ~n3575 & n3577 ) | ( ~n3575 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = x233 & ~x237 ;
  assign n3581 = n3563 & n3580 ;
  assign n3582 = x206 | n3580 ;
  assign n3583 = ( x206 & n3570 ) | ( x206 & n3582 ) | ( n3570 & n3582 ) ;
  assign n3584 = n3569 | n3583 ;
  assign n3585 = ~n3581 & n3584 ;
  assign n3586 = x710 & n3518 ;
  assign n3587 = x207 | n3515 ;
  assign n3588 = ~n3586 & n3587 ;
  assign n3589 = x623 & n3516 ;
  assign n3590 = n3588 & ~n3589 ;
  assign n3591 = x638 & n3518 ;
  assign n3592 = x208 | n3515 ;
  assign n3593 = ~n3591 & n3592 ;
  assign n3594 = x607 & n3516 ;
  assign n3595 = n3593 & ~n3594 ;
  assign n3596 = x639 & n3518 ;
  assign n3597 = x209 | n3515 ;
  assign n3598 = ~n3596 & n3597 ;
  assign n3599 = x622 & n3516 ;
  assign n3600 = n3598 & ~n3599 ;
  assign n3601 = n3251 & n3515 ;
  assign n3602 = x634 & n3601 ;
  assign n3603 = x210 | n3515 ;
  assign n3604 = x947 & n3515 ;
  assign n3605 = x633 & n3604 ;
  assign n3606 = n3515 & ~n3605 ;
  assign n3607 = ( n3602 & n3603 ) | ( n3602 & ~n3606 ) | ( n3603 & ~n3606 ) ;
  assign n3608 = x606 & n3604 ;
  assign n3609 = x211 & ~n3515 ;
  assign n3610 = x643 & n3601 ;
  assign n3611 = ( ~n3608 & n3609 ) | ( ~n3608 & n3610 ) | ( n3609 & n3610 ) ;
  assign n3612 = n3608 | n3611 ;
  assign n3613 = x607 & n3604 ;
  assign n3614 = x638 & n3601 ;
  assign n3615 = x212 | n3515 ;
  assign n3616 = ~n3614 & n3615 ;
  assign n3617 = ~n3613 & n3616 ;
  assign n3618 = x622 & n3604 ;
  assign n3619 = x639 & n3601 ;
  assign n3620 = x213 | n3515 ;
  assign n3621 = ~n3619 & n3620 ;
  assign n3622 = ~n3618 & n3621 ;
  assign n3623 = x623 & n3604 ;
  assign n3624 = x710 & n3601 ;
  assign n3625 = x214 | n3515 ;
  assign n3626 = ~n3624 & n3625 ;
  assign n3627 = ~n3623 & n3626 ;
  assign n3628 = x642 & n3604 ;
  assign n3629 = x215 & ~n3515 ;
  assign n3630 = x681 & n3601 ;
  assign n3631 = ( ~n3628 & n3629 ) | ( ~n3628 & n3630 ) | ( n3629 & n3630 ) ;
  assign n3632 = n3628 | n3631 ;
  assign n3633 = x614 & n3604 ;
  assign n3634 = x216 & ~n3515 ;
  assign n3635 = x662 & n3601 ;
  assign n3636 = ( ~n3633 & n3634 ) | ( ~n3633 & n3635 ) | ( n3634 & n3635 ) ;
  assign n3637 = n3633 | n3636 ;
  assign n3638 = ~x695 & n3518 ;
  assign n3639 = x217 | n3515 ;
  assign n3640 = ~n3638 & n3639 ;
  assign n3641 = x612 & n3516 ;
  assign n3642 = n3640 & ~n3641 ;
  assign n3643 = ~n3557 & n3563 ;
  assign n3644 = ~n3557 & n3570 ;
  assign n3645 = n3569 | n3644 ;
  assign n3646 = x218 & ~n3643 ;
  assign n3647 = ( ~n3643 & n3645 ) | ( ~n3643 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = x617 & n3604 ;
  assign n3649 = x219 & ~n3515 ;
  assign n3650 = x637 & n3601 ;
  assign n3651 = ( ~n3648 & n3649 ) | ( ~n3648 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = n3648 | n3651 ;
  assign n3653 = n3534 & n3580 ;
  assign n3654 = x220 | n3580 ;
  assign n3655 = ( x220 & n3546 ) | ( x220 & n3654 ) | ( n3546 & n3654 ) ;
  assign n3656 = n3541 | n3655 ;
  assign n3657 = ~n3653 & n3656 ;
  assign n3658 = x616 & n3604 ;
  assign n3659 = x221 & ~n3515 ;
  assign n3660 = x661 & n3601 ;
  assign n3661 = ( ~n3658 & n3659 ) | ( ~n3658 & n3660 ) | ( n3659 & n3660 ) ;
  assign n3662 = n3658 | n3661 ;
  assign n3663 = x661 & n3518 ;
  assign n3664 = x222 & ~n3515 ;
  assign n3665 = n3663 | n3664 ;
  assign n3666 = x616 & n3516 ;
  assign n3667 = n3665 | n3666 ;
  assign n3668 = x681 & n3518 ;
  assign n3669 = x223 & ~n3515 ;
  assign n3670 = n3668 | n3669 ;
  assign n3671 = x642 & n3516 ;
  assign n3672 = n3670 | n3671 ;
  assign n3673 = x662 & n3518 ;
  assign n3674 = x224 & ~n3515 ;
  assign n3675 = n3673 | n3674 ;
  assign n3676 = x614 & n3516 ;
  assign n3677 = n3675 | n3676 ;
  assign n3678 = n1239 | n1431 ;
  assign n3679 = ~n1450 & n2653 ;
  assign n3680 = ~n3678 & n3679 ;
  assign n3681 = x228 & x231 ;
  assign n3682 = x228 & ~x231 ;
  assign n3683 = ( n3680 & n3681 ) | ( n3680 & ~n3682 ) | ( n3681 & ~n3682 ) ;
  assign n3684 = x47 | x91 ;
  assign n3685 = ( n2493 & n2830 ) | ( n2493 & ~n3684 ) | ( n2830 & ~n3684 ) ;
  assign n3686 = n3684 | n3685 ;
  assign n3687 = ( n2488 & n2830 ) | ( n2488 & n3686 ) | ( n2830 & n3686 ) ;
  assign n3688 = n1854 | n3687 ;
  assign n3689 = ( n2599 & n3687 ) | ( n2599 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3690 = ~x39 & x228 ;
  assign n3691 = x96 | x97 ;
  assign n3692 = x1091 & x1093 ;
  assign n3693 = ( n1731 & n3691 ) | ( n1731 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3694 = n3690 | n3693 ;
  assign n3695 = ( n1485 & n3690 ) | ( n1485 & n3694 ) | ( n3690 & n3694 ) ;
  assign n3696 = x1091 | n3695 ;
  assign n3697 = ( n2769 & n3695 ) | ( n2769 & n3696 ) | ( n3695 & n3696 ) ;
  assign n3698 = n2342 | n2588 ;
  assign n3699 = ~n2488 & n3698 ;
  assign n3700 = ( n2488 & n3031 ) | ( n2488 & ~n3699 ) | ( n3031 & ~n3699 ) ;
  assign n3701 = x1143 & n2458 ;
  assign n3702 = x1144 & n2455 ;
  assign n3703 = ~x211 & x219 ;
  assign n3704 = ( x219 & n2457 ) | ( x219 & ~n3703 ) | ( n2457 & ~n3703 ) ;
  assign n3705 = ( n2439 & n2454 ) | ( n2439 & ~n3704 ) | ( n2454 & ~n3704 ) ;
  assign n3706 = ~x1142 & n3705 ;
  assign n3707 = ( n3702 & n3705 ) | ( n3702 & ~n3706 ) | ( n3705 & ~n3706 ) ;
  assign n3708 = n3701 | n3707 ;
  assign n3709 = x230 & n1421 ;
  assign n3710 = x213 & n3709 ;
  assign n3711 = ~n3708 & n3710 ;
  assign n3712 = x207 & ~x208 ;
  assign n3713 = x199 & ~x200 ;
  assign n3714 = x1155 & n3713 ;
  assign n3715 = ~x200 & x1157 ;
  assign n3716 = x200 & x1156 ;
  assign n3717 = ( ~x199 & n3715 ) | ( ~x199 & n3716 ) | ( n3715 & n3716 ) ;
  assign n3718 = n3714 | n3717 ;
  assign n3719 = n3712 & n3718 ;
  assign n3720 = x230 & ~n1421 ;
  assign n3721 = ~x209 & n3720 ;
  assign n3722 = ~x200 & x1156 ;
  assign n3723 = x200 & x1155 ;
  assign n3724 = ( ~x199 & n3722 ) | ( ~x199 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = x1154 & n3713 ;
  assign n3726 = n3724 | n3725 ;
  assign n3727 = n3712 & n3726 ;
  assign n3728 = n3721 & n3727 ;
  assign n3729 = x207 | x208 ;
  assign n3730 = n3726 & n3729 ;
  assign n3731 = ~x207 & n3730 ;
  assign n3732 = ( n3721 & n3728 ) | ( n3721 & ~n3731 ) | ( n3728 & ~n3731 ) ;
  assign n3733 = n3719 & n3732 ;
  assign n3734 = ~x200 & x1155 ;
  assign n3735 = x200 & x1154 ;
  assign n3736 = ( ~x199 & n3734 ) | ( ~x199 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = n2430 & n3736 ;
  assign n3738 = x199 & n2430 ;
  assign n3739 = ~n2430 & n3729 ;
  assign n3740 = ( ~x199 & n2432 ) | ( ~x199 & n3713 ) | ( n2432 & n3713 ) ;
  assign n3741 = ( n2430 & n3739 ) | ( n2430 & n3740 ) | ( n3739 & n3740 ) ;
  assign n3742 = x1153 & n3741 ;
  assign n3743 = n3738 & n3742 ;
  assign n3744 = n3737 | n3743 ;
  assign n3745 = ( n3732 & n3733 ) | ( n3732 & ~n3744 ) | ( n3733 & ~n3744 ) ;
  assign n3746 = ( n3711 & ~n3733 ) | ( n3711 & n3745 ) | ( ~n3733 & n3745 ) ;
  assign n3747 = ~x230 & x233 ;
  assign n3748 = x1142 & n3741 ;
  assign n3749 = ~n2431 & n3739 ;
  assign n3750 = x1144 & n3749 ;
  assign n3751 = ~n2432 & n3729 ;
  assign n3752 = ( x200 & n2461 ) | ( x200 & n3751 ) | ( n2461 & n3751 ) ;
  assign n3753 = x1143 & n3752 ;
  assign n3754 = ( ~n3748 & n3750 ) | ( ~n3748 & n3753 ) | ( n3750 & n3753 ) ;
  assign n3755 = n3748 | n3754 ;
  assign n3756 = x209 & n3720 ;
  assign n3757 = ~n3755 & n3756 ;
  assign n3758 = n3747 | n3757 ;
  assign n3759 = x1155 & n2458 ;
  assign n3760 = x1156 & n2455 ;
  assign n3761 = x1154 & n3705 ;
  assign n3762 = n3760 | n3761 ;
  assign n3763 = n3759 | n3762 ;
  assign n3764 = ( x212 & ~x214 ) | ( x212 & n2456 ) | ( ~x214 & n2456 ) ;
  assign n3765 = n3763 & n3764 ;
  assign n3766 = ~x213 & n3709 ;
  assign n3767 = x1157 & ~n2452 ;
  assign n3768 = x1156 & n2619 ;
  assign n3769 = x1155 & n3703 ;
  assign n3770 = ( ~n3767 & n3768 ) | ( ~n3767 & n3769 ) | ( n3768 & n3769 ) ;
  assign n3771 = n3767 | n3770 ;
  assign n3772 = n2439 & n3703 ;
  assign n3773 = x1153 & n3772 ;
  assign n3774 = ~x212 & x214 ;
  assign n3775 = n3773 | n3774 ;
  assign n3776 = ( n3771 & n3773 ) | ( n3771 & n3775 ) | ( n3773 & n3775 ) ;
  assign n3777 = n3766 & ~n3776 ;
  assign n3778 = n3765 | n3777 ;
  assign n3779 = ( n3758 & ~n3765 ) | ( n3758 & n3778 ) | ( ~n3765 & n3778 ) ;
  assign n3780 = n3746 | n3779 ;
  assign n3781 = n2458 | n3705 ;
  assign n3782 = n3741 | n3752 ;
  assign n3783 = n1421 | n3782 ;
  assign n3784 = ~n1421 & n3782 ;
  assign n3785 = ( n3781 & n3783 ) | ( n3781 & n3784 ) | ( n3783 & n3784 ) ;
  assign n3786 = ~n1421 & n3751 ;
  assign n3787 = n1421 & n2457 ;
  assign n3788 = n3786 | n3787 ;
  assign n3789 = x1152 & ~n3788 ;
  assign n3790 = ( x1153 & n3786 ) | ( x1153 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3791 = ( n3785 & n3789 ) | ( n3785 & n3790 ) | ( n3789 & n3790 ) ;
  assign n3792 = ~n3785 & n3788 ;
  assign n3793 = x1154 & n3792 ;
  assign n3794 = n3791 | n3793 ;
  assign n3795 = ~x230 & x234 ;
  assign n3796 = n3710 | n3756 ;
  assign n3797 = x230 & ~n3796 ;
  assign n3798 = n3795 | n3797 ;
  assign n3799 = ( n3794 & n3795 ) | ( n3794 & n3798 ) | ( n3795 & n3798 ) ;
  assign n3800 = n1421 & n3763 ;
  assign n3801 = n2430 & n3724 ;
  assign n3802 = ~n3737 & n3801 ;
  assign n3803 = ( n3730 & n3737 ) | ( n3730 & ~n3802 ) | ( n3737 & ~n3802 ) ;
  assign n3804 = ~n1421 & n3803 ;
  assign n3805 = ( n3796 & n3800 ) | ( n3796 & n3804 ) | ( n3800 & n3804 ) ;
  assign n3806 = n3799 | n3805 ;
  assign n3807 = ~x230 & x235 ;
  assign n3808 = n3739 | n3801 ;
  assign n3809 = ( n3718 & n3801 ) | ( n3718 & n3808 ) | ( n3801 & n3808 ) ;
  assign n3810 = n3807 | n3809 ;
  assign n3811 = ( n3756 & n3807 ) | ( n3756 & n3810 ) | ( n3807 & n3810 ) ;
  assign n3812 = x1155 & n2439 ;
  assign n3813 = n2619 & n3812 ;
  assign n3814 = n2454 | n3813 ;
  assign n3815 = ( n3771 & n3813 ) | ( n3771 & n3814 ) | ( n3813 & n3814 ) ;
  assign n3816 = x1156 & n2458 ;
  assign n3817 = n3815 | n3816 ;
  assign n3818 = n3710 & n3817 ;
  assign n3819 = x1154 & n2461 ;
  assign n3820 = n3736 & n3739 ;
  assign n3821 = ( n3742 & ~n3819 ) | ( n3742 & n3820 ) | ( ~n3819 & n3820 ) ;
  assign n3822 = n3819 | n3821 ;
  assign n3823 = n3738 & n3822 ;
  assign n3824 = ( n3721 & n3822 ) | ( n3721 & n3823 ) | ( n3822 & n3823 ) ;
  assign n3825 = ( n3818 & ~n3823 ) | ( n3818 & n3824 ) | ( ~n3823 & n3824 ) ;
  assign n3826 = n3766 & ~n3772 ;
  assign n3827 = x1154 & n2458 ;
  assign n3828 = x1155 & n2455 ;
  assign n3829 = x1153 & n3705 ;
  assign n3830 = n3828 | n3829 ;
  assign n3831 = n3827 | n3830 ;
  assign n3832 = n3826 & n3831 ;
  assign n3833 = ( ~n3811 & n3825 ) | ( ~n3811 & n3832 ) | ( n3825 & n3832 ) ;
  assign n3834 = n3811 | n3833 ;
  assign n3835 = x1144 & n2458 ;
  assign n3836 = x1145 & n2455 ;
  assign n3837 = x1143 & n3705 ;
  assign n3838 = n3836 | n3837 ;
  assign n3839 = n3835 | n3838 ;
  assign n3840 = x213 & n3839 ;
  assign n3841 = ~x211 & x1158 ;
  assign n3842 = x211 & x1157 ;
  assign n3843 = ( ~x219 & n3841 ) | ( ~x219 & n3842 ) | ( n3841 & n3842 ) ;
  assign n3844 = x1156 & n3703 ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = n3774 & n3845 ;
  assign n3847 = x212 | n3846 ;
  assign n3848 = ( n3817 & n3846 ) | ( n3817 & n3847 ) | ( n3846 & n3847 ) ;
  assign n3849 = ~x213 & x1154 ;
  assign n3850 = n3772 & n3849 ;
  assign n3851 = ( ~x213 & n3848 ) | ( ~x213 & n3850 ) | ( n3848 & n3850 ) ;
  assign n3852 = ( n3709 & n3840 ) | ( n3709 & n3851 ) | ( n3840 & n3851 ) ;
  assign n3853 = n2430 & n3726 ;
  assign n3854 = ~x199 & x1158 ;
  assign n3855 = x199 & x1156 ;
  assign n3856 = ( ~x200 & n3854 ) | ( ~x200 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = x1157 & n2621 ;
  assign n3858 = n3856 | n3857 ;
  assign n3859 = n3712 & n3858 ;
  assign n3860 = x208 & n3718 ;
  assign n3861 = ( n3739 & n3859 ) | ( n3739 & n3860 ) | ( n3859 & n3860 ) ;
  assign n3862 = ( n3721 & n3853 ) | ( n3721 & n3861 ) | ( n3853 & n3861 ) ;
  assign n3863 = x230 | x237 ;
  assign n3864 = ~n3756 & n3863 ;
  assign n3865 = x1145 & n3749 ;
  assign n3866 = x1143 & n3741 ;
  assign n3867 = x1144 & n3752 ;
  assign n3868 = ( ~n3865 & n3866 ) | ( ~n3865 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = n3865 | n3868 ;
  assign n3870 = n3756 & ~n3869 ;
  assign n3871 = ( ~n3862 & n3864 ) | ( ~n3862 & n3870 ) | ( n3864 & n3870 ) ;
  assign n3872 = ~n3852 & n3871 ;
  assign n3873 = ( x1152 & n3786 ) | ( x1152 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3874 = x1151 & ~n3788 ;
  assign n3875 = ( n3785 & n3873 ) | ( n3785 & n3874 ) | ( n3873 & n3874 ) ;
  assign n3876 = x1153 & n3792 ;
  assign n3877 = n3875 | n3876 ;
  assign n3878 = n3797 & n3877 ;
  assign n3879 = n3720 & n3822 ;
  assign n3880 = ~x230 & x238 ;
  assign n3881 = n3709 | n3880 ;
  assign n3882 = ( n3831 & n3880 ) | ( n3831 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = n3879 | n3882 ;
  assign n3884 = n3797 | n3883 ;
  assign n3885 = ( ~n3797 & n3878 ) | ( ~n3797 & n3884 ) | ( n3878 & n3884 ) ;
  assign n3886 = n3756 & n3859 ;
  assign n3887 = ~x230 & x239 ;
  assign n3888 = n3846 | n3887 ;
  assign n3889 = ( n3710 & n3887 ) | ( n3710 & n3888 ) | ( n3887 & n3888 ) ;
  assign n3890 = ( n3728 & ~n3886 ) | ( n3728 & n3889 ) | ( ~n3886 & n3889 ) ;
  assign n3891 = n3886 | n3890 ;
  assign n3892 = ~x212 & n3766 ;
  assign n3893 = n3763 & n3892 ;
  assign n3894 = n3891 | n3893 ;
  assign n3895 = x1147 & ~n3788 ;
  assign n3896 = ( x1148 & n3786 ) | ( x1148 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3897 = ( n3785 & n3895 ) | ( n3785 & n3896 ) | ( n3895 & n3896 ) ;
  assign n3898 = x1149 & n3792 ;
  assign n3899 = n3897 | n3898 ;
  assign n3900 = n3796 & ~n3899 ;
  assign n3901 = x1147 & n2455 ;
  assign n3902 = x1145 & n3705 ;
  assign n3903 = n3901 | n3902 ;
  assign n3904 = x1146 & n2458 ;
  assign n3905 = n3903 | n3904 ;
  assign n3906 = n3709 & n3905 ;
  assign n3907 = n3796 | n3906 ;
  assign n3908 = x1147 & n3749 ;
  assign n3909 = x1145 & n3741 ;
  assign n3910 = x1146 & n3752 ;
  assign n3911 = ( ~n3908 & n3909 ) | ( ~n3908 & n3910 ) | ( n3909 & n3910 ) ;
  assign n3912 = n3908 | n3911 ;
  assign n3913 = n3721 & n3912 ;
  assign n3914 = ( x230 & x240 ) | ( x230 & n3709 ) | ( x240 & n3709 ) ;
  assign n3915 = ( x240 & n3913 ) | ( x240 & ~n3914 ) | ( n3913 & ~n3914 ) ;
  assign n3916 = ( ~n3900 & n3907 ) | ( ~n3900 & n3915 ) | ( n3907 & n3915 ) ;
  assign n3917 = n3796 & n3877 ;
  assign n3918 = x1149 & ~n3788 ;
  assign n3919 = ( x1150 & n3786 ) | ( x1150 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3920 = ( n3785 & n3918 ) | ( n3785 & n3919 ) | ( n3918 & n3919 ) ;
  assign n3921 = x1151 & n3792 ;
  assign n3922 = n3920 | n3921 ;
  assign n3923 = ~x230 & x241 ;
  assign n3924 = n3797 | n3923 ;
  assign n3925 = ( n3922 & n3923 ) | ( n3922 & n3924 ) | ( n3923 & n3924 ) ;
  assign n3926 = n3917 | n3925 ;
  assign n3927 = x1146 & n3749 ;
  assign n3928 = x1144 & n3741 ;
  assign n3929 = x1145 & n3752 ;
  assign n3930 = ( ~n3927 & n3928 ) | ( ~n3927 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3931 = n3927 | n3930 ;
  assign n3932 = x209 & n3931 ;
  assign n3933 = ~x209 & n3755 ;
  assign n3934 = ( n3720 & n3932 ) | ( n3720 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3935 = ~x213 & n3708 ;
  assign n3936 = x1145 & n2458 ;
  assign n3937 = x1146 & n2455 ;
  assign n3938 = x1144 & n3705 ;
  assign n3939 = n3937 | n3938 ;
  assign n3940 = n3936 | n3939 ;
  assign n3941 = x213 & n3940 ;
  assign n3942 = ( n3709 & n3935 ) | ( n3709 & n3941 ) | ( n3935 & n3941 ) ;
  assign n3943 = ~x230 & x242 ;
  assign n3944 = ( ~n3934 & n3942 ) | ( ~n3934 & n3943 ) | ( n3942 & n3943 ) ;
  assign n3945 = n3934 | n3944 ;
  assign n3946 = x230 | x1091 ;
  assign n3947 = n2623 & n3946 ;
  assign n3948 = x1156 & n3947 ;
  assign n3949 = n1421 & n3703 ;
  assign n3950 = ~n1421 & n3713 ;
  assign n3951 = ( n3946 & n3949 ) | ( n3946 & n3950 ) | ( n3949 & n3950 ) ;
  assign n3952 = x1157 & n3951 ;
  assign n3953 = ~n2730 & n3946 ;
  assign n3954 = x1155 & n3953 ;
  assign n3955 = ( ~n3948 & n3952 ) | ( ~n3948 & n3954 ) | ( n3952 & n3954 ) ;
  assign n3956 = n3948 | n3955 ;
  assign n3957 = x83 | x85 ;
  assign n3958 = x81 | n3957 ;
  assign n3959 = ( ~n2593 & n3957 ) | ( ~n2593 & n3958 ) | ( n3957 & n3958 ) ;
  assign n3960 = x314 & n3959 ;
  assign n3961 = x802 & n3960 ;
  assign n3962 = x276 & n3961 ;
  assign n3963 = x271 & n3962 ;
  assign n3964 = x273 & n3963 ;
  assign n3965 = x283 & n3964 ;
  assign n3966 = x272 & n3965 ;
  assign n3967 = x275 & n3966 ;
  assign n3968 = x268 & n3967 ;
  assign n3969 = x253 & n3968 ;
  assign n3970 = x254 & n3969 ;
  assign n3971 = x267 & n3970 ;
  assign n3972 = ~x263 & n3971 ;
  assign n3973 = ( ~x243 & n3946 ) | ( ~x243 & n3972 ) | ( n3946 & n3972 ) ;
  assign n3974 = x243 & ~n3972 ;
  assign n3975 = ( ~n3956 & n3973 ) | ( ~n3956 & n3974 ) | ( n3973 & n3974 ) ;
  assign n3976 = n3721 & n3869 ;
  assign n3977 = ~x230 & x244 ;
  assign n3978 = ( ~n3906 & n3976 ) | ( ~n3906 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3979 = n3756 & n3912 ;
  assign n3980 = n3906 | n3979 ;
  assign n3981 = n3978 | n3980 ;
  assign n3982 = n3766 & ~n3839 ;
  assign n3983 = n3766 & n3839 ;
  assign n3984 = ( n3981 & ~n3982 ) | ( n3981 & n3983 ) | ( ~n3982 & n3983 ) ;
  assign n3985 = ( x1147 & n3786 ) | ( x1147 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3986 = x1146 & ~n3788 ;
  assign n3987 = ( n3785 & n3985 ) | ( n3785 & n3986 ) | ( n3985 & n3986 ) ;
  assign n3988 = x1148 & n3792 ;
  assign n3989 = n3987 | n3988 ;
  assign n3990 = ~x230 & x245 ;
  assign n3991 = n3796 | n3990 ;
  assign n3992 = ( n3989 & n3990 ) | ( n3989 & n3991 ) | ( n3990 & n3991 ) ;
  assign n3993 = n3766 & n3940 ;
  assign n3994 = n3721 & n3931 ;
  assign n3995 = n3993 | n3994 ;
  assign n3996 = n3992 | n3995 ;
  assign n3997 = ( x1149 & n3786 ) | ( x1149 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3998 = x1148 & ~n3788 ;
  assign n3999 = ( n3785 & n3997 ) | ( n3785 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4000 = x1150 & n3792 ;
  assign n4001 = n3999 | n4000 ;
  assign n4002 = n3796 & ~n4001 ;
  assign n4003 = x230 | x246 ;
  assign n4004 = ~n3797 & n4003 ;
  assign n4005 = ( n3989 & n4003 ) | ( n3989 & n4004 ) | ( n4003 & n4004 ) ;
  assign n4006 = ~n4002 & n4005 ;
  assign n4007 = n3796 & ~n3922 ;
  assign n4008 = n3797 & ~n3899 ;
  assign n4009 = x230 | x247 ;
  assign n4010 = ( n4007 & ~n4008 ) | ( n4007 & n4009 ) | ( ~n4008 & n4009 ) ;
  assign n4011 = ~n4007 & n4010 ;
  assign n4012 = ~x230 & x248 ;
  assign n4013 = n3797 | n4012 ;
  assign n4014 = ( n4001 & n4012 ) | ( n4001 & n4013 ) | ( n4012 & n4013 ) ;
  assign n4015 = ( x1151 & n3786 ) | ( x1151 & n3787 ) | ( n3786 & n3787 ) ;
  assign n4016 = x1150 & ~n3788 ;
  assign n4017 = ( n3785 & n4015 ) | ( n3785 & n4016 ) | ( n4015 & n4016 ) ;
  assign n4018 = x1152 & n3792 ;
  assign n4019 = n4017 | n4018 ;
  assign n4020 = n3796 & n4019 ;
  assign n4021 = n4014 | n4020 ;
  assign n4022 = ~n3794 & n3796 ;
  assign n4023 = n3797 & ~n4019 ;
  assign n4024 = x230 | x249 ;
  assign n4025 = ( n4022 & ~n4023 ) | ( n4022 & n4024 ) | ( ~n4023 & n4024 ) ;
  assign n4026 = ~n4022 & n4025 ;
  assign n4027 = n1373 | n2486 ;
  assign n4028 = ( ~n1416 & n2486 ) | ( ~n1416 & n4027 ) | ( n2486 & n4027 ) ;
  assign n4029 = ~x250 & n4028 ;
  assign n4030 = x897 & ~n2431 ;
  assign n4031 = ~x476 & n2621 ;
  assign n4032 = n4030 | n4031 ;
  assign n4033 = x251 & ~n4032 ;
  assign n4034 = x1053 & n4030 ;
  assign n4035 = x1039 & n4031 ;
  assign n4036 = n4034 | n4035 ;
  assign n4037 = n4033 | n4036 ;
  assign n4038 = x252 & x1092 ;
  assign n4039 = ~x1093 & n4038 ;
  assign n4040 = ( ~n2144 & n4038 ) | ( ~n2144 & n4039 ) | ( n4038 & n4039 ) ;
  assign n4041 = n2598 | n4040 ;
  assign n4042 = x1152 & n3947 ;
  assign n4043 = x1153 & n3951 ;
  assign n4044 = x1151 & n3953 ;
  assign n4045 = n4043 | n4044 ;
  assign n4046 = n4042 | n4045 ;
  assign n4047 = ( x253 & n3946 ) | ( x253 & n3968 ) | ( n3946 & n3968 ) ;
  assign n4048 = x253 | n3968 ;
  assign n4049 = ( n4046 & ~n4047 ) | ( n4046 & n4048 ) | ( ~n4047 & n4048 ) ;
  assign n4050 = x1153 & n3947 ;
  assign n4051 = x1154 & n3951 ;
  assign n4052 = x1152 & n3953 ;
  assign n4053 = n4051 | n4052 ;
  assign n4054 = n4050 | n4053 ;
  assign n4055 = ( x254 & n3946 ) | ( x254 & n3969 ) | ( n3946 & n3969 ) ;
  assign n4056 = x254 | n3969 ;
  assign n4057 = ( n4054 & ~n4055 ) | ( n4054 & n4056 ) | ( ~n4055 & n4056 ) ;
  assign n4058 = x1036 & n4031 ;
  assign n4059 = x1049 & n4030 ;
  assign n4060 = n4058 | n4059 ;
  assign n4061 = x255 & ~n4032 ;
  assign n4062 = n4060 | n4061 ;
  assign n4063 = x1070 & n4031 ;
  assign n4064 = x1048 & n4030 ;
  assign n4065 = n4063 | n4064 ;
  assign n4066 = x256 & ~n4032 ;
  assign n4067 = n4065 | n4066 ;
  assign n4068 = x1065 & n2431 ;
  assign n4069 = x1084 & ~n2431 ;
  assign n4070 = n4068 | n4069 ;
  assign n4071 = x257 & ~n4032 ;
  assign n4072 = x257 | n4032 ;
  assign n4073 = ( n4070 & n4071 ) | ( n4070 & n4072 ) | ( n4071 & n4072 ) ;
  assign n4074 = x1062 & n4031 ;
  assign n4075 = x1072 & n4030 ;
  assign n4076 = n4074 | n4075 ;
  assign n4077 = x258 & ~n4032 ;
  assign n4078 = n4076 | n4077 ;
  assign n4079 = x1069 & n4031 ;
  assign n4080 = x1059 & n4030 ;
  assign n4081 = n4079 | n4080 ;
  assign n4082 = x259 & ~n4032 ;
  assign n4083 = n4081 | n4082 ;
  assign n4084 = x1067 & n4031 ;
  assign n4085 = x1044 & n4030 ;
  assign n4086 = n4084 | n4085 ;
  assign n4087 = x260 & ~n4032 ;
  assign n4088 = n4086 | n4087 ;
  assign n4089 = x1040 & n4031 ;
  assign n4090 = x1037 & n4030 ;
  assign n4091 = n4089 | n4090 ;
  assign n4092 = x261 & ~n4032 ;
  assign n4093 = n4091 | n4092 ;
  assign n4094 = x1142 & n3788 ;
  assign n4095 = ~x123 & x228 ;
  assign n4096 = ~x228 & x1093 ;
  assign n4097 = n4095 | n4096 ;
  assign n4098 = x262 | n4097 ;
  assign n4099 = x262 & ~n4097 ;
  assign n4100 = ( ~n4094 & n4098 ) | ( ~n4094 & n4099 ) | ( n4098 & n4099 ) ;
  assign n4101 = x1155 & n3947 ;
  assign n4102 = x1156 & n3951 ;
  assign n4103 = x1154 & n3953 ;
  assign n4104 = n4102 | n4103 ;
  assign n4105 = n4101 | n4104 ;
  assign n4106 = ( ~x263 & n3946 ) | ( ~x263 & n3971 ) | ( n3946 & n3971 ) ;
  assign n4107 = x263 & ~n3971 ;
  assign n4108 = ( ~n4105 & n4106 ) | ( ~n4105 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = x1142 & n3947 ;
  assign n4110 = n3946 | n3960 ;
  assign n4111 = x264 & ~n4109 ;
  assign n4112 = ( ~n4109 & n4110 ) | ( ~n4109 & n4111 ) | ( n4110 & n4111 ) ;
  assign n4113 = x1143 & n3951 ;
  assign n4114 = x1141 & n3953 ;
  assign n4115 = ~n3946 & n3960 ;
  assign n4116 = x796 | n4114 ;
  assign n4117 = ( n4114 & n4115 ) | ( n4114 & n4116 ) | ( n4115 & n4116 ) ;
  assign n4118 = n4113 | n4117 ;
  assign n4119 = n4112 & ~n4118 ;
  assign n4120 = x1143 & n3947 ;
  assign n4121 = x265 & ~n4120 ;
  assign n4122 = ( n4110 & ~n4120 ) | ( n4110 & n4121 ) | ( ~n4120 & n4121 ) ;
  assign n4123 = x1142 & n3953 ;
  assign n4124 = x1144 & n3951 ;
  assign n4125 = x819 | n4124 ;
  assign n4126 = ( n4115 & n4124 ) | ( n4115 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = ( n4122 & n4123 ) | ( n4122 & n4126 ) | ( n4123 & n4126 ) ;
  assign n4128 = n4122 & ~n4127 ;
  assign n4129 = x1136 & n3951 ;
  assign n4130 = x948 | n4129 ;
  assign n4131 = ( n4115 & n4129 ) | ( n4115 & n4130 ) | ( n4129 & n4130 ) ;
  assign n4132 = x1134 & n3953 ;
  assign n4133 = x1135 & n3947 ;
  assign n4134 = x266 | n4133 ;
  assign n4135 = ( ~n4110 & n4133 ) | ( ~n4110 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4136 = ( ~n4131 & n4132 ) | ( ~n4131 & n4135 ) | ( n4132 & n4135 ) ;
  assign n4137 = n4131 | n4136 ;
  assign n4138 = x1154 & n3947 ;
  assign n4139 = x1155 & n3951 ;
  assign n4140 = x1153 & n3953 ;
  assign n4141 = n4139 | n4140 ;
  assign n4142 = n4138 | n4141 ;
  assign n4143 = ( x267 & n3946 ) | ( x267 & n3970 ) | ( n3946 & n3970 ) ;
  assign n4144 = x267 | n3970 ;
  assign n4145 = ( n4142 & ~n4143 ) | ( n4142 & n4144 ) | ( ~n4143 & n4144 ) ;
  assign n4146 = x1151 & n3947 ;
  assign n4147 = x1152 & n3951 ;
  assign n4148 = x1150 & n3953 ;
  assign n4149 = n4147 | n4148 ;
  assign n4150 = n4146 | n4149 ;
  assign n4151 = ( x268 & n3946 ) | ( x268 & n3967 ) | ( n3946 & n3967 ) ;
  assign n4152 = x268 | n3967 ;
  assign n4153 = ( n4150 & ~n4151 ) | ( n4150 & n4152 ) | ( ~n4151 & n4152 ) ;
  assign n4154 = x1137 & n3947 ;
  assign n4155 = x269 & ~n4154 ;
  assign n4156 = ( n4110 & ~n4154 ) | ( n4110 & n4155 ) | ( ~n4154 & n4155 ) ;
  assign n4157 = x1136 & n3953 ;
  assign n4158 = x1138 & n3951 ;
  assign n4159 = x817 | n4158 ;
  assign n4160 = ( n4115 & n4158 ) | ( n4115 & n4159 ) | ( n4158 & n4159 ) ;
  assign n4161 = ( n4156 & n4157 ) | ( n4156 & n4160 ) | ( n4157 & n4160 ) ;
  assign n4162 = n4156 & ~n4161 ;
  assign n4163 = x1140 & n3947 ;
  assign n4164 = x270 & ~n4163 ;
  assign n4165 = ( n4110 & ~n4163 ) | ( n4110 & n4164 ) | ( ~n4163 & n4164 ) ;
  assign n4166 = x1139 & n3953 ;
  assign n4167 = x1141 & n3951 ;
  assign n4168 = x805 | n4167 ;
  assign n4169 = ( n4115 & n4167 ) | ( n4115 & n4168 ) | ( n4167 & n4168 ) ;
  assign n4170 = ( n4165 & n4166 ) | ( n4165 & n4169 ) | ( n4166 & n4169 ) ;
  assign n4171 = n4165 & ~n4170 ;
  assign n4172 = x1147 & n3951 ;
  assign n4173 = x1145 & n3953 ;
  assign n4174 = n4172 | n4173 ;
  assign n4175 = x1146 & n3947 ;
  assign n4176 = n4174 | n4175 ;
  assign n4177 = ( x271 & n3946 ) | ( x271 & n3962 ) | ( n3946 & n3962 ) ;
  assign n4178 = x271 | n3962 ;
  assign n4179 = ( n4176 & ~n4177 ) | ( n4176 & n4178 ) | ( ~n4177 & n4178 ) ;
  assign n4180 = x1150 & n3951 ;
  assign n4181 = x1148 & n3953 ;
  assign n4182 = n4180 | n4181 ;
  assign n4183 = x1149 & n3947 ;
  assign n4184 = n4182 | n4183 ;
  assign n4185 = ( x272 & n3946 ) | ( x272 & n3965 ) | ( n3946 & n3965 ) ;
  assign n4186 = x272 | n3965 ;
  assign n4187 = ( n4184 & ~n4185 ) | ( n4184 & n4186 ) | ( ~n4185 & n4186 ) ;
  assign n4188 = x1147 & n3947 ;
  assign n4189 = x1146 & n3953 ;
  assign n4190 = x1148 & n3951 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = n4188 | n4191 ;
  assign n4193 = ( x273 & n3946 ) | ( x273 & n3963 ) | ( n3946 & n3963 ) ;
  assign n4194 = x273 | n3963 ;
  assign n4195 = ( n4192 & ~n4193 ) | ( n4192 & n4194 ) | ( ~n4193 & n4194 ) ;
  assign n4196 = x1143 & n3953 ;
  assign n4197 = x659 | n4196 ;
  assign n4198 = ( n4115 & n4196 ) | ( n4115 & n4197 ) | ( n4196 & n4197 ) ;
  assign n4199 = x1144 & n3947 ;
  assign n4200 = x1145 & n3951 ;
  assign n4201 = x274 & ~n4200 ;
  assign n4202 = ( n4110 & ~n4200 ) | ( n4110 & n4201 ) | ( ~n4200 & n4201 ) ;
  assign n4203 = ( n4198 & ~n4199 ) | ( n4198 & n4202 ) | ( ~n4199 & n4202 ) ;
  assign n4204 = ~n4198 & n4203 ;
  assign n4205 = x1150 & n3947 ;
  assign n4206 = x1151 & n3951 ;
  assign n4207 = x1149 & n3953 ;
  assign n4208 = n4206 | n4207 ;
  assign n4209 = n4205 | n4208 ;
  assign n4210 = ( x275 & n3946 ) | ( x275 & n3966 ) | ( n3946 & n3966 ) ;
  assign n4211 = x275 | n3966 ;
  assign n4212 = ( n4209 & ~n4210 ) | ( n4209 & n4211 ) | ( ~n4210 & n4211 ) ;
  assign n4213 = x1145 & n3947 ;
  assign n4214 = x1144 & n3953 ;
  assign n4215 = x1146 & n3951 ;
  assign n4216 = n4214 | n4215 ;
  assign n4217 = n4213 | n4216 ;
  assign n4218 = ( x276 & n3946 ) | ( x276 & n3961 ) | ( n3946 & n3961 ) ;
  assign n4219 = x276 | n3961 ;
  assign n4220 = ( n4217 & ~n4218 ) | ( n4217 & n4219 ) | ( ~n4218 & n4219 ) ;
  assign n4221 = x1141 & n3947 ;
  assign n4222 = x277 & ~n4221 ;
  assign n4223 = ( n4110 & ~n4221 ) | ( n4110 & n4222 ) | ( ~n4221 & n4222 ) ;
  assign n4224 = x1140 & n3953 ;
  assign n4225 = x1142 & n3951 ;
  assign n4226 = x820 | n4225 ;
  assign n4227 = ( n4115 & n4225 ) | ( n4115 & n4226 ) | ( n4225 & n4226 ) ;
  assign n4228 = ( n4223 & n4224 ) | ( n4223 & n4227 ) | ( n4224 & n4227 ) ;
  assign n4229 = n4223 & ~n4228 ;
  assign n4230 = x1132 & n3953 ;
  assign n4231 = x976 | n4230 ;
  assign n4232 = ( n4115 & n4230 ) | ( n4115 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = x1133 & n3947 ;
  assign n4234 = x1134 & n3951 ;
  assign n4235 = x278 | n4234 ;
  assign n4236 = ( ~n4110 & n4234 ) | ( ~n4110 & n4235 ) | ( n4234 & n4235 ) ;
  assign n4237 = ( ~n4232 & n4233 ) | ( ~n4232 & n4236 ) | ( n4233 & n4236 ) ;
  assign n4238 = n4232 | n4237 ;
  assign n4239 = x958 & n4115 ;
  assign n4240 = x1134 & n3947 ;
  assign n4241 = x1133 & n3953 ;
  assign n4242 = x1135 & n3951 ;
  assign n4243 = n4241 | n4242 ;
  assign n4244 = n4240 | n4243 ;
  assign n4245 = x279 & ~n4110 ;
  assign n4246 = ( ~n4239 & n4244 ) | ( ~n4239 & n4245 ) | ( n4244 & n4245 ) ;
  assign n4247 = n4239 | n4246 ;
  assign n4248 = x1136 & n3947 ;
  assign n4249 = x280 & ~n4248 ;
  assign n4250 = ( n4110 & ~n4248 ) | ( n4110 & n4249 ) | ( ~n4248 & n4249 ) ;
  assign n4251 = x1135 & n3953 ;
  assign n4252 = x1137 & n3951 ;
  assign n4253 = x914 | n4252 ;
  assign n4254 = ( n4115 & n4252 ) | ( n4115 & n4253 ) | ( n4252 & n4253 ) ;
  assign n4255 = ( n4250 & n4251 ) | ( n4250 & n4254 ) | ( n4251 & n4254 ) ;
  assign n4256 = n4250 & ~n4255 ;
  assign n4257 = x1137 & n3953 ;
  assign n4258 = x830 | n4257 ;
  assign n4259 = ( n4115 & n4257 ) | ( n4115 & n4258 ) | ( n4257 & n4258 ) ;
  assign n4260 = x1138 & n3947 ;
  assign n4261 = x1139 & n3951 ;
  assign n4262 = x281 & ~n4261 ;
  assign n4263 = ( n4110 & ~n4261 ) | ( n4110 & n4262 ) | ( ~n4261 & n4262 ) ;
  assign n4264 = ( n4259 & ~n4260 ) | ( n4259 & n4263 ) | ( ~n4260 & n4263 ) ;
  assign n4265 = ~n4259 & n4264 ;
  assign n4266 = x1139 & n3947 ;
  assign n4267 = x282 & ~n4266 ;
  assign n4268 = ( n4110 & ~n4266 ) | ( n4110 & n4267 ) | ( ~n4266 & n4267 ) ;
  assign n4269 = x1138 & n3953 ;
  assign n4270 = x1140 & n3951 ;
  assign n4271 = x836 | n4270 ;
  assign n4272 = ( n4115 & n4270 ) | ( n4115 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4273 = ( n4268 & n4269 ) | ( n4268 & n4272 ) | ( n4269 & n4272 ) ;
  assign n4274 = n4268 & ~n4273 ;
  assign n4275 = x1149 & n3951 ;
  assign n4276 = x1147 & n3953 ;
  assign n4277 = n4275 | n4276 ;
  assign n4278 = x1148 & n3947 ;
  assign n4279 = n4277 | n4278 ;
  assign n4280 = ( x283 & n3946 ) | ( x283 & n3964 ) | ( n3946 & n3964 ) ;
  assign n4281 = x283 | n3964 ;
  assign n4282 = ( n4279 & ~n4280 ) | ( n4279 & n4281 ) | ( ~n4280 & n4281 ) ;
  assign n4283 = x1143 & n3792 ;
  assign n4284 = x284 | n4097 ;
  assign n4285 = x284 & ~n4097 ;
  assign n4286 = ( ~n4283 & n4284 ) | ( ~n4283 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = n2413 & n2804 ;
  assign n4288 = x122 | n1873 ;
  assign n4289 = n1872 & ~n4288 ;
  assign n4290 = ~n4287 & n4289 ;
  assign n4291 = x289 | x793 ;
  assign n4292 = x285 & ~n4291 ;
  assign n4293 = ~n4290 & n4292 ;
  assign n4294 = x289 & ~x793 ;
  assign n4295 = ( x288 & n1877 ) | ( x288 & ~n4287 ) | ( n1877 & ~n4287 ) ;
  assign n4296 = x286 & x288 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4298 = ( x285 & ~n4294 ) | ( x285 & n4297 ) | ( ~n4294 & n4297 ) ;
  assign n4299 = x285 | n4297 ;
  assign n4300 = ( n4293 & ~n4298 ) | ( n4293 & n4299 ) | ( ~n4298 & n4299 ) ;
  assign n4301 = n1873 & ~n4296 ;
  assign n4302 = ( x793 & n4295 ) | ( x793 & n4301 ) | ( n4295 & n4301 ) ;
  assign n4303 = ( ~x793 & n4295 ) | ( ~x793 & n4301 ) | ( n4295 & n4301 ) ;
  assign n4304 = ~n4302 & n4303 ;
  assign n4305 = ~x287 & x457 ;
  assign n4306 = x332 | n4305 ;
  assign n4307 = ( ~x288 & n1877 ) | ( ~x288 & n4287 ) | ( n1877 & n4287 ) ;
  assign n4308 = ( ~n1877 & n4295 ) | ( ~n1877 & n4307 ) | ( n4295 & n4307 ) ;
  assign n4309 = ~x793 & n4308 ;
  assign n4310 = n4290 & n4292 ;
  assign n4311 = ~n4290 & n4294 ;
  assign n4312 = n4297 | n4311 ;
  assign n4313 = n4291 & n4297 ;
  assign n4314 = ( n4310 & n4312 ) | ( n4310 & ~n4313 ) | ( n4312 & ~n4313 ) ;
  assign n4315 = x290 & x476 ;
  assign n4316 = ~x476 & x1048 ;
  assign n4317 = n4315 | n4316 ;
  assign n4318 = x291 & x476 ;
  assign n4319 = ~x476 & x1049 ;
  assign n4320 = n4318 | n4319 ;
  assign n4321 = x292 & x476 ;
  assign n4322 = ~x476 & x1084 ;
  assign n4323 = n4321 | n4322 ;
  assign n4324 = x293 & x476 ;
  assign n4325 = ~x476 & x1059 ;
  assign n4326 = n4324 | n4325 ;
  assign n4327 = x294 & x476 ;
  assign n4328 = ~x476 & x1072 ;
  assign n4329 = n4327 | n4328 ;
  assign n4330 = x295 & x476 ;
  assign n4331 = ~x476 & x1053 ;
  assign n4332 = n4330 | n4331 ;
  assign n4333 = x296 & x476 ;
  assign n4334 = ~x476 & x1037 ;
  assign n4335 = n4333 | n4334 ;
  assign n4336 = x297 & x476 ;
  assign n4337 = ~x476 & x1044 ;
  assign n4338 = n4336 | n4337 ;
  assign n4339 = x298 & x478 ;
  assign n4340 = ~x478 & x1044 ;
  assign n4341 = n4339 | n4340 ;
  assign n4342 = n2536 | n2540 ;
  assign n4343 = n2337 | n4342 ;
  assign n4344 = ~n1394 & n2578 ;
  assign n4345 = ~x312 & n4344 ;
  assign n4346 = ( x55 & ~x300 ) | ( x55 & n4345 ) | ( ~x300 & n4345 ) ;
  assign n4347 = ( x55 & x300 ) | ( x55 & ~n4345 ) | ( x300 & ~n4345 ) ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = ~x300 & n4345 ;
  assign n4350 = ( x55 & ~x301 ) | ( x55 & n4349 ) | ( ~x301 & n4349 ) ;
  assign n4351 = ( x55 & x301 ) | ( x55 & ~n4349 ) | ( x301 & ~n4349 ) ;
  assign n4352 = n4350 | n4351 ;
  assign n4353 = n1517 | n1520 ;
  assign n4354 = x237 | n4353 ;
  assign n4355 = x937 & n1502 ;
  assign n4356 = x1148 & ~n1502 ;
  assign n4357 = ( n1517 & n4355 ) | ( n1517 & n4356 ) | ( n4355 & n4356 ) ;
  assign n4358 = x273 & n1520 ;
  assign n4359 = n4357 | n4358 ;
  assign n4360 = n4354 & ~n4359 ;
  assign n4361 = x303 & x478 ;
  assign n4362 = ~x478 & x1049 ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = x304 & x478 ;
  assign n4365 = ~x478 & x1048 ;
  assign n4366 = n4364 | n4365 ;
  assign n4367 = x305 & x478 ;
  assign n4368 = ~x478 & x1084 ;
  assign n4369 = n4367 | n4368 ;
  assign n4370 = x306 & x478 ;
  assign n4371 = ~x478 & x1059 ;
  assign n4372 = n4370 | n4371 ;
  assign n4373 = x307 & x478 ;
  assign n4374 = ~x478 & x1053 ;
  assign n4375 = n4373 | n4374 ;
  assign n4376 = x308 & x478 ;
  assign n4377 = ~x478 & x1037 ;
  assign n4378 = n4376 | n4377 ;
  assign n4379 = x309 & x478 ;
  assign n4380 = ~x478 & x1072 ;
  assign n4381 = n4379 | n4380 ;
  assign n4382 = ~x271 & n1520 ;
  assign n4383 = ~x934 & n1517 ;
  assign n4384 = x233 | n4383 ;
  assign n4385 = ( ~n4353 & n4383 ) | ( ~n4353 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4386 = n4382 | n4385 ;
  assign n4387 = x1147 & n1523 ;
  assign n4388 = ~x1147 & n1523 ;
  assign n4389 = ( n4386 & ~n4387 ) | ( n4386 & n4388 ) | ( ~n4387 & n4388 ) ;
  assign n4390 = x301 & n4349 ;
  assign n4391 = ( x55 & ~x311 ) | ( x55 & n4390 ) | ( ~x311 & n4390 ) ;
  assign n4392 = ( x55 & x311 ) | ( x55 & ~n4390 ) | ( x311 & ~n4390 ) ;
  assign n4393 = n4391 | n4392 ;
  assign n4394 = ( ~x55 & x312 ) | ( ~x55 & n4344 ) | ( x312 & n4344 ) ;
  assign n4395 = x312 & n4344 ;
  assign n4396 = n4394 & ~n4395 ;
  assign n4397 = ~n1732 & n2810 ;
  assign n4398 = x314 & n1732 ;
  assign n4399 = ( n2827 & n4397 ) | ( n2827 & ~n4398 ) | ( n4397 & ~n4398 ) ;
  assign n4400 = ~x313 & x954 ;
  assign n4401 = x313 & x954 ;
  assign n4402 = ( n4399 & n4400 ) | ( n4399 & ~n4401 ) | ( n4400 & ~n4401 ) ;
  assign n4403 = n2949 | n2961 ;
  assign n4404 = n1713 | n4403 ;
  assign n4405 = ~x340 & n4287 ;
  assign n4406 = ~x1080 & n4405 ;
  assign n4407 = x315 | n4405 ;
  assign n4408 = ~n4406 & n4407 ;
  assign n4409 = x316 & ~n4405 ;
  assign n4410 = x1047 & n4405 ;
  assign n4411 = n4409 | n4410 ;
  assign n4412 = ~x330 & n4287 ;
  assign n4413 = ~x1078 & n4412 ;
  assign n4414 = x317 | n4412 ;
  assign n4415 = ~n4413 & n4414 ;
  assign n4416 = ~x341 & n4287 ;
  assign n4417 = ~x1074 & n4416 ;
  assign n4418 = x318 | n4416 ;
  assign n4419 = ~n4417 & n4418 ;
  assign n4420 = x319 & ~n4416 ;
  assign n4421 = x1072 & n4416 ;
  assign n4422 = n4420 | n4421 ;
  assign n4423 = x320 & ~n4405 ;
  assign n4424 = x1048 & n4405 ;
  assign n4425 = n4423 | n4424 ;
  assign n4426 = x321 & ~n4405 ;
  assign n4427 = x1058 & n4405 ;
  assign n4428 = n4426 | n4427 ;
  assign n4429 = x322 & ~n4405 ;
  assign n4430 = x1051 & n4405 ;
  assign n4431 = n4429 | n4430 ;
  assign n4432 = x323 & ~n4405 ;
  assign n4433 = x1065 & n4405 ;
  assign n4434 = n4432 | n4433 ;
  assign n4435 = x324 & ~n4416 ;
  assign n4436 = x1086 & n4416 ;
  assign n4437 = n4435 | n4436 ;
  assign n4438 = x325 & ~n4416 ;
  assign n4439 = x1063 & n4416 ;
  assign n4440 = n4438 | n4439 ;
  assign n4441 = x326 & ~n4416 ;
  assign n4442 = x1057 & n4416 ;
  assign n4443 = n4441 | n4442 ;
  assign n4444 = x327 & ~n4405 ;
  assign n4445 = x1040 & n4405 ;
  assign n4446 = n4444 | n4445 ;
  assign n4447 = x328 & ~n4416 ;
  assign n4448 = x1058 & n4416 ;
  assign n4449 = n4447 | n4448 ;
  assign n4450 = x329 & ~n4416 ;
  assign n4451 = x1043 & n4416 ;
  assign n4452 = n4450 | n4451 ;
  assign n4453 = x1092 & ~n3692 ;
  assign n4454 = x330 | n4287 ;
  assign n4455 = ( n4405 & n4453 ) | ( n4405 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = x331 | n4287 ;
  assign n4457 = ( n4416 & n4453 ) | ( n4416 & ~n4456 ) | ( n4453 & ~n4456 ) ;
  assign n4458 = n1398 & ~n2475 ;
  assign n4459 = ~n1237 & n2357 ;
  assign n4460 = ~n1355 & n4459 ;
  assign n4461 = x46 | n1480 ;
  assign n4462 = n1224 & ~n4461 ;
  assign n4463 = ( n4460 & n4461 ) | ( n4460 & ~n4462 ) | ( n4461 & ~n4462 ) ;
  assign n4464 = ~n1301 & n4463 ;
  assign n4465 = n4458 | n4464 ;
  assign n4466 = ~n1417 & n4465 ;
  assign n4467 = x333 & ~n4416 ;
  assign n4468 = x1040 & n4416 ;
  assign n4469 = n4467 | n4468 ;
  assign n4470 = x334 & ~n4416 ;
  assign n4471 = x1065 & n4416 ;
  assign n4472 = n4470 | n4471 ;
  assign n4473 = x335 & ~n4416 ;
  assign n4474 = x1069 & n4416 ;
  assign n4475 = n4473 | n4474 ;
  assign n4476 = x336 & ~n4412 ;
  assign n4477 = x1070 & n4412 ;
  assign n4478 = n4476 | n4477 ;
  assign n4479 = x337 & ~n4412 ;
  assign n4480 = x1044 & n4412 ;
  assign n4481 = n4479 | n4480 ;
  assign n4482 = x338 & ~n4412 ;
  assign n4483 = x1072 & n4412 ;
  assign n4484 = n4482 | n4483 ;
  assign n4485 = x339 & ~n4412 ;
  assign n4486 = x1086 & n4412 ;
  assign n4487 = n4485 | n4486 ;
  assign n4488 = x331 & n4287 ;
  assign n4489 = x340 & ~n4287 ;
  assign n4490 = ( n4453 & n4488 ) | ( n4453 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = x341 | n4287 ;
  assign n4492 = ( n4412 & n4453 ) | ( n4412 & ~n4491 ) | ( n4453 & ~n4491 ) ;
  assign n4493 = x342 & ~n4405 ;
  assign n4494 = x1049 & n4405 ;
  assign n4495 = n4493 | n4494 ;
  assign n4496 = x343 & ~n4405 ;
  assign n4497 = x1062 & n4405 ;
  assign n4498 = n4496 | n4497 ;
  assign n4499 = x344 & ~n4405 ;
  assign n4500 = x1069 & n4405 ;
  assign n4501 = n4499 | n4500 ;
  assign n4502 = x345 & ~n4405 ;
  assign n4503 = x1039 & n4405 ;
  assign n4504 = n4502 | n4503 ;
  assign n4505 = x346 & ~n4405 ;
  assign n4506 = x1067 & n4405 ;
  assign n4507 = n4505 | n4506 ;
  assign n4508 = x347 & ~n4405 ;
  assign n4509 = x1055 & n4405 ;
  assign n4510 = n4508 | n4509 ;
  assign n4511 = x348 & ~n4405 ;
  assign n4512 = x1087 & n4405 ;
  assign n4513 = n4511 | n4512 ;
  assign n4514 = x349 & ~n4405 ;
  assign n4515 = x1043 & n4405 ;
  assign n4516 = n4514 | n4515 ;
  assign n4517 = x350 & ~n4405 ;
  assign n4518 = x1035 & n4405 ;
  assign n4519 = n4517 | n4518 ;
  assign n4520 = x351 & ~n4405 ;
  assign n4521 = x1079 & n4405 ;
  assign n4522 = n4520 | n4521 ;
  assign n4523 = x352 & ~n4405 ;
  assign n4524 = x1078 & n4405 ;
  assign n4525 = n4523 | n4524 ;
  assign n4526 = x353 & ~n4405 ;
  assign n4527 = x1063 & n4405 ;
  assign n4528 = n4526 | n4527 ;
  assign n4529 = x354 & ~n4405 ;
  assign n4530 = x1045 & n4405 ;
  assign n4531 = n4529 | n4530 ;
  assign n4532 = x355 & ~n4405 ;
  assign n4533 = x1084 & n4405 ;
  assign n4534 = n4532 | n4533 ;
  assign n4535 = x356 & ~n4405 ;
  assign n4536 = x1081 & n4405 ;
  assign n4537 = n4535 | n4536 ;
  assign n4538 = x357 & ~n4405 ;
  assign n4539 = x1076 & n4405 ;
  assign n4540 = n4538 | n4539 ;
  assign n4541 = x358 & ~n4405 ;
  assign n4542 = x1071 & n4405 ;
  assign n4543 = n4541 | n4542 ;
  assign n4544 = x359 & ~n4405 ;
  assign n4545 = x1068 & n4405 ;
  assign n4546 = n4544 | n4545 ;
  assign n4547 = x360 & ~n4405 ;
  assign n4548 = x1042 & n4405 ;
  assign n4549 = n4547 | n4548 ;
  assign n4550 = x361 & ~n4405 ;
  assign n4551 = x1059 & n4405 ;
  assign n4552 = n4550 | n4551 ;
  assign n4553 = x362 & ~n4405 ;
  assign n4554 = x1070 & n4405 ;
  assign n4555 = n4553 | n4554 ;
  assign n4556 = x363 & ~n4412 ;
  assign n4557 = x1049 & n4412 ;
  assign n4558 = n4556 | n4557 ;
  assign n4559 = x364 & ~n4412 ;
  assign n4560 = x1062 & n4412 ;
  assign n4561 = n4559 | n4560 ;
  assign n4562 = x365 & ~n4412 ;
  assign n4563 = x1065 & n4412 ;
  assign n4564 = n4562 | n4563 ;
  assign n4565 = x366 & ~n4412 ;
  assign n4566 = x1069 & n4412 ;
  assign n4567 = n4565 | n4566 ;
  assign n4568 = x367 & ~n4412 ;
  assign n4569 = x1039 & n4412 ;
  assign n4570 = n4568 | n4569 ;
  assign n4571 = x368 & ~n4412 ;
  assign n4572 = x1067 & n4412 ;
  assign n4573 = n4571 | n4572 ;
  assign n4574 = x369 & ~n4412 ;
  assign n4575 = x1080 & n4412 ;
  assign n4576 = n4574 | n4575 ;
  assign n4577 = x370 & ~n4412 ;
  assign n4578 = x1055 & n4412 ;
  assign n4579 = n4577 | n4578 ;
  assign n4580 = x371 & ~n4412 ;
  assign n4581 = x1051 & n4412 ;
  assign n4582 = n4580 | n4581 ;
  assign n4583 = x372 & ~n4412 ;
  assign n4584 = x1048 & n4412 ;
  assign n4585 = n4583 | n4584 ;
  assign n4586 = x373 & ~n4412 ;
  assign n4587 = x1087 & n4412 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = x374 & ~n4412 ;
  assign n4590 = x1035 & n4412 ;
  assign n4591 = n4589 | n4590 ;
  assign n4592 = x375 & ~n4412 ;
  assign n4593 = x1047 & n4412 ;
  assign n4594 = n4592 | n4593 ;
  assign n4595 = x376 & ~n4412 ;
  assign n4596 = x1079 & n4412 ;
  assign n4597 = n4595 | n4596 ;
  assign n4598 = x377 & ~n4412 ;
  assign n4599 = x1074 & n4412 ;
  assign n4600 = n4598 | n4599 ;
  assign n4601 = x378 & ~n4412 ;
  assign n4602 = x1063 & n4412 ;
  assign n4603 = n4601 | n4602 ;
  assign n4604 = x379 & ~n4412 ;
  assign n4605 = x1045 & n4412 ;
  assign n4606 = n4604 | n4605 ;
  assign n4607 = x380 & ~n4412 ;
  assign n4608 = x1084 & n4412 ;
  assign n4609 = n4607 | n4608 ;
  assign n4610 = x381 & ~n4412 ;
  assign n4611 = x1081 & n4412 ;
  assign n4612 = n4610 | n4611 ;
  assign n4613 = x382 & ~n4412 ;
  assign n4614 = x1076 & n4412 ;
  assign n4615 = n4613 | n4614 ;
  assign n4616 = x383 & ~n4412 ;
  assign n4617 = x1071 & n4412 ;
  assign n4618 = n4616 | n4617 ;
  assign n4619 = x384 & ~n4412 ;
  assign n4620 = x1068 & n4412 ;
  assign n4621 = n4619 | n4620 ;
  assign n4622 = x385 & ~n4412 ;
  assign n4623 = x1042 & n4412 ;
  assign n4624 = n4622 | n4623 ;
  assign n4625 = x386 & ~n4412 ;
  assign n4626 = x1059 & n4412 ;
  assign n4627 = n4625 | n4626 ;
  assign n4628 = x387 & ~n4412 ;
  assign n4629 = x1053 & n4412 ;
  assign n4630 = n4628 | n4629 ;
  assign n4631 = x388 & ~n4412 ;
  assign n4632 = x1037 & n4412 ;
  assign n4633 = n4631 | n4632 ;
  assign n4634 = x389 & ~n4412 ;
  assign n4635 = x1036 & n4412 ;
  assign n4636 = n4634 | n4635 ;
  assign n4637 = x390 & ~n4416 ;
  assign n4638 = x1049 & n4416 ;
  assign n4639 = n4637 | n4638 ;
  assign n4640 = x391 & ~n4416 ;
  assign n4641 = x1062 & n4416 ;
  assign n4642 = n4640 | n4641 ;
  assign n4643 = x392 & ~n4416 ;
  assign n4644 = x1039 & n4416 ;
  assign n4645 = n4643 | n4644 ;
  assign n4646 = x393 & ~n4416 ;
  assign n4647 = x1067 & n4416 ;
  assign n4648 = n4646 | n4647 ;
  assign n4649 = x394 & ~n4416 ;
  assign n4650 = x1080 & n4416 ;
  assign n4651 = n4649 | n4650 ;
  assign n4652 = x395 & ~n4416 ;
  assign n4653 = x1055 & n4416 ;
  assign n4654 = n4652 | n4653 ;
  assign n4655 = x396 & ~n4416 ;
  assign n4656 = x1051 & n4416 ;
  assign n4657 = n4655 | n4656 ;
  assign n4658 = x397 & ~n4416 ;
  assign n4659 = x1048 & n4416 ;
  assign n4660 = n4658 | n4659 ;
  assign n4661 = x398 & ~n4416 ;
  assign n4662 = x1087 & n4416 ;
  assign n4663 = n4661 | n4662 ;
  assign n4664 = x399 & ~n4416 ;
  assign n4665 = x1047 & n4416 ;
  assign n4666 = n4664 | n4665 ;
  assign n4667 = x400 & ~n4416 ;
  assign n4668 = x1035 & n4416 ;
  assign n4669 = n4667 | n4668 ;
  assign n4670 = x401 & ~n4416 ;
  assign n4671 = x1079 & n4416 ;
  assign n4672 = n4670 | n4671 ;
  assign n4673 = x402 & ~n4416 ;
  assign n4674 = x1078 & n4416 ;
  assign n4675 = n4673 | n4674 ;
  assign n4676 = x403 & ~n4416 ;
  assign n4677 = x1045 & n4416 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = x404 & ~n4416 ;
  assign n4680 = x1084 & n4416 ;
  assign n4681 = n4679 | n4680 ;
  assign n4682 = x405 & ~n4416 ;
  assign n4683 = x1081 & n4416 ;
  assign n4684 = n4682 | n4683 ;
  assign n4685 = x406 & ~n4416 ;
  assign n4686 = x1076 & n4416 ;
  assign n4687 = n4685 | n4686 ;
  assign n4688 = x407 & ~n4416 ;
  assign n4689 = x1071 & n4416 ;
  assign n4690 = n4688 | n4689 ;
  assign n4691 = x408 & ~n4416 ;
  assign n4692 = x1068 & n4416 ;
  assign n4693 = n4691 | n4692 ;
  assign n4694 = x409 & ~n4416 ;
  assign n4695 = x1042 & n4416 ;
  assign n4696 = n4694 | n4695 ;
  assign n4697 = x410 & ~n4416 ;
  assign n4698 = x1059 & n4416 ;
  assign n4699 = n4697 | n4698 ;
  assign n4700 = x411 & ~n4416 ;
  assign n4701 = x1053 & n4416 ;
  assign n4702 = n4700 | n4701 ;
  assign n4703 = x412 & ~n4416 ;
  assign n4704 = x1037 & n4416 ;
  assign n4705 = n4703 | n4704 ;
  assign n4706 = x413 & ~n4416 ;
  assign n4707 = x1036 & n4416 ;
  assign n4708 = n4706 | n4707 ;
  assign n4709 = ~x331 & n4287 ;
  assign n4710 = ~x1049 & n4709 ;
  assign n4711 = x414 | n4709 ;
  assign n4712 = ~n4710 & n4711 ;
  assign n4713 = x415 & ~n4709 ;
  assign n4714 = x1062 & n4709 ;
  assign n4715 = n4713 | n4714 ;
  assign n4716 = x416 & ~n4709 ;
  assign n4717 = x1069 & n4709 ;
  assign n4718 = n4716 | n4717 ;
  assign n4719 = x417 & ~n4709 ;
  assign n4720 = x1039 & n4709 ;
  assign n4721 = n4719 | n4720 ;
  assign n4722 = x418 & ~n4709 ;
  assign n4723 = x1067 & n4709 ;
  assign n4724 = n4722 | n4723 ;
  assign n4725 = x419 & ~n4709 ;
  assign n4726 = x1080 & n4709 ;
  assign n4727 = n4725 | n4726 ;
  assign n4728 = x420 & ~n4709 ;
  assign n4729 = x1055 & n4709 ;
  assign n4730 = n4728 | n4729 ;
  assign n4731 = x421 & ~n4709 ;
  assign n4732 = x1051 & n4709 ;
  assign n4733 = n4731 | n4732 ;
  assign n4734 = x422 & ~n4709 ;
  assign n4735 = x1048 & n4709 ;
  assign n4736 = n4734 | n4735 ;
  assign n4737 = x423 & ~n4709 ;
  assign n4738 = x1087 & n4709 ;
  assign n4739 = n4737 | n4738 ;
  assign n4740 = x424 & ~n4709 ;
  assign n4741 = x1047 & n4709 ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = x425 & ~n4709 ;
  assign n4744 = x1035 & n4709 ;
  assign n4745 = n4743 | n4744 ;
  assign n4746 = x426 & ~n4709 ;
  assign n4747 = x1079 & n4709 ;
  assign n4748 = n4746 | n4747 ;
  assign n4749 = x427 & ~n4709 ;
  assign n4750 = x1078 & n4709 ;
  assign n4751 = n4749 | n4750 ;
  assign n4752 = x428 & ~n4709 ;
  assign n4753 = x1045 & n4709 ;
  assign n4754 = n4752 | n4753 ;
  assign n4755 = x429 & ~n4709 ;
  assign n4756 = x1084 & n4709 ;
  assign n4757 = n4755 | n4756 ;
  assign n4758 = x430 & ~n4709 ;
  assign n4759 = x1076 & n4709 ;
  assign n4760 = n4758 | n4759 ;
  assign n4761 = x431 & ~n4709 ;
  assign n4762 = x1071 & n4709 ;
  assign n4763 = n4761 | n4762 ;
  assign n4764 = x432 & ~n4709 ;
  assign n4765 = x1068 & n4709 ;
  assign n4766 = n4764 | n4765 ;
  assign n4767 = x433 & ~n4709 ;
  assign n4768 = x1042 & n4709 ;
  assign n4769 = n4767 | n4768 ;
  assign n4770 = x434 & ~n4709 ;
  assign n4771 = x1059 & n4709 ;
  assign n4772 = n4770 | n4771 ;
  assign n4773 = x435 & ~n4709 ;
  assign n4774 = x1053 & n4709 ;
  assign n4775 = n4773 | n4774 ;
  assign n4776 = x436 & ~n4709 ;
  assign n4777 = x1037 & n4709 ;
  assign n4778 = n4776 | n4777 ;
  assign n4779 = x437 & ~n4709 ;
  assign n4780 = x1070 & n4709 ;
  assign n4781 = n4779 | n4780 ;
  assign n4782 = x438 & ~n4709 ;
  assign n4783 = x1036 & n4709 ;
  assign n4784 = n4782 | n4783 ;
  assign n4785 = x439 & ~n4412 ;
  assign n4786 = x1057 & n4412 ;
  assign n4787 = n4785 | n4786 ;
  assign n4788 = x440 & ~n4412 ;
  assign n4789 = x1043 & n4412 ;
  assign n4790 = n4788 | n4789 ;
  assign n4791 = x441 & ~n4405 ;
  assign n4792 = x1044 & n4405 ;
  assign n4793 = n4791 | n4792 ;
  assign n4794 = x442 & ~n4412 ;
  assign n4795 = x1058 & n4412 ;
  assign n4796 = n4794 | n4795 ;
  assign n4797 = x443 & ~n4709 ;
  assign n4798 = x1044 & n4709 ;
  assign n4799 = n4797 | n4798 ;
  assign n4800 = x444 & ~n4709 ;
  assign n4801 = x1072 & n4709 ;
  assign n4802 = n4800 | n4801 ;
  assign n4803 = x445 & ~n4709 ;
  assign n4804 = x1081 & n4709 ;
  assign n4805 = n4803 | n4804 ;
  assign n4806 = x446 & ~n4709 ;
  assign n4807 = x1086 & n4709 ;
  assign n4808 = n4806 | n4807 ;
  assign n4809 = x447 & ~n4412 ;
  assign n4810 = x1040 & n4412 ;
  assign n4811 = n4809 | n4810 ;
  assign n4812 = x448 & ~n4709 ;
  assign n4813 = x1074 & n4709 ;
  assign n4814 = n4812 | n4813 ;
  assign n4815 = x449 & ~n4709 ;
  assign n4816 = x1057 & n4709 ;
  assign n4817 = n4815 | n4816 ;
  assign n4818 = x450 & ~n4405 ;
  assign n4819 = x1036 & n4405 ;
  assign n4820 = n4818 | n4819 ;
  assign n4821 = x451 & ~n4709 ;
  assign n4822 = x1063 & n4709 ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = x452 & ~n4405 ;
  assign n4825 = x1053 & n4405 ;
  assign n4826 = n4824 | n4825 ;
  assign n4827 = x453 & ~n4709 ;
  assign n4828 = x1040 & n4709 ;
  assign n4829 = n4827 | n4828 ;
  assign n4830 = x454 & ~n4709 ;
  assign n4831 = x1043 & n4709 ;
  assign n4832 = n4830 | n4831 ;
  assign n4833 = x455 & ~n4405 ;
  assign n4834 = x1037 & n4405 ;
  assign n4835 = n4833 | n4834 ;
  assign n4836 = x456 & ~n4416 ;
  assign n4837 = x1044 & n4416 ;
  assign n4838 = n4836 | n4837 ;
  assign n4839 = x594 & x597 ;
  assign n4840 = x601 & x605 ;
  assign n4841 = ( x600 & ~n4839 ) | ( x600 & n4840 ) | ( ~n4839 & n4840 ) ;
  assign n4842 = n4839 & n4841 ;
  assign n4843 = x804 & x810 ;
  assign n4844 = ~x599 & n4843 ;
  assign n4845 = ( ~x596 & x804 ) | ( ~x596 & n4844 ) | ( x804 & n4844 ) ;
  assign n4846 = x804 | x810 ;
  assign n4847 = x595 & x815 ;
  assign n4848 = n4846 & ~n4847 ;
  assign n4849 = n4845 | n4848 ;
  assign n4850 = n4842 & ~n4849 ;
  assign n4851 = n4840 | n4843 ;
  assign n4852 = x594 & x990 ;
  assign n4853 = x600 & ~x810 ;
  assign n4854 = ( x600 & n4852 ) | ( x600 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4855 = n4851 & n4854 ;
  assign n4856 = x605 & ~n4846 ;
  assign n4857 = ( ~x804 & n4840 ) | ( ~x804 & n4856 ) | ( n4840 & n4856 ) ;
  assign n4858 = n4855 | n4857 ;
  assign n4859 = ~x815 & x821 ;
  assign n4860 = n4858 & n4859 ;
  assign n4861 = ( x821 & n4850 ) | ( x821 & n4860 ) | ( n4850 & n4860 ) ;
  assign n4862 = x458 & ~n4405 ;
  assign n4863 = x1072 & n4405 ;
  assign n4864 = n4862 | n4863 ;
  assign n4865 = x459 & ~n4709 ;
  assign n4866 = x1058 & n4709 ;
  assign n4867 = n4865 | n4866 ;
  assign n4868 = x460 & ~n4405 ;
  assign n4869 = x1086 & n4405 ;
  assign n4870 = n4868 | n4869 ;
  assign n4871 = x461 & ~n4405 ;
  assign n4872 = x1057 & n4405 ;
  assign n4873 = n4871 | n4872 ;
  assign n4874 = x462 & ~n4405 ;
  assign n4875 = x1074 & n4405 ;
  assign n4876 = n4874 | n4875 ;
  assign n4877 = x463 & ~n4416 ;
  assign n4878 = x1070 & n4416 ;
  assign n4879 = n4877 | n4878 ;
  assign n4880 = x464 & ~n4709 ;
  assign n4881 = x1065 & n4709 ;
  assign n4882 = n4880 | n4881 ;
  assign n4883 = x1157 & n1523 ;
  assign n4884 = ~x243 & n1520 ;
  assign n4885 = x926 & n1518 ;
  assign n4886 = ( ~n4883 & n4884 ) | ( ~n4883 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4887 = n4883 | n4886 ;
  assign n4888 = x1151 & n1523 ;
  assign n4889 = x275 & n1520 ;
  assign n4890 = x943 & n1518 ;
  assign n4891 = ( ~n4888 & n4889 ) | ( ~n4888 & n4890 ) | ( n4889 & n4890 ) ;
  assign n4892 = n4888 | n4891 ;
  assign n4893 = x40 & ~x287 ;
  assign n4894 = ( ~x1001 & n1683 ) | ( ~x1001 & n4893 ) | ( n1683 & n4893 ) ;
  assign n4895 = n4893 & ~n4894 ;
  assign n4896 = ~n1691 & n4895 ;
  assign n4897 = n1254 | n4896 ;
  assign n4898 = ( n2804 & n4896 ) | ( n2804 & n4897 ) | ( n4896 & n4897 ) ;
  assign n4899 = x468 & ~n2149 ;
  assign n4900 = ( x468 & n1416 ) | ( x468 & n4899 ) | ( n1416 & n4899 ) ;
  assign n4901 = n2569 | n4900 ;
  assign n4902 = x1156 & n1523 ;
  assign n4903 = ~x263 & n1520 ;
  assign n4904 = x942 & n1518 ;
  assign n4905 = ( ~n4902 & n4903 ) | ( ~n4902 & n4904 ) | ( n4903 & n4904 ) ;
  assign n4906 = n4902 | n4905 ;
  assign n4907 = x1155 & n1523 ;
  assign n4908 = x267 & n1520 ;
  assign n4909 = x925 & n1518 ;
  assign n4910 = ( ~n4907 & n4908 ) | ( ~n4907 & n4909 ) | ( n4908 & n4909 ) ;
  assign n4911 = n4907 | n4910 ;
  assign n4912 = x1153 & n1523 ;
  assign n4913 = x253 & n1520 ;
  assign n4914 = x941 & n1518 ;
  assign n4915 = ( ~n4912 & n4913 ) | ( ~n4912 & n4914 ) | ( n4913 & n4914 ) ;
  assign n4916 = n4912 | n4915 ;
  assign n4917 = x1154 & n1523 ;
  assign n4918 = x254 & n1520 ;
  assign n4919 = x923 & n1518 ;
  assign n4920 = ( ~n4917 & n4918 ) | ( ~n4917 & n4919 ) | ( n4918 & n4919 ) ;
  assign n4921 = n4917 | n4920 ;
  assign n4922 = x1152 & n1523 ;
  assign n4923 = x268 & n1520 ;
  assign n4924 = x922 & n1518 ;
  assign n4925 = ( ~n4922 & n4923 ) | ( ~n4922 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4926 = n4922 | n4925 ;
  assign n4927 = x1150 & n1523 ;
  assign n4928 = x272 & n1520 ;
  assign n4929 = x931 & n1518 ;
  assign n4930 = ( ~n4927 & n4928 ) | ( ~n4927 & n4929 ) | ( n4928 & n4929 ) ;
  assign n4931 = n4927 | n4930 ;
  assign n4932 = x1149 & n1523 ;
  assign n4933 = x283 & n1520 ;
  assign n4934 = x936 & n1518 ;
  assign n4935 = ( ~n4932 & n4933 ) | ( ~n4932 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4936 = n4932 | n4935 ;
  assign n4937 = x71 & n2623 ;
  assign n4938 = x84 | n4937 ;
  assign n4939 = ( n2351 & n4937 ) | ( n2351 & n4938 ) | ( n4937 & n4938 ) ;
  assign n4940 = ( x71 & n2520 ) | ( x71 & ~n2521 ) | ( n2520 & ~n2521 ) ;
  assign n4941 = x248 & n3536 ;
  assign n4942 = x481 & ~n3536 ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = x249 & n3558 ;
  assign n4945 = x482 & ~n3558 ;
  assign n4946 = n4944 | n4945 ;
  assign n4947 = x242 & n3581 ;
  assign n4948 = x483 & ~n3581 ;
  assign n4949 = n4947 | n4948 ;
  assign n4950 = x249 & n3581 ;
  assign n4951 = x484 & ~n3581 ;
  assign n4952 = n4950 | n4951 ;
  assign n4953 = x234 & n3643 ;
  assign n4954 = x485 & ~n3643 ;
  assign n4955 = n4953 | n4954 ;
  assign n4956 = x244 & n3643 ;
  assign n4957 = x486 & ~n3643 ;
  assign n4958 = n4956 | n4957 ;
  assign n4959 = x246 & n3536 ;
  assign n4960 = x487 & ~n3536 ;
  assign n4961 = n4959 | n4960 ;
  assign n4962 = ~x239 & n3536 ;
  assign n4963 = x488 & ~n3536 ;
  assign n4964 = n4962 | n4963 ;
  assign n4965 = x242 & n3643 ;
  assign n4966 = x489 & ~n3643 ;
  assign n4967 = n4965 | n4966 ;
  assign n4968 = x241 & n3581 ;
  assign n4969 = x490 & ~n3581 ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = x238 & n3581 ;
  assign n4972 = x491 & ~n3581 ;
  assign n4973 = n4971 | n4972 ;
  assign n4974 = x240 & n3581 ;
  assign n4975 = x492 & ~n3581 ;
  assign n4976 = n4974 | n4975 ;
  assign n4977 = x244 & n3581 ;
  assign n4978 = x493 & ~n3581 ;
  assign n4979 = n4977 | n4978 ;
  assign n4980 = ~x239 & n3581 ;
  assign n4981 = x494 & ~n3581 ;
  assign n4982 = n4980 | n4981 ;
  assign n4983 = x235 & n3581 ;
  assign n4984 = x495 & ~n3581 ;
  assign n4985 = n4983 | n4984 ;
  assign n4986 = x249 & n3575 ;
  assign n4987 = x496 & ~n3575 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = ~x239 & n3575 ;
  assign n4990 = x497 & ~n3575 ;
  assign n4991 = n4989 | n4990 ;
  assign n4992 = x238 & n3558 ;
  assign n4993 = x498 & ~n3558 ;
  assign n4994 = n4992 | n4993 ;
  assign n4995 = x246 & n3575 ;
  assign n4996 = x499 & ~n3575 ;
  assign n4997 = n4995 | n4996 ;
  assign n4998 = x241 & n3575 ;
  assign n4999 = x500 & ~n3575 ;
  assign n5000 = n4998 | n4999 ;
  assign n5001 = x248 & n3575 ;
  assign n5002 = x501 & ~n3575 ;
  assign n5003 = n5001 | n5002 ;
  assign n5004 = x247 & n3575 ;
  assign n5005 = x502 & ~n3575 ;
  assign n5006 = n5004 | n5005 ;
  assign n5007 = x245 & n3575 ;
  assign n5008 = x503 & ~n3575 ;
  assign n5009 = n5007 | n5008 ;
  assign n5010 = x242 & n3564 ;
  assign n5011 = x504 & ~n3564 ;
  assign n5012 = n5010 | n5011 ;
  assign n5013 = x234 & n3575 ;
  assign n5014 = x505 & ~n3575 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = x241 & n3564 ;
  assign n5017 = x506 & ~n3564 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = x238 & n3564 ;
  assign n5020 = x507 & ~n3564 ;
  assign n5021 = n5019 | n5020 ;
  assign n5022 = x247 & n3564 ;
  assign n5023 = x508 & ~n3564 ;
  assign n5024 = n5022 | n5023 ;
  assign n5025 = x245 & n3564 ;
  assign n5026 = x509 & ~n3564 ;
  assign n5027 = n5025 | n5026 ;
  assign n5028 = x242 & n3536 ;
  assign n5029 = x510 & ~n3536 ;
  assign n5030 = n5028 | n5029 ;
  assign n5031 = x234 & n3536 ;
  assign n5032 = x511 & ~n3536 ;
  assign n5033 = n5031 | n5032 ;
  assign n5034 = x235 & n3536 ;
  assign n5035 = x512 & ~n3536 ;
  assign n5036 = n5034 | n5035 ;
  assign n5037 = x244 & n3536 ;
  assign n5038 = x513 & ~n3536 ;
  assign n5039 = n5037 | n5038 ;
  assign n5040 = x245 & n3536 ;
  assign n5041 = x514 & ~n3536 ;
  assign n5042 = n5040 | n5041 ;
  assign n5043 = x240 & n3536 ;
  assign n5044 = x515 & ~n3536 ;
  assign n5045 = n5043 | n5044 ;
  assign n5046 = x247 & n3536 ;
  assign n5047 = x516 & ~n3536 ;
  assign n5048 = n5046 | n5047 ;
  assign n5049 = x238 & n3536 ;
  assign n5050 = x517 & ~n3536 ;
  assign n5051 = n5049 | n5050 ;
  assign n5052 = x234 & n3552 ;
  assign n5053 = x518 & ~n3552 ;
  assign n5054 = n5052 | n5053 ;
  assign n5055 = ~x239 & n3552 ;
  assign n5056 = x519 & ~n3552 ;
  assign n5057 = n5055 | n5056 ;
  assign n5058 = x246 & n3552 ;
  assign n5059 = x520 & ~n3552 ;
  assign n5060 = n5058 | n5059 ;
  assign n5061 = x248 & n3552 ;
  assign n5062 = x521 & ~n3552 ;
  assign n5063 = n5061 | n5062 ;
  assign n5064 = x238 & n3552 ;
  assign n5065 = x522 & ~n3552 ;
  assign n5066 = n5064 | n5065 ;
  assign n5067 = x234 & n3653 ;
  assign n5068 = x523 & ~n3653 ;
  assign n5069 = n5067 | n5068 ;
  assign n5070 = ~x239 & n3653 ;
  assign n5071 = x524 & ~n3653 ;
  assign n5072 = n5070 | n5071 ;
  assign n5073 = x245 & n3653 ;
  assign n5074 = x525 & ~n3653 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = x246 & n3653 ;
  assign n5077 = x526 & ~n3653 ;
  assign n5078 = n5076 | n5077 ;
  assign n5079 = x247 & n3653 ;
  assign n5080 = x527 & ~n3653 ;
  assign n5081 = n5079 | n5080 ;
  assign n5082 = x249 & n3653 ;
  assign n5083 = x528 & ~n3653 ;
  assign n5084 = n5082 | n5083 ;
  assign n5085 = x238 & n3653 ;
  assign n5086 = x529 & ~n3653 ;
  assign n5087 = n5085 | n5086 ;
  assign n5088 = x240 & n3653 ;
  assign n5089 = x530 & ~n3653 ;
  assign n5090 = n5088 | n5089 ;
  assign n5091 = x235 & n3558 ;
  assign n5092 = x531 & ~n3558 ;
  assign n5093 = n5091 | n5092 ;
  assign n5094 = x247 & n3558 ;
  assign n5095 = x532 & ~n3558 ;
  assign n5096 = n5094 | n5095 ;
  assign n5097 = x235 & n3564 ;
  assign n5098 = x533 & ~n3564 ;
  assign n5099 = n5097 | n5098 ;
  assign n5100 = ~x239 & n3564 ;
  assign n5101 = x534 & ~n3564 ;
  assign n5102 = n5100 | n5101 ;
  assign n5103 = x240 & n3564 ;
  assign n5104 = x535 & ~n3564 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = x246 & n3564 ;
  assign n5107 = x536 & ~n3564 ;
  assign n5108 = n5106 | n5107 ;
  assign n5109 = x248 & n3564 ;
  assign n5110 = x537 & ~n3564 ;
  assign n5111 = n5109 | n5110 ;
  assign n5112 = x249 & n3564 ;
  assign n5113 = x538 & ~n3564 ;
  assign n5114 = n5112 | n5113 ;
  assign n5115 = x242 & n3575 ;
  assign n5116 = x539 & ~n3575 ;
  assign n5117 = n5115 | n5116 ;
  assign n5118 = x235 & n3575 ;
  assign n5119 = x540 & ~n3575 ;
  assign n5120 = n5118 | n5119 ;
  assign n5121 = x244 & n3575 ;
  assign n5122 = x541 & ~n3575 ;
  assign n5123 = n5121 | n5122 ;
  assign n5124 = x240 & n3575 ;
  assign n5125 = x542 & ~n3575 ;
  assign n5126 = n5124 | n5125 ;
  assign n5127 = x238 & n3575 ;
  assign n5128 = x543 & ~n3575 ;
  assign n5129 = n5127 | n5128 ;
  assign n5130 = x234 & n3581 ;
  assign n5131 = x544 & ~n3581 ;
  assign n5132 = n5130 | n5131 ;
  assign n5133 = x245 & n3581 ;
  assign n5134 = x545 & ~n3581 ;
  assign n5135 = n5133 | n5134 ;
  assign n5136 = x246 & n3581 ;
  assign n5137 = x546 & ~n3581 ;
  assign n5138 = n5136 | n5137 ;
  assign n5139 = x247 & n3581 ;
  assign n5140 = x547 & ~n3581 ;
  assign n5141 = n5139 | n5140 ;
  assign n5142 = x248 & n3581 ;
  assign n5143 = x548 & ~n3581 ;
  assign n5144 = n5142 | n5143 ;
  assign n5145 = x235 & n3643 ;
  assign n5146 = x549 & ~n3643 ;
  assign n5147 = n5145 | n5146 ;
  assign n5148 = ~x239 & n3643 ;
  assign n5149 = x550 & ~n3643 ;
  assign n5150 = n5148 | n5149 ;
  assign n5151 = x240 & n3643 ;
  assign n5152 = x551 & ~n3643 ;
  assign n5153 = n5151 | n5152 ;
  assign n5154 = x247 & n3643 ;
  assign n5155 = x552 & ~n3643 ;
  assign n5156 = n5154 | n5155 ;
  assign n5157 = x241 & n3643 ;
  assign n5158 = x553 & ~n3643 ;
  assign n5159 = n5157 | n5158 ;
  assign n5160 = x248 & n3643 ;
  assign n5161 = x554 & ~n3643 ;
  assign n5162 = n5160 | n5161 ;
  assign n5163 = x249 & n3643 ;
  assign n5164 = x555 & ~n3643 ;
  assign n5165 = n5163 | n5164 ;
  assign n5166 = x242 & n3558 ;
  assign n5167 = x556 & ~n3558 ;
  assign n5168 = n5166 | n5167 ;
  assign n5169 = x234 & n3564 ;
  assign n5170 = x557 & ~n3564 ;
  assign n5171 = n5169 | n5170 ;
  assign n5172 = x244 & n3564 ;
  assign n5173 = x558 & ~n3564 ;
  assign n5174 = n5172 | n5173 ;
  assign n5175 = x241 & n3536 ;
  assign n5176 = x559 & ~n3536 ;
  assign n5177 = n5175 | n5176 ;
  assign n5178 = x240 & n3558 ;
  assign n5179 = x560 & ~n3558 ;
  assign n5180 = n5178 | n5179 ;
  assign n5181 = x247 & n3552 ;
  assign n5182 = x561 & ~n3552 ;
  assign n5183 = n5181 | n5182 ;
  assign n5184 = x241 & n3558 ;
  assign n5185 = x562 & ~n3558 ;
  assign n5186 = n5184 | n5185 ;
  assign n5187 = x246 & n3643 ;
  assign n5188 = x563 & ~n3643 ;
  assign n5189 = n5187 | n5188 ;
  assign n5190 = x246 & n3558 ;
  assign n5191 = x564 & ~n3558 ;
  assign n5192 = n5190 | n5191 ;
  assign n5193 = x248 & n3558 ;
  assign n5194 = x565 & ~n3558 ;
  assign n5195 = n5193 | n5194 ;
  assign n5196 = x244 & n3558 ;
  assign n5197 = x566 & ~n3558 ;
  assign n5198 = n5196 | n5197 ;
  assign n5199 = x230 & n1841 ;
  assign n5200 = ( ~x567 & x1092 ) | ( ~x567 & n5199 ) | ( x1092 & n5199 ) ;
  assign n5201 = n3217 & n3218 ;
  assign n5202 = n5199 & ~n5201 ;
  assign n5203 = n3185 & n3186 ;
  assign n5204 = n5200 & n5203 ;
  assign n5205 = ( n5200 & ~n5202 ) | ( n5200 & n5204 ) | ( ~n5202 & n5204 ) ;
  assign n5206 = x245 & n3558 ;
  assign n5207 = x568 & ~n3558 ;
  assign n5208 = n5206 | n5207 ;
  assign n5209 = ~x239 & n3558 ;
  assign n5210 = x569 & ~n3558 ;
  assign n5211 = n5209 | n5210 ;
  assign n5212 = x234 & n3558 ;
  assign n5213 = x570 & ~n3558 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = x241 & n3653 ;
  assign n5216 = x571 & ~n3653 ;
  assign n5217 = n5215 | n5216 ;
  assign n5218 = x244 & n3653 ;
  assign n5219 = x572 & ~n3653 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = x242 & n3653 ;
  assign n5222 = x573 & ~n3653 ;
  assign n5223 = n5221 | n5222 ;
  assign n5224 = x241 & n3552 ;
  assign n5225 = x574 & ~n3552 ;
  assign n5226 = n5224 | n5225 ;
  assign n5227 = x235 & n3653 ;
  assign n5228 = x575 & ~n3653 ;
  assign n5229 = n5227 | n5228 ;
  assign n5230 = x248 & n3653 ;
  assign n5231 = x576 & ~n3653 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = x238 & n3643 ;
  assign n5234 = x577 & ~n3643 ;
  assign n5235 = n5233 | n5234 ;
  assign n5236 = x249 & n3552 ;
  assign n5237 = x578 & ~n3552 ;
  assign n5238 = n5236 | n5237 ;
  assign n5239 = x249 & n3536 ;
  assign n5240 = x579 & ~n3536 ;
  assign n5241 = n5239 | n5240 ;
  assign n5242 = x245 & n3643 ;
  assign n5243 = x580 & ~n3643 ;
  assign n5244 = n5242 | n5243 ;
  assign n5245 = x235 & n3552 ;
  assign n5246 = x581 & ~n3552 ;
  assign n5247 = n5245 | n5246 ;
  assign n5248 = x240 & n3552 ;
  assign n5249 = x582 & ~n3552 ;
  assign n5250 = n5248 | n5249 ;
  assign n5251 = x245 & n3552 ;
  assign n5252 = x584 & ~n3552 ;
  assign n5253 = n5251 | n5252 ;
  assign n5254 = x244 & n3552 ;
  assign n5255 = x585 & ~n3552 ;
  assign n5256 = n5254 | n5255 ;
  assign n5257 = x242 & n3552 ;
  assign n5258 = x586 & ~n3552 ;
  assign n5259 = n5257 | n5258 ;
  assign n5260 = ~x230 & x587 ;
  assign n5261 = x230 | x587 ;
  assign n5262 = ( n3187 & n5260 ) | ( n3187 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = ~x123 & n1870 ;
  assign n5264 = x588 & ~n5263 ;
  assign n5265 = x591 & n5263 ;
  assign n5266 = ( n4453 & n5264 ) | ( n4453 & n5265 ) | ( n5264 & n5265 ) ;
  assign n5267 = x220 & n3580 ;
  assign n5268 = x203 & ~n3557 ;
  assign n5269 = x201 & n3535 ;
  assign n5270 = ( ~n5267 & n5268 ) | ( ~n5267 & n5269 ) | ( n5268 & n5269 ) ;
  assign n5271 = x202 & n3551 ;
  assign n5272 = n5267 | n5271 ;
  assign n5273 = n5270 | n5272 ;
  assign n5274 = n1797 & ~n5273 ;
  assign n5275 = x204 & x233 ;
  assign n5276 = x205 & ~x233 ;
  assign n5277 = ( x237 & n5275 ) | ( x237 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5278 = x218 & ~x233 ;
  assign n5279 = x206 & x233 ;
  assign n5280 = ( ~x237 & n5278 ) | ( ~x237 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = n5277 | n5280 ;
  assign n5282 = n1791 & ~n5281 ;
  assign n5283 = n5274 | n5282 ;
  assign n5284 = x590 | n5263 ;
  assign n5285 = ~x588 & n5263 ;
  assign n5286 = ( n4453 & ~n5284 ) | ( n4453 & n5285 ) | ( ~n5284 & n5285 ) ;
  assign n5287 = x591 & ~n5263 ;
  assign n5288 = x592 & n5263 ;
  assign n5289 = ( n4453 & n5287 ) | ( n4453 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5290 = x592 & ~n5263 ;
  assign n5291 = x590 & n5263 ;
  assign n5292 = ( n4453 & n5290 ) | ( n4453 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5293 = ~x247 & x532 ;
  assign n5294 = ( ~x245 & x568 ) | ( ~x245 & n5293 ) | ( x568 & n5293 ) ;
  assign n5295 = x247 & ~x532 ;
  assign n5296 = ( x245 & ~x568 ) | ( x245 & n5295 ) | ( ~x568 & n5295 ) ;
  assign n5297 = n5294 | n5296 ;
  assign n5298 = ~x240 & x560 ;
  assign n5299 = ( ~x238 & x498 ) | ( ~x238 & n5298 ) | ( x498 & n5298 ) ;
  assign n5300 = x240 & ~x560 ;
  assign n5301 = ( x238 & ~x498 ) | ( x238 & n5300 ) | ( ~x498 & n5300 ) ;
  assign n5302 = n5299 | n5301 ;
  assign n5303 = ~x242 & x556 ;
  assign n5304 = ( ~x235 & x531 ) | ( ~x235 & n5303 ) | ( x531 & n5303 ) ;
  assign n5305 = x242 & ~x556 ;
  assign n5306 = ( x235 & ~x531 ) | ( x235 & n5305 ) | ( ~x531 & n5305 ) ;
  assign n5307 = n5304 | n5306 ;
  assign n5308 = ( ~n5297 & n5302 ) | ( ~n5297 & n5307 ) | ( n5302 & n5307 ) ;
  assign n5309 = n5297 | n5308 ;
  assign n5310 = ~x249 & x482 ;
  assign n5311 = ( ~x248 & x565 ) | ( ~x248 & n5310 ) | ( x565 & n5310 ) ;
  assign n5312 = x249 & ~x482 ;
  assign n5313 = ( x248 & ~x565 ) | ( x248 & n5312 ) | ( ~x565 & n5312 ) ;
  assign n5314 = n5311 | n5313 ;
  assign n5315 = ~x244 & x566 ;
  assign n5316 = ( ~x241 & x562 ) | ( ~x241 & n5315 ) | ( x562 & n5315 ) ;
  assign n5317 = x244 & ~x566 ;
  assign n5318 = ( x241 & ~x562 ) | ( x241 & n5317 ) | ( ~x562 & n5317 ) ;
  assign n5319 = n5316 | n5318 ;
  assign n5320 = n5314 | n5319 ;
  assign n5321 = ( ~x234 & x570 ) | ( ~x234 & n5320 ) | ( x570 & n5320 ) ;
  assign n5322 = ~x246 & x564 ;
  assign n5323 = ( x239 & x569 ) | ( x239 & n5322 ) | ( x569 & n5322 ) ;
  assign n5324 = x246 & ~x564 ;
  assign n5325 = ( x239 & x569 ) | ( x239 & ~n5324 ) | ( x569 & ~n5324 ) ;
  assign n5326 = ~n5323 & n5325 ;
  assign n5327 = ( ~x234 & x570 ) | ( ~x234 & n5326 ) | ( x570 & n5326 ) ;
  assign n5328 = ( n5309 & ~n5321 ) | ( n5309 & n5327 ) | ( ~n5321 & n5327 ) ;
  assign n5329 = ( n1797 & n5309 ) | ( n1797 & ~n5328 ) | ( n5309 & ~n5328 ) ;
  assign n5330 = n1797 | n3557 ;
  assign n5331 = ( n3557 & ~n5329 ) | ( n3557 & n5330 ) | ( ~n5329 & n5330 ) ;
  assign n5332 = ~x248 & x554 ;
  assign n5333 = ( ~x234 & x485 ) | ( ~x234 & n5332 ) | ( x485 & n5332 ) ;
  assign n5334 = x248 & ~x554 ;
  assign n5335 = ( x234 & ~x485 ) | ( x234 & n5334 ) | ( ~x485 & n5334 ) ;
  assign n5336 = n5333 | n5335 ;
  assign n5337 = ~x242 & x489 ;
  assign n5338 = ( ~x235 & x549 ) | ( ~x235 & n5337 ) | ( x549 & n5337 ) ;
  assign n5339 = x242 & ~x489 ;
  assign n5340 = ( x235 & ~x549 ) | ( x235 & n5339 ) | ( ~x549 & n5339 ) ;
  assign n5341 = n5338 | n5340 ;
  assign n5342 = x239 & x550 ;
  assign n5343 = ( ~x238 & x577 ) | ( ~x238 & n5342 ) | ( x577 & n5342 ) ;
  assign n5344 = x239 | x550 ;
  assign n5345 = ( ~x238 & x577 ) | ( ~x238 & n5344 ) | ( x577 & n5344 ) ;
  assign n5346 = ~n5343 & n5345 ;
  assign n5347 = ( n5336 & ~n5341 ) | ( n5336 & n5346 ) | ( ~n5341 & n5346 ) ;
  assign n5348 = ~x241 & x553 ;
  assign n5349 = ( ~x240 & x551 ) | ( ~x240 & n5348 ) | ( x551 & n5348 ) ;
  assign n5350 = x241 & ~x553 ;
  assign n5351 = ( x240 & ~x551 ) | ( x240 & n5350 ) | ( ~x551 & n5350 ) ;
  assign n5352 = n5349 | n5351 ;
  assign n5353 = n5336 | n5352 ;
  assign n5354 = n5347 & ~n5353 ;
  assign n5355 = ~x247 & x552 ;
  assign n5356 = ( ~x244 & x486 ) | ( ~x244 & n5355 ) | ( x486 & n5355 ) ;
  assign n5357 = x247 & ~x552 ;
  assign n5358 = ( x244 & ~x486 ) | ( x244 & n5357 ) | ( ~x486 & n5357 ) ;
  assign n5359 = n5356 | n5358 ;
  assign n5360 = ( x249 & ~x555 ) | ( x249 & n5359 ) | ( ~x555 & n5359 ) ;
  assign n5361 = ~x246 & x563 ;
  assign n5362 = ( ~x245 & x580 ) | ( ~x245 & n5361 ) | ( x580 & n5361 ) ;
  assign n5363 = x246 & ~x563 ;
  assign n5364 = ( x245 & ~x580 ) | ( x245 & n5363 ) | ( ~x580 & n5363 ) ;
  assign n5365 = n5362 | n5364 ;
  assign n5366 = ( ~x249 & x555 ) | ( ~x249 & n5365 ) | ( x555 & n5365 ) ;
  assign n5367 = n5360 | n5366 ;
  assign n5368 = ( ~n1791 & n5354 ) | ( ~n1791 & n5367 ) | ( n5354 & n5367 ) ;
  assign n5369 = n5354 & ~n5368 ;
  assign n5370 = n5331 | n5369 ;
  assign n5371 = ~x244 & x572 ;
  assign n5372 = ( ~x242 & x573 ) | ( ~x242 & n5371 ) | ( x573 & n5371 ) ;
  assign n5373 = x244 & ~x572 ;
  assign n5374 = ( x242 & ~x573 ) | ( x242 & n5373 ) | ( ~x573 & n5373 ) ;
  assign n5375 = n5372 | n5374 ;
  assign n5376 = n3580 & n5375 ;
  assign n5377 = ~x246 & x526 ;
  assign n5378 = ( ~x238 & x529 ) | ( ~x238 & n5377 ) | ( x529 & n5377 ) ;
  assign n5379 = x246 & ~x526 ;
  assign n5380 = ( x238 & ~x529 ) | ( x238 & n5379 ) | ( ~x529 & n5379 ) ;
  assign n5381 = n5378 | n5380 ;
  assign n5382 = ~x241 & x571 ;
  assign n5383 = ( x239 & x524 ) | ( x239 & n5382 ) | ( x524 & n5382 ) ;
  assign n5384 = x241 & ~x571 ;
  assign n5385 = ( x239 & x524 ) | ( x239 & ~n5384 ) | ( x524 & ~n5384 ) ;
  assign n5386 = ~n5383 & n5385 ;
  assign n5387 = ~x249 & x528 ;
  assign n5388 = ( ~x235 & x575 ) | ( ~x235 & n5387 ) | ( x575 & n5387 ) ;
  assign n5389 = x249 & ~x528 ;
  assign n5390 = ( x235 & ~x575 ) | ( x235 & n5389 ) | ( ~x575 & n5389 ) ;
  assign n5391 = n5388 | n5390 ;
  assign n5392 = ( n5381 & n5386 ) | ( n5381 & ~n5391 ) | ( n5386 & ~n5391 ) ;
  assign n5393 = ~x245 & x525 ;
  assign n5394 = ( ~x234 & x523 ) | ( ~x234 & n5393 ) | ( x523 & n5393 ) ;
  assign n5395 = x245 & ~x525 ;
  assign n5396 = ( x234 & ~x523 ) | ( x234 & n5395 ) | ( ~x523 & n5395 ) ;
  assign n5397 = n5394 | n5396 ;
  assign n5398 = n5381 | n5397 ;
  assign n5399 = n5392 & ~n5398 ;
  assign n5400 = ( x248 & ~x576 ) | ( x248 & n5399 ) | ( ~x576 & n5399 ) ;
  assign n5401 = ~x247 & x527 ;
  assign n5402 = ( ~x240 & x530 ) | ( ~x240 & n5401 ) | ( x530 & n5401 ) ;
  assign n5403 = x247 & ~x527 ;
  assign n5404 = ( x240 & ~x530 ) | ( x240 & n5403 ) | ( ~x530 & n5403 ) ;
  assign n5405 = n5402 | n5404 ;
  assign n5406 = ( x248 & ~x576 ) | ( x248 & n5405 ) | ( ~x576 & n5405 ) ;
  assign n5407 = n5400 & ~n5406 ;
  assign n5408 = n1797 & n5407 ;
  assign n5409 = ( n3580 & n5376 ) | ( n3580 & ~n5408 ) | ( n5376 & ~n5408 ) ;
  assign n5410 = ~x241 & x490 ;
  assign n5411 = ( ~x235 & x495 ) | ( ~x235 & n5410 ) | ( x495 & n5410 ) ;
  assign n5412 = x241 & ~x490 ;
  assign n5413 = ( x235 & ~x495 ) | ( x235 & n5412 ) | ( ~x495 & n5412 ) ;
  assign n5414 = n5411 | n5413 ;
  assign n5415 = ~x248 & x548 ;
  assign n5416 = ( ~x246 & x546 ) | ( ~x246 & n5415 ) | ( x546 & n5415 ) ;
  assign n5417 = x248 & ~x548 ;
  assign n5418 = ( x246 & ~x546 ) | ( x246 & n5417 ) | ( ~x546 & n5417 ) ;
  assign n5419 = n5416 | n5418 ;
  assign n5420 = ~x238 & x491 ;
  assign n5421 = ( ~x234 & x544 ) | ( ~x234 & n5420 ) | ( x544 & n5420 ) ;
  assign n5422 = x238 & ~x491 ;
  assign n5423 = ( x234 & ~x544 ) | ( x234 & n5422 ) | ( ~x544 & n5422 ) ;
  assign n5424 = n5421 | n5423 ;
  assign n5425 = ( ~n5414 & n5419 ) | ( ~n5414 & n5424 ) | ( n5419 & n5424 ) ;
  assign n5426 = ~x249 & x484 ;
  assign n5427 = ( ~x242 & x483 ) | ( ~x242 & n5426 ) | ( x483 & n5426 ) ;
  assign n5428 = x249 & ~x484 ;
  assign n5429 = ( x242 & ~x483 ) | ( x242 & n5428 ) | ( ~x483 & n5428 ) ;
  assign n5430 = n5427 | n5429 ;
  assign n5431 = n5414 | n5430 ;
  assign n5432 = n5425 | n5431 ;
  assign n5433 = ( ~x247 & x547 ) | ( ~x247 & n5432 ) | ( x547 & n5432 ) ;
  assign n5434 = ~x240 & x492 ;
  assign n5435 = ( x239 & x494 ) | ( x239 & n5434 ) | ( x494 & n5434 ) ;
  assign n5436 = x240 & ~x492 ;
  assign n5437 = ( x239 & x494 ) | ( x239 & ~n5436 ) | ( x494 & ~n5436 ) ;
  assign n5438 = ~n5435 & n5437 ;
  assign n5439 = ( ~x247 & x547 ) | ( ~x247 & n5438 ) | ( x547 & n5438 ) ;
  assign n5440 = ~n5433 & n5439 ;
  assign n5441 = ~x245 & x545 ;
  assign n5442 = ( ~x244 & x493 ) | ( ~x244 & n5441 ) | ( x493 & n5441 ) ;
  assign n5443 = x245 & ~x545 ;
  assign n5444 = ( x244 & ~x493 ) | ( x244 & n5443 ) | ( ~x493 & n5443 ) ;
  assign n5445 = n5442 | n5444 ;
  assign n5446 = ( n1791 & ~n5440 ) | ( n1791 & n5445 ) | ( ~n5440 & n5445 ) ;
  assign n5447 = ( n1791 & ~n5409 ) | ( n1791 & n5446 ) | ( ~n5409 & n5446 ) ;
  assign n5448 = n1791 & ~n5447 ;
  assign n5449 = ( n5370 & ~n5409 ) | ( n5370 & n5448 ) | ( ~n5409 & n5448 ) ;
  assign n5450 = ~x249 & x578 ;
  assign n5451 = ( ~x234 & x518 ) | ( ~x234 & n5450 ) | ( x518 & n5450 ) ;
  assign n5452 = x249 & ~x578 ;
  assign n5453 = ( x234 & ~x518 ) | ( x234 & n5452 ) | ( ~x518 & n5452 ) ;
  assign n5454 = n5451 | n5453 ;
  assign n5455 = n3551 & n5454 ;
  assign n5456 = ~x248 & x521 ;
  assign n5457 = ( ~x246 & x520 ) | ( ~x246 & n5456 ) | ( x520 & n5456 ) ;
  assign n5458 = x248 & ~x521 ;
  assign n5459 = ( x246 & ~x520 ) | ( x246 & n5458 ) | ( ~x520 & n5458 ) ;
  assign n5460 = n5457 | n5459 ;
  assign n5461 = ~x245 & x584 ;
  assign n5462 = ( ~x241 & x574 ) | ( ~x241 & n5461 ) | ( x574 & n5461 ) ;
  assign n5463 = x245 & ~x584 ;
  assign n5464 = ( x241 & ~x574 ) | ( x241 & n5463 ) | ( ~x574 & n5463 ) ;
  assign n5465 = n5462 | n5464 ;
  assign n5466 = ~x247 & x561 ;
  assign n5467 = ( ~x238 & x522 ) | ( ~x238 & n5466 ) | ( x522 & n5466 ) ;
  assign n5468 = x247 & ~x561 ;
  assign n5469 = ( x238 & ~x522 ) | ( x238 & n5468 ) | ( ~x522 & n5468 ) ;
  assign n5470 = n5467 | n5469 ;
  assign n5471 = ( ~n5460 & n5465 ) | ( ~n5460 & n5470 ) | ( n5465 & n5470 ) ;
  assign n5472 = ~x242 & x586 ;
  assign n5473 = ( ~x240 & x582 ) | ( ~x240 & n5472 ) | ( x582 & n5472 ) ;
  assign n5474 = x242 & ~x586 ;
  assign n5475 = ( x240 & ~x582 ) | ( x240 & n5474 ) | ( ~x582 & n5474 ) ;
  assign n5476 = n5473 | n5475 ;
  assign n5477 = n5460 | n5476 ;
  assign n5478 = n5471 | n5477 ;
  assign n5479 = ( ~x235 & x581 ) | ( ~x235 & n5478 ) | ( x581 & n5478 ) ;
  assign n5480 = ~x244 & x585 ;
  assign n5481 = ( x239 & x519 ) | ( x239 & n5480 ) | ( x519 & n5480 ) ;
  assign n5482 = x244 & ~x585 ;
  assign n5483 = ( x239 & x519 ) | ( x239 & ~n5482 ) | ( x519 & ~n5482 ) ;
  assign n5484 = ~n5481 & n5483 ;
  assign n5485 = ( ~x235 & x581 ) | ( ~x235 & n5484 ) | ( x581 & n5484 ) ;
  assign n5486 = ~n5479 & n5485 ;
  assign n5487 = n1797 & n5486 ;
  assign n5488 = ( n3551 & n5455 ) | ( n3551 & ~n5487 ) | ( n5455 & ~n5487 ) ;
  assign n5489 = ~x248 & x501 ;
  assign n5490 = ( ~x242 & x539 ) | ( ~x242 & n5489 ) | ( x539 & n5489 ) ;
  assign n5491 = x248 & ~x501 ;
  assign n5492 = ( x242 & ~x539 ) | ( x242 & n5491 ) | ( ~x539 & n5491 ) ;
  assign n5493 = n5490 | n5492 ;
  assign n5494 = n1791 & ~n5493 ;
  assign n5495 = ~x247 & x502 ;
  assign n5496 = ( ~x235 & x540 ) | ( ~x235 & n5495 ) | ( x540 & n5495 ) ;
  assign n5497 = x247 & ~x502 ;
  assign n5498 = ( x235 & ~x540 ) | ( x235 & n5497 ) | ( ~x540 & n5497 ) ;
  assign n5499 = n5496 | n5498 ;
  assign n5500 = ~x244 & x541 ;
  assign n5501 = ( x239 & x497 ) | ( x239 & n5500 ) | ( x497 & n5500 ) ;
  assign n5502 = x244 & ~x541 ;
  assign n5503 = ( x239 & x497 ) | ( x239 & ~n5502 ) | ( x497 & ~n5502 ) ;
  assign n5504 = ~n5501 & n5503 ;
  assign n5505 = ~x240 & x542 ;
  assign n5506 = ( ~x234 & x505 ) | ( ~x234 & n5505 ) | ( x505 & n5505 ) ;
  assign n5507 = x240 & ~x542 ;
  assign n5508 = ( x234 & ~x505 ) | ( x234 & n5507 ) | ( ~x505 & n5507 ) ;
  assign n5509 = n5506 | n5508 ;
  assign n5510 = ( n5499 & n5504 ) | ( n5499 & ~n5509 ) | ( n5504 & ~n5509 ) ;
  assign n5511 = ~x249 & x496 ;
  assign n5512 = ( ~x246 & x499 ) | ( ~x246 & n5511 ) | ( x499 & n5511 ) ;
  assign n5513 = x249 & ~x496 ;
  assign n5514 = ( x246 & ~x499 ) | ( x246 & n5513 ) | ( ~x499 & n5513 ) ;
  assign n5515 = n5512 | n5514 ;
  assign n5516 = n5499 | n5515 ;
  assign n5517 = n5510 & ~n5516 ;
  assign n5518 = ( x238 & ~x543 ) | ( x238 & n5517 ) | ( ~x543 & n5517 ) ;
  assign n5519 = ~x245 & x503 ;
  assign n5520 = ( ~x241 & x500 ) | ( ~x241 & n5519 ) | ( x500 & n5519 ) ;
  assign n5521 = x245 & ~x503 ;
  assign n5522 = ( x241 & ~x500 ) | ( x241 & n5521 ) | ( ~x500 & n5521 ) ;
  assign n5523 = n5520 | n5522 ;
  assign n5524 = ( x238 & ~x543 ) | ( x238 & n5523 ) | ( ~x543 & n5523 ) ;
  assign n5525 = n5518 & ~n5524 ;
  assign n5526 = n5494 & n5525 ;
  assign n5527 = n5488 & ~n5526 ;
  assign n5528 = ~x241 & x506 ;
  assign n5529 = ( ~x238 & x507 ) | ( ~x238 & n5528 ) | ( x507 & n5528 ) ;
  assign n5530 = x241 & ~x506 ;
  assign n5531 = ( x238 & ~x507 ) | ( x238 & n5530 ) | ( ~x507 & n5530 ) ;
  assign n5532 = n5529 | n5531 ;
  assign n5533 = n1791 & ~n5532 ;
  assign n5534 = ~x247 & x508 ;
  assign n5535 = ( ~x245 & x509 ) | ( ~x245 & n5534 ) | ( x509 & n5534 ) ;
  assign n5536 = x247 & ~x508 ;
  assign n5537 = ( x245 & ~x509 ) | ( x245 & n5536 ) | ( ~x509 & n5536 ) ;
  assign n5538 = n5535 | n5537 ;
  assign n5539 = x239 & x534 ;
  assign n5540 = ( ~x235 & x533 ) | ( ~x235 & n5539 ) | ( x533 & n5539 ) ;
  assign n5541 = x239 | x534 ;
  assign n5542 = ( ~x235 & x533 ) | ( ~x235 & n5541 ) | ( x533 & n5541 ) ;
  assign n5543 = ~n5540 & n5542 ;
  assign n5544 = ~x244 & x558 ;
  assign n5545 = ( ~x240 & x535 ) | ( ~x240 & n5544 ) | ( x535 & n5544 ) ;
  assign n5546 = x244 & ~x558 ;
  assign n5547 = ( x240 & ~x535 ) | ( x240 & n5546 ) | ( ~x535 & n5546 ) ;
  assign n5548 = n5545 | n5547 ;
  assign n5549 = ( n5538 & n5543 ) | ( n5538 & ~n5548 ) | ( n5543 & ~n5548 ) ;
  assign n5550 = ~x246 & x536 ;
  assign n5551 = ( ~x242 & x504 ) | ( ~x242 & n5550 ) | ( x504 & n5550 ) ;
  assign n5552 = x246 & ~x536 ;
  assign n5553 = ( x242 & ~x504 ) | ( x242 & n5552 ) | ( ~x504 & n5552 ) ;
  assign n5554 = n5551 | n5553 ;
  assign n5555 = n5538 | n5554 ;
  assign n5556 = n5549 & ~n5555 ;
  assign n5557 = ( x249 & ~x538 ) | ( x249 & n5556 ) | ( ~x538 & n5556 ) ;
  assign n5558 = ~x248 & x537 ;
  assign n5559 = ( ~x234 & x557 ) | ( ~x234 & n5558 ) | ( x557 & n5558 ) ;
  assign n5560 = x248 & ~x537 ;
  assign n5561 = ( x234 & ~x557 ) | ( x234 & n5560 ) | ( ~x557 & n5560 ) ;
  assign n5562 = n5559 | n5561 ;
  assign n5563 = ( x249 & ~x538 ) | ( x249 & n5562 ) | ( ~x538 & n5562 ) ;
  assign n5564 = n5557 & ~n5563 ;
  assign n5565 = n5533 & n5564 ;
  assign n5566 = ~x247 & x516 ;
  assign n5567 = ( ~x234 & x511 ) | ( ~x234 & n5566 ) | ( x511 & n5566 ) ;
  assign n5568 = x247 & ~x516 ;
  assign n5569 = ( x234 & ~x511 ) | ( x234 & n5568 ) | ( ~x511 & n5568 ) ;
  assign n5570 = n5567 | n5569 ;
  assign n5571 = n3535 & n5570 ;
  assign n5572 = ~x245 & x514 ;
  assign n5573 = ( ~x242 & x510 ) | ( ~x242 & n5572 ) | ( x510 & n5572 ) ;
  assign n5574 = x245 & ~x514 ;
  assign n5575 = ( x242 & ~x510 ) | ( x242 & n5574 ) | ( ~x510 & n5574 ) ;
  assign n5576 = n5573 | n5575 ;
  assign n5577 = ~x249 & x579 ;
  assign n5578 = ( ~x240 & x515 ) | ( ~x240 & n5577 ) | ( x515 & n5577 ) ;
  assign n5579 = x249 & ~x579 ;
  assign n5580 = ( x240 & ~x515 ) | ( x240 & n5579 ) | ( ~x515 & n5579 ) ;
  assign n5581 = n5578 | n5580 ;
  assign n5582 = ~x241 & x559 ;
  assign n5583 = ( ~x238 & x517 ) | ( ~x238 & n5582 ) | ( x517 & n5582 ) ;
  assign n5584 = x241 & ~x559 ;
  assign n5585 = ( x238 & ~x517 ) | ( x238 & n5584 ) | ( ~x517 & n5584 ) ;
  assign n5586 = n5583 | n5585 ;
  assign n5587 = ( ~n5576 & n5581 ) | ( ~n5576 & n5586 ) | ( n5581 & n5586 ) ;
  assign n5588 = ~x248 & x481 ;
  assign n5589 = ( ~x246 & x487 ) | ( ~x246 & n5588 ) | ( x487 & n5588 ) ;
  assign n5590 = x248 & ~x481 ;
  assign n5591 = ( x246 & ~x487 ) | ( x246 & n5590 ) | ( ~x487 & n5590 ) ;
  assign n5592 = n5589 | n5591 ;
  assign n5593 = n5576 | n5592 ;
  assign n5594 = n5587 | n5593 ;
  assign n5595 = ( x239 & x488 ) | ( x239 & ~n5594 ) | ( x488 & ~n5594 ) ;
  assign n5596 = ~x244 & x513 ;
  assign n5597 = ( ~x235 & x512 ) | ( ~x235 & n5596 ) | ( x512 & n5596 ) ;
  assign n5598 = x244 & ~x513 ;
  assign n5599 = ( x235 & ~x512 ) | ( x235 & n5598 ) | ( ~x512 & n5598 ) ;
  assign n5600 = n5597 | n5599 ;
  assign n5601 = ( x239 & x488 ) | ( x239 & n5600 ) | ( x488 & n5600 ) ;
  assign n5602 = n5595 & ~n5601 ;
  assign n5603 = n1797 & n5602 ;
  assign n5604 = ( n3535 & n5571 ) | ( n3535 & ~n5603 ) | ( n5571 & ~n5603 ) ;
  assign n5605 = n5565 | n5604 ;
  assign n5606 = ( n5527 & ~n5565 ) | ( n5527 & n5605 ) | ( ~n5565 & n5605 ) ;
  assign n5607 = n5449 & ~n5606 ;
  assign n5608 = ~x806 & x990 ;
  assign n5609 = x600 & n5608 ;
  assign n5610 = ( x332 & x594 ) | ( x332 & n5609 ) | ( x594 & n5609 ) ;
  assign n5611 = ( ~x332 & x594 ) | ( ~x332 & n5609 ) | ( x594 & n5609 ) ;
  assign n5612 = ~n5610 & n5611 ;
  assign n5613 = ~x806 & n4842 ;
  assign n5614 = ( x332 & x595 ) | ( x332 & n5613 ) | ( x595 & n5613 ) ;
  assign n5615 = ( ~x332 & x595 ) | ( ~x332 & n5613 ) | ( x595 & n5613 ) ;
  assign n5616 = ~n5614 & n5615 ;
  assign n5617 = x594 & n5609 ;
  assign n5618 = x595 & x597 ;
  assign n5619 = n5617 & n5618 ;
  assign n5620 = ( x332 & x596 ) | ( x332 & n5619 ) | ( x596 & n5619 ) ;
  assign n5621 = ( ~x332 & x596 ) | ( ~x332 & n5619 ) | ( x596 & n5619 ) ;
  assign n5622 = ~n5620 & n5621 ;
  assign n5623 = ( x332 & x597 ) | ( x332 & n5617 ) | ( x597 & n5617 ) ;
  assign n5624 = ( ~x332 & x597 ) | ( ~x332 & n5617 ) | ( x597 & n5617 ) ;
  assign n5625 = ~n5623 & n5624 ;
  assign n5626 = x882 | n1380 ;
  assign n5627 = x947 & ~n5626 ;
  assign n5628 = x740 & x780 ;
  assign n5629 = n1659 & n5628 ;
  assign n5630 = x598 | n5629 ;
  assign n5631 = ( ~n5627 & n5629 ) | ( ~n5627 & n5630 ) | ( n5629 & n5630 ) ;
  assign n5632 = x596 & n5619 ;
  assign n5633 = ( x332 & x599 ) | ( x332 & n5632 ) | ( x599 & n5632 ) ;
  assign n5634 = ( ~x332 & x599 ) | ( ~x332 & n5632 ) | ( x599 & n5632 ) ;
  assign n5635 = ~n5633 & n5634 ;
  assign n5636 = ( ~x332 & x600 ) | ( ~x332 & n5608 ) | ( x600 & n5608 ) ;
  assign n5637 = ~n5609 & n5636 ;
  assign n5638 = x601 & x806 ;
  assign n5639 = ~x806 & x989 ;
  assign n5640 = ( ~x332 & n5638 ) | ( ~x332 & n5639 ) | ( n5638 & n5639 ) ;
  assign n5641 = ~x230 & x602 ;
  assign n5642 = x230 | x602 ;
  assign n5643 = ( n3219 & n5641 ) | ( n3219 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5644 = ~x871 & x966 ;
  assign n5645 = ~x872 & n5644 ;
  assign n5646 = x1038 & x1060 ;
  assign n5647 = ( x832 & x980 ) | ( x832 & x1061 ) | ( x980 & x1061 ) ;
  assign n5648 = ( x832 & ~n5646 ) | ( x832 & n5647 ) | ( ~n5646 & n5647 ) ;
  assign n5649 = x832 & ~n5648 ;
  assign n5650 = x952 & n5649 ;
  assign n5651 = ~x966 & n5650 ;
  assign n5652 = ( x603 & x966 ) | ( x603 & ~n5651 ) | ( x966 & ~n5651 ) ;
  assign n5653 = x1100 & n5651 ;
  assign n5654 = ( ~n5645 & n5652 ) | ( ~n5645 & n5653 ) | ( n5652 & n5653 ) ;
  assign n5655 = ~x779 & x823 ;
  assign n5656 = ~x299 & x983 ;
  assign n5657 = x604 & ~x907 ;
  assign n5658 = ( x604 & ~n5656 ) | ( x604 & n5657 ) | ( ~n5656 & n5657 ) ;
  assign n5659 = n1655 & ~n5658 ;
  assign n5660 = ( ~x823 & n1655 ) | ( ~x823 & n5658 ) | ( n1655 & n5658 ) ;
  assign n5661 = ( n5655 & ~n5659 ) | ( n5655 & n5660 ) | ( ~n5659 & n5660 ) ;
  assign n5662 = ( x332 & ~x605 ) | ( x332 & x806 ) | ( ~x605 & x806 ) ;
  assign n5663 = ( x332 & x605 ) | ( x332 & ~x806 ) | ( x605 & ~x806 ) ;
  assign n5664 = n5662 | n5663 ;
  assign n5665 = x966 | n5650 ;
  assign n5666 = x837 & x966 ;
  assign n5667 = x606 | n5666 ;
  assign n5668 = ( ~n5665 & n5666 ) | ( ~n5665 & n5667 ) | ( n5666 & n5667 ) ;
  assign n5669 = x1104 & n5651 ;
  assign n5670 = n5668 | n5669 ;
  assign n5671 = x607 & ~n5650 ;
  assign n5672 = x1107 & n5650 ;
  assign n5673 = ( ~x966 & n5671 ) | ( ~x966 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5674 = x608 & ~n5650 ;
  assign n5675 = x1116 & n5650 ;
  assign n5676 = ( ~x966 & n5674 ) | ( ~x966 & n5675 ) | ( n5674 & n5675 ) ;
  assign n5677 = x609 & ~n5650 ;
  assign n5678 = x1118 & n5650 ;
  assign n5679 = ( ~x966 & n5677 ) | ( ~x966 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5680 = x610 & ~n5650 ;
  assign n5681 = x1113 & n5650 ;
  assign n5682 = ( ~x966 & n5680 ) | ( ~x966 & n5681 ) | ( n5680 & n5681 ) ;
  assign n5683 = x611 & ~n5650 ;
  assign n5684 = x1114 & n5650 ;
  assign n5685 = ( ~x966 & n5683 ) | ( ~x966 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5686 = x612 & ~n5650 ;
  assign n5687 = x1111 & n5650 ;
  assign n5688 = ( ~x966 & n5686 ) | ( ~x966 & n5687 ) | ( n5686 & n5687 ) ;
  assign n5689 = x613 & ~n5650 ;
  assign n5690 = x1115 & n5650 ;
  assign n5691 = ( ~x966 & n5689 ) | ( ~x966 & n5690 ) | ( n5689 & n5690 ) ;
  assign n5692 = x1102 & ~n5644 ;
  assign n5693 = ( n5644 & n5651 ) | ( n5644 & ~n5692 ) | ( n5651 & ~n5692 ) ;
  assign n5694 = x614 | n5665 ;
  assign n5695 = ~n5693 & n5694 ;
  assign n5696 = x907 & ~n5626 ;
  assign n5697 = x779 & x797 ;
  assign n5698 = n1656 & n5697 ;
  assign n5699 = x615 & ~n5698 ;
  assign n5700 = ( n5696 & ~n5698 ) | ( n5696 & n5699 ) | ( ~n5698 & n5699 ) ;
  assign n5701 = x616 | n5650 ;
  assign n5702 = x872 & x966 ;
  assign n5703 = ~x1101 & n5650 ;
  assign n5704 = ( x966 & ~n5702 ) | ( x966 & n5703 ) | ( ~n5702 & n5703 ) ;
  assign n5705 = ( n5701 & n5702 ) | ( n5701 & ~n5704 ) | ( n5702 & ~n5704 ) ;
  assign n5706 = x850 & x966 ;
  assign n5707 = x617 | n5706 ;
  assign n5708 = ( ~n5665 & n5706 ) | ( ~n5665 & n5707 ) | ( n5706 & n5707 ) ;
  assign n5709 = x1105 & n5651 ;
  assign n5710 = n5708 | n5709 ;
  assign n5711 = x618 & ~n5650 ;
  assign n5712 = x1117 & n5650 ;
  assign n5713 = ( ~x966 & n5711 ) | ( ~x966 & n5712 ) | ( n5711 & n5712 ) ;
  assign n5714 = x619 & ~n5650 ;
  assign n5715 = x1122 & n5650 ;
  assign n5716 = ( ~x966 & n5714 ) | ( ~x966 & n5715 ) | ( n5714 & n5715 ) ;
  assign n5717 = x620 & ~n5650 ;
  assign n5718 = x1112 & n5650 ;
  assign n5719 = ( ~x966 & n5717 ) | ( ~x966 & n5718 ) | ( n5717 & n5718 ) ;
  assign n5720 = x621 & ~n5650 ;
  assign n5721 = x1108 & n5650 ;
  assign n5722 = ( ~x966 & n5720 ) | ( ~x966 & n5721 ) | ( n5720 & n5721 ) ;
  assign n5723 = x622 & ~n5650 ;
  assign n5724 = x1109 & n5650 ;
  assign n5725 = ( ~x966 & n5723 ) | ( ~x966 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5726 = x623 & ~n5650 ;
  assign n5727 = x1106 & n5650 ;
  assign n5728 = ( ~x966 & n5726 ) | ( ~x966 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5729 = ~x780 & x831 ;
  assign n5730 = x624 & ~x947 ;
  assign n5731 = ( x624 & ~n5656 ) | ( x624 & n5730 ) | ( ~n5656 & n5730 ) ;
  assign n5732 = n1658 & ~n5731 ;
  assign n5733 = ( ~x831 & n1658 ) | ( ~x831 & n5731 ) | ( n1658 & n5731 ) ;
  assign n5734 = ( n5729 & ~n5732 ) | ( n5729 & n5733 ) | ( ~n5732 & n5733 ) ;
  assign n5735 = ~x1054 & x1066 ;
  assign n5736 = ( x832 & x973 ) | ( x832 & ~x1088 ) | ( x973 & ~x1088 ) ;
  assign n5737 = ( x832 & ~n5735 ) | ( x832 & n5736 ) | ( ~n5735 & n5736 ) ;
  assign n5738 = x832 & ~n5737 ;
  assign n5739 = ~x953 & n5738 ;
  assign n5740 = x625 & ~n5739 ;
  assign n5741 = x1116 & n5739 ;
  assign n5742 = ( ~x962 & n5740 ) | ( ~x962 & n5741 ) | ( n5740 & n5741 ) ;
  assign n5743 = x626 & ~n5650 ;
  assign n5744 = x1121 & n5650 ;
  assign n5745 = ( ~x966 & n5743 ) | ( ~x966 & n5744 ) | ( n5743 & n5744 ) ;
  assign n5746 = x627 & ~n5739 ;
  assign n5747 = x1117 & n5739 ;
  assign n5748 = ( ~x962 & n5746 ) | ( ~x962 & n5747 ) | ( n5746 & n5747 ) ;
  assign n5749 = x628 & ~n5739 ;
  assign n5750 = x1119 & n5739 ;
  assign n5751 = ( ~x962 & n5749 ) | ( ~x962 & n5750 ) | ( n5749 & n5750 ) ;
  assign n5752 = x629 & ~n5650 ;
  assign n5753 = x1119 & n5650 ;
  assign n5754 = ( ~x966 & n5752 ) | ( ~x966 & n5753 ) | ( n5752 & n5753 ) ;
  assign n5755 = x630 & ~n5650 ;
  assign n5756 = x1120 & n5650 ;
  assign n5757 = ( ~x966 & n5755 ) | ( ~x966 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5758 = x631 | n5739 ;
  assign n5759 = x1113 & n5739 ;
  assign n5760 = ( x962 & n5758 ) | ( x962 & ~n5759 ) | ( n5758 & ~n5759 ) ;
  assign n5761 = x632 | n5739 ;
  assign n5762 = x1115 & n5739 ;
  assign n5763 = ( x962 & n5761 ) | ( x962 & ~n5762 ) | ( n5761 & ~n5762 ) ;
  assign n5764 = x633 & ~n5650 ;
  assign n5765 = x1110 & n5650 ;
  assign n5766 = ( ~x966 & n5764 ) | ( ~x966 & n5765 ) | ( n5764 & n5765 ) ;
  assign n5767 = x634 & ~n5739 ;
  assign n5768 = x1110 & n5739 ;
  assign n5769 = ( ~x962 & n5767 ) | ( ~x962 & n5768 ) | ( n5767 & n5768 ) ;
  assign n5770 = x635 | n5739 ;
  assign n5771 = x1112 & n5739 ;
  assign n5772 = ( x962 & n5770 ) | ( x962 & ~n5771 ) | ( n5770 & ~n5771 ) ;
  assign n5773 = x636 & ~n5650 ;
  assign n5774 = x1127 & n5650 ;
  assign n5775 = ( ~x966 & n5773 ) | ( ~x966 & n5774 ) | ( n5773 & n5774 ) ;
  assign n5776 = x637 & ~n5739 ;
  assign n5777 = x1105 & n5739 ;
  assign n5778 = ( ~x962 & n5776 ) | ( ~x962 & n5777 ) | ( n5776 & n5777 ) ;
  assign n5779 = x638 & ~n5739 ;
  assign n5780 = x1107 & n5739 ;
  assign n5781 = ( ~x962 & n5779 ) | ( ~x962 & n5780 ) | ( n5779 & n5780 ) ;
  assign n5782 = x639 & ~n5739 ;
  assign n5783 = x1109 & n5739 ;
  assign n5784 = ( ~x962 & n5782 ) | ( ~x962 & n5783 ) | ( n5782 & n5783 ) ;
  assign n5785 = x640 & ~n5650 ;
  assign n5786 = x1128 & n5650 ;
  assign n5787 = ( ~x966 & n5785 ) | ( ~x966 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5788 = x641 & ~n5739 ;
  assign n5789 = x1121 & n5739 ;
  assign n5790 = ( ~x962 & n5788 ) | ( ~x962 & n5789 ) | ( n5788 & n5789 ) ;
  assign n5791 = x642 & ~n5650 ;
  assign n5792 = x1103 & n5650 ;
  assign n5793 = ( ~x966 & n5791 ) | ( ~x966 & n5792 ) | ( n5791 & n5792 ) ;
  assign n5794 = x643 & ~n5739 ;
  assign n5795 = x1104 & n5739 ;
  assign n5796 = ( ~x962 & n5794 ) | ( ~x962 & n5795 ) | ( n5794 & n5795 ) ;
  assign n5797 = x644 & ~n5650 ;
  assign n5798 = x1123 & n5650 ;
  assign n5799 = ( ~x966 & n5797 ) | ( ~x966 & n5798 ) | ( n5797 & n5798 ) ;
  assign n5800 = x645 & ~n5650 ;
  assign n5801 = x1125 & n5650 ;
  assign n5802 = ( ~x966 & n5800 ) | ( ~x966 & n5801 ) | ( n5800 & n5801 ) ;
  assign n5803 = x646 | n5739 ;
  assign n5804 = x1114 & n5739 ;
  assign n5805 = ( x962 & n5803 ) | ( x962 & ~n5804 ) | ( n5803 & ~n5804 ) ;
  assign n5806 = x647 & ~n5739 ;
  assign n5807 = x1120 & n5739 ;
  assign n5808 = ( ~x962 & n5806 ) | ( ~x962 & n5807 ) | ( n5806 & n5807 ) ;
  assign n5809 = x648 & ~n5739 ;
  assign n5810 = x1122 & n5739 ;
  assign n5811 = ( ~x962 & n5809 ) | ( ~x962 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5812 = x649 | n5739 ;
  assign n5813 = x1126 & n5739 ;
  assign n5814 = ( x962 & n5812 ) | ( x962 & ~n5813 ) | ( n5812 & ~n5813 ) ;
  assign n5815 = x650 | n5739 ;
  assign n5816 = x1127 & n5739 ;
  assign n5817 = ( x962 & n5815 ) | ( x962 & ~n5816 ) | ( n5815 & ~n5816 ) ;
  assign n5818 = x651 & ~n5650 ;
  assign n5819 = x1130 & n5650 ;
  assign n5820 = ( ~x966 & n5818 ) | ( ~x966 & n5819 ) | ( n5818 & n5819 ) ;
  assign n5821 = x652 & ~n5650 ;
  assign n5822 = x1131 & n5650 ;
  assign n5823 = ( ~x966 & n5821 ) | ( ~x966 & n5822 ) | ( n5821 & n5822 ) ;
  assign n5824 = x653 & ~n5650 ;
  assign n5825 = x1129 & n5650 ;
  assign n5826 = ( ~x966 & n5824 ) | ( ~x966 & n5825 ) | ( n5824 & n5825 ) ;
  assign n5827 = x654 | n5739 ;
  assign n5828 = x1130 & n5739 ;
  assign n5829 = ( x962 & n5827 ) | ( x962 & ~n5828 ) | ( n5827 & ~n5828 ) ;
  assign n5830 = x655 | n5739 ;
  assign n5831 = x1124 & n5739 ;
  assign n5832 = ( x962 & n5830 ) | ( x962 & ~n5831 ) | ( n5830 & ~n5831 ) ;
  assign n5833 = x656 & ~n5650 ;
  assign n5834 = x1126 & n5650 ;
  assign n5835 = ( ~x966 & n5833 ) | ( ~x966 & n5834 ) | ( n5833 & n5834 ) ;
  assign n5836 = x657 | n5739 ;
  assign n5837 = x1131 & n5739 ;
  assign n5838 = ( x962 & n5836 ) | ( x962 & ~n5837 ) | ( n5836 & ~n5837 ) ;
  assign n5839 = x658 & ~n5650 ;
  assign n5840 = x1124 & n5650 ;
  assign n5841 = ( ~x966 & n5839 ) | ( ~x966 & n5840 ) | ( n5839 & n5840 ) ;
  assign n5842 = x266 & x992 ;
  assign n5843 = ~x280 & n5842 ;
  assign n5844 = ~x269 & n5843 ;
  assign n5845 = x270 | x277 ;
  assign n5846 = x281 | x282 ;
  assign n5847 = n5845 | n5846 ;
  assign n5848 = x264 | n5847 ;
  assign n5849 = n5844 & ~n5848 ;
  assign n5850 = ~x265 & n5849 ;
  assign n5851 = ~x274 & n5850 ;
  assign n5852 = x274 & ~n5850 ;
  assign n5853 = n5851 | n5852 ;
  assign n5854 = x660 & ~n5739 ;
  assign n5855 = x1118 & n5739 ;
  assign n5856 = ( ~x962 & n5854 ) | ( ~x962 & n5855 ) | ( n5854 & n5855 ) ;
  assign n5857 = x661 & ~n5739 ;
  assign n5858 = x1101 & n5739 ;
  assign n5859 = ( ~x962 & n5857 ) | ( ~x962 & n5858 ) | ( n5857 & n5858 ) ;
  assign n5860 = x662 & ~n5739 ;
  assign n5861 = x1102 & n5739 ;
  assign n5862 = ( ~x962 & n5860 ) | ( ~x962 & n5861 ) | ( n5860 & n5861 ) ;
  assign n5863 = x1137 | x1138 ;
  assign n5864 = n2144 & ~n5863 ;
  assign n5865 = ~x1134 & n5864 ;
  assign n5866 = x1135 & ~x1136 ;
  assign n5867 = n5865 & n5866 ;
  assign n5868 = x784 & n5867 ;
  assign n5869 = ~x1135 & x1136 ;
  assign n5870 = x1134 & n5864 ;
  assign n5871 = n5869 & n5870 ;
  assign n5872 = x766 & n5871 ;
  assign n5873 = n5868 | n5872 ;
  assign n5874 = x1135 & x1136 ;
  assign n5875 = n5870 & n5874 ;
  assign n5876 = x700 & n5875 ;
  assign n5877 = n1499 | n2144 ;
  assign n5878 = n1881 | n5877 ;
  assign n5879 = n1945 & ~n5878 ;
  assign n5880 = x334 & n5879 ;
  assign n5881 = n5876 | n5880 ;
  assign n5882 = x1135 | x1136 ;
  assign n5883 = n5870 & ~n5882 ;
  assign n5884 = x855 & n5883 ;
  assign n5885 = ( ~n5873 & n5881 ) | ( ~n5873 & n5884 ) | ( n5881 & n5884 ) ;
  assign n5886 = n5865 & ~n5882 ;
  assign n5887 = x815 & n5886 ;
  assign n5888 = n5873 | n5887 ;
  assign n5889 = n5885 | n5888 ;
  assign n5890 = n2136 & ~n5877 ;
  assign n5891 = x365 & n5890 ;
  assign n5892 = n2013 & ~n5877 ;
  assign n5893 = x323 & n5892 ;
  assign n5894 = n5891 | n5893 ;
  assign n5895 = n1882 & ~n5878 ;
  assign n5896 = x199 & x1065 ;
  assign n5897 = n1499 & ~n2144 ;
  assign n5898 = ~x199 & x257 ;
  assign n5899 = ( n5896 & n5897 ) | ( n5896 & n5898 ) | ( n5897 & n5898 ) ;
  assign n5900 = x464 | n5899 ;
  assign n5901 = ( n5895 & n5899 ) | ( n5895 & n5900 ) | ( n5899 & n5900 ) ;
  assign n5902 = n5894 | n5901 ;
  assign n5903 = n5865 & n5869 ;
  assign n5904 = x633 & n5903 ;
  assign n5905 = n5865 & n5874 ;
  assign n5906 = x634 & ~n5905 ;
  assign n5907 = ( x634 & n5904 ) | ( x634 & ~n5906 ) | ( n5904 & ~n5906 ) ;
  assign n5908 = n5902 | n5907 ;
  assign n5909 = n5889 | n5908 ;
  assign n5910 = x727 & n5875 ;
  assign n5911 = ~x662 & x1135 ;
  assign n5912 = x614 | x1135 ;
  assign n5913 = ( x1136 & n5911 ) | ( x1136 & ~n5912 ) | ( n5911 & ~n5912 ) ;
  assign n5914 = x811 | x1135 ;
  assign n5915 = ~x785 & x1135 ;
  assign n5916 = ( x1136 & n5914 ) | ( x1136 & ~n5915 ) | ( n5914 & ~n5915 ) ;
  assign n5917 = ~n5913 & n5916 ;
  assign n5918 = n5865 & n5917 ;
  assign n5919 = ~x355 & n5892 ;
  assign n5920 = ( n5892 & n5918 ) | ( n5892 & ~n5919 ) | ( n5918 & ~n5919 ) ;
  assign n5921 = x199 & x1084 ;
  assign n5922 = ~x199 & x292 ;
  assign n5923 = ( n5897 & n5921 ) | ( n5897 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5924 = x872 | n5923 ;
  assign n5925 = ( n5883 & n5923 ) | ( n5883 & n5924 ) | ( n5923 & n5924 ) ;
  assign n5926 = ( ~n5910 & n5920 ) | ( ~n5910 & n5925 ) | ( n5920 & n5925 ) ;
  assign n5927 = x380 & n5890 ;
  assign n5928 = n5910 | n5927 ;
  assign n5929 = n5926 | n5928 ;
  assign n5930 = x429 & n5895 ;
  assign n5931 = x404 & n5879 ;
  assign n5932 = x772 & n5871 ;
  assign n5933 = ( ~n5930 & n5931 ) | ( ~n5930 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5934 = n5930 | n5933 ;
  assign n5935 = n5929 | n5934 ;
  assign n5936 = x665 & ~n5739 ;
  assign n5937 = x1108 & n5739 ;
  assign n5938 = ( ~x962 & n5936 ) | ( ~x962 & n5937 ) | ( n5936 & n5937 ) ;
  assign n5939 = x199 & x1044 ;
  assign n5940 = ~x199 & x297 ;
  assign n5941 = ( n5897 & n5939 ) | ( n5897 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5942 = x441 & n5892 ;
  assign n5943 = n5941 | n5942 ;
  assign n5944 = x764 & n5871 ;
  assign n5945 = x443 & n5895 ;
  assign n5946 = ( ~n5943 & n5944 ) | ( ~n5943 & n5945 ) | ( n5944 & n5945 ) ;
  assign n5947 = n5943 | n5946 ;
  assign n5948 = x691 & n5875 ;
  assign n5949 = x873 & n5883 ;
  assign n5950 = n5948 | n5949 ;
  assign n5951 = ~x790 & n5866 ;
  assign n5952 = x799 & ~n5882 ;
  assign n5953 = ~x638 & n5874 ;
  assign n5954 = ( ~n5951 & n5952 ) | ( ~n5951 & n5953 ) | ( n5952 & n5953 ) ;
  assign n5955 = ~x607 & n5869 ;
  assign n5956 = n5951 | n5955 ;
  assign n5957 = n5954 | n5956 ;
  assign n5958 = n5865 & ~n5957 ;
  assign n5959 = ~x337 & n5890 ;
  assign n5960 = ( n5890 & n5958 ) | ( n5890 & ~n5959 ) | ( n5958 & ~n5959 ) ;
  assign n5961 = x456 & n5879 ;
  assign n5962 = ( ~n5950 & n5960 ) | ( ~n5950 & n5961 ) | ( n5960 & n5961 ) ;
  assign n5963 = n5950 | n5962 ;
  assign n5964 = n5947 | n5963 ;
  assign n5965 = x199 & n5897 ;
  assign n5966 = x1072 & n5965 ;
  assign n5967 = ~x871 & n5883 ;
  assign n5968 = ( n5883 & n5966 ) | ( n5883 & ~n5967 ) | ( n5966 & ~n5967 ) ;
  assign n5969 = x699 & n5875 ;
  assign n5970 = x763 & n5871 ;
  assign n5971 = x444 & n5895 ;
  assign n5972 = ( ~n5969 & n5970 ) | ( ~n5969 & n5971 ) | ( n5970 & n5971 ) ;
  assign n5973 = x319 & n5879 ;
  assign n5974 = n5969 | n5973 ;
  assign n5975 = n5972 | n5974 ;
  assign n5976 = x792 & ~x1136 ;
  assign n5977 = x681 & x1136 ;
  assign n5978 = ( x1135 & n5976 ) | ( x1135 & n5977 ) | ( n5976 & n5977 ) ;
  assign n5979 = x809 | x1136 ;
  assign n5980 = x642 & x1136 ;
  assign n5981 = ( x1135 & n5979 ) | ( x1135 & ~n5980 ) | ( n5979 & ~n5980 ) ;
  assign n5982 = ~n5978 & n5981 ;
  assign n5983 = n5865 & ~n5982 ;
  assign n5984 = ~x338 & n5890 ;
  assign n5985 = ( n5890 & n5983 ) | ( n5890 & ~n5984 ) | ( n5983 & ~n5984 ) ;
  assign n5986 = x458 & n5892 ;
  assign n5987 = ~x199 & n5897 ;
  assign n5988 = x294 & n5987 ;
  assign n5989 = ( ~n5985 & n5986 ) | ( ~n5985 & n5988 ) | ( n5986 & n5988 ) ;
  assign n5990 = n5985 | n5989 ;
  assign n5991 = ( ~n5968 & n5975 ) | ( ~n5968 & n5990 ) | ( n5975 & n5990 ) ;
  assign n5992 = n5968 | n5991 ;
  assign n5993 = x363 & n5890 ;
  assign n5994 = x291 & n5987 ;
  assign n5995 = x342 & n5892 ;
  assign n5996 = ( ~n5993 & n5994 ) | ( ~n5993 & n5995 ) | ( n5994 & n5995 ) ;
  assign n5997 = n5993 | n5996 ;
  assign n5998 = x981 & ~x1136 ;
  assign n5999 = x603 & x1136 ;
  assign n6000 = ( ~x1135 & n5998 ) | ( ~x1135 & n5999 ) | ( n5998 & n5999 ) ;
  assign n6001 = x778 & ~x1136 ;
  assign n6002 = x680 & x1136 ;
  assign n6003 = ( x1135 & n6001 ) | ( x1135 & n6002 ) | ( n6001 & n6002 ) ;
  assign n6004 = n6000 | n6003 ;
  assign n6005 = n5865 & n6004 ;
  assign n6006 = ~x1049 & n5965 ;
  assign n6007 = ( n5965 & n6005 ) | ( n5965 & ~n6006 ) | ( n6005 & ~n6006 ) ;
  assign n6008 = x837 & n5883 ;
  assign n6009 = ( ~n5997 & n6007 ) | ( ~n5997 & n6008 ) | ( n6007 & n6008 ) ;
  assign n6010 = n5997 | n6009 ;
  assign n6011 = x414 & n5895 ;
  assign n6012 = x759 & n5871 ;
  assign n6013 = x696 & n5875 ;
  assign n6014 = ( ~n6011 & n6012 ) | ( ~n6011 & n6013 ) | ( n6012 & n6013 ) ;
  assign n6015 = x390 & n5879 ;
  assign n6016 = n6011 | n6015 ;
  assign n6017 = n6014 | n6016 ;
  assign n6018 = n6010 | n6017 ;
  assign n6019 = x669 | n5739 ;
  assign n6020 = x1125 & n5739 ;
  assign n6021 = ( x962 & n6019 ) | ( x962 & ~n6020 ) | ( n6019 & ~n6020 ) ;
  assign n6022 = x364 & n5890 ;
  assign n6023 = x1062 & n5965 ;
  assign n6024 = x343 & n5892 ;
  assign n6025 = ( ~n6022 & n6023 ) | ( ~n6022 & n6024 ) | ( n6023 & n6024 ) ;
  assign n6026 = x258 & n5987 ;
  assign n6027 = n6022 | n6026 ;
  assign n6028 = n6025 | n6027 ;
  assign n6029 = x852 & n5883 ;
  assign n6030 = ~x695 & n5905 ;
  assign n6031 = ( ~n6028 & n6029 ) | ( ~n6028 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6032 = n6028 | n6031 ;
  assign n6033 = x391 & n5879 ;
  assign n6034 = x612 & n5903 ;
  assign n6035 = ( ~n6028 & n6033 ) | ( ~n6028 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6036 = ~x745 & n5871 ;
  assign n6037 = ~x723 & n5875 ;
  assign n6038 = x415 & n5895 ;
  assign n6039 = ( ~n6036 & n6037 ) | ( ~n6036 & n6038 ) | ( n6037 & n6038 ) ;
  assign n6040 = n6036 | n6039 ;
  assign n6041 = n6035 | n6040 ;
  assign n6042 = n6032 | n6041 ;
  assign n6043 = x447 & n5890 ;
  assign n6044 = x1040 & n5965 ;
  assign n6045 = x327 & n5892 ;
  assign n6046 = ( ~n6043 & n6044 ) | ( ~n6043 & n6045 ) | ( n6044 & n6045 ) ;
  assign n6047 = x261 & n5987 ;
  assign n6048 = n6043 | n6047 ;
  assign n6049 = n6046 | n6048 ;
  assign n6050 = x333 & n5879 ;
  assign n6051 = n6049 | n6050 ;
  assign n6052 = x865 & n5883 ;
  assign n6053 = ~x724 & n5875 ;
  assign n6054 = ~x741 & n5871 ;
  assign n6055 = ( ~n6052 & n6053 ) | ( ~n6052 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6056 = n6052 | n6055 ;
  assign n6057 = x611 & n5903 ;
  assign n6058 = x453 & n5895 ;
  assign n6059 = ~x646 & n5905 ;
  assign n6060 = ( ~n6057 & n6058 ) | ( ~n6057 & n6059 ) | ( n6058 & n6059 ) ;
  assign n6061 = n6057 | n6060 ;
  assign n6062 = ( ~n6051 & n6056 ) | ( ~n6051 & n6061 ) | ( n6056 & n6061 ) ;
  assign n6063 = n6051 | n6062 ;
  assign n6064 = x1048 & n5965 ;
  assign n6065 = x422 & n5895 ;
  assign n6066 = x758 & n5871 ;
  assign n6067 = ( ~n6064 & n6065 ) | ( ~n6064 & n6066 ) | ( n6065 & n6066 ) ;
  assign n6068 = n6064 | n6067 ;
  assign n6069 = x850 & n5883 ;
  assign n6070 = x397 & n5879 ;
  assign n6071 = x736 & n5875 ;
  assign n6072 = ( ~n6069 & n6070 ) | ( ~n6069 & n6071 ) | ( n6070 & n6071 ) ;
  assign n6073 = n6069 | n6072 ;
  assign n6074 = x808 | x1136 ;
  assign n6075 = ~x616 & x1136 ;
  assign n6076 = ( x1135 & n6074 ) | ( x1135 & ~n6075 ) | ( n6074 & ~n6075 ) ;
  assign n6077 = x781 | x1136 ;
  assign n6078 = ~x661 & x1136 ;
  assign n6079 = ( x1135 & ~n6077 ) | ( x1135 & n6078 ) | ( ~n6077 & n6078 ) ;
  assign n6080 = n6076 & ~n6079 ;
  assign n6081 = n5865 & n6080 ;
  assign n6082 = ~x372 & n5890 ;
  assign n6083 = ( n5890 & n6081 ) | ( n5890 & ~n6082 ) | ( n6081 & ~n6082 ) ;
  assign n6084 = x290 & n5987 ;
  assign n6085 = x320 & n5892 ;
  assign n6086 = ( ~n6083 & n6084 ) | ( ~n6083 & n6085 ) | ( n6084 & n6085 ) ;
  assign n6087 = n6083 | n6086 ;
  assign n6088 = ( ~n6068 & n6073 ) | ( ~n6068 & n6087 ) | ( n6073 & n6087 ) ;
  assign n6089 = n6068 | n6088 ;
  assign n6090 = x1053 & n5965 ;
  assign n6091 = x452 & n5892 ;
  assign n6092 = x295 & n5987 ;
  assign n6093 = ( ~n6090 & n6091 ) | ( ~n6090 & n6092 ) | ( n6091 & n6092 ) ;
  assign n6094 = x387 & n5890 ;
  assign n6095 = n6090 | n6094 ;
  assign n6096 = n6093 | n6095 ;
  assign n6097 = x866 & n5883 ;
  assign n6098 = x617 & n5903 ;
  assign n6099 = ( ~n6096 & n6097 ) | ( ~n6096 & n6098 ) | ( n6097 & n6098 ) ;
  assign n6100 = n6096 | n6099 ;
  assign n6101 = x435 & n5895 ;
  assign n6102 = x788 & n5867 ;
  assign n6103 = x749 & n5871 ;
  assign n6104 = ( ~n6101 & n6102 ) | ( ~n6101 & n6103 ) | ( n6102 & n6103 ) ;
  assign n6105 = x411 & n5879 ;
  assign n6106 = n6101 | n6105 ;
  assign n6107 = n6104 | n6106 ;
  assign n6108 = ~x814 & n5886 ;
  assign n6109 = x637 & n5905 ;
  assign n6110 = x706 & n5875 ;
  assign n6111 = ( ~n6108 & n6109 ) | ( ~n6108 & n6110 ) | ( n6109 & n6110 ) ;
  assign n6112 = n6108 | n6111 ;
  assign n6113 = n6107 | n6112 ;
  assign n6114 = n6100 | n6113 ;
  assign n6115 = x437 & n5895 ;
  assign n6116 = x362 & n5892 ;
  assign n6117 = x735 & n5875 ;
  assign n6118 = ( ~n6115 & n6116 ) | ( ~n6115 & n6117 ) | ( n6116 & n6117 ) ;
  assign n6119 = n6115 | n6118 ;
  assign n6120 = x743 & n5871 ;
  assign n6121 = x463 & n5879 ;
  assign n6122 = x859 & n5883 ;
  assign n6123 = ( ~n6120 & n6121 ) | ( ~n6120 & n6122 ) | ( n6121 & n6122 ) ;
  assign n6124 = n6120 | n6123 ;
  assign n6125 = x804 | x1136 ;
  assign n6126 = ~x622 & x1136 ;
  assign n6127 = ( x1135 & n6125 ) | ( x1135 & ~n6126 ) | ( n6125 & ~n6126 ) ;
  assign n6128 = x783 | x1136 ;
  assign n6129 = ~x639 & x1136 ;
  assign n6130 = ( x1135 & ~n6128 ) | ( x1135 & n6129 ) | ( ~n6128 & n6129 ) ;
  assign n6131 = n6127 & ~n6130 ;
  assign n6132 = n5865 & n6131 ;
  assign n6133 = ~x256 & n5987 ;
  assign n6134 = ( n5987 & n6132 ) | ( n5987 & ~n6133 ) | ( n6132 & ~n6133 ) ;
  assign n6135 = x336 & n5890 ;
  assign n6136 = x1070 & n5965 ;
  assign n6137 = ( ~n6134 & n6135 ) | ( ~n6134 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = n6134 | n6137 ;
  assign n6139 = ( ~n6119 & n6124 ) | ( ~n6119 & n6138 ) | ( n6124 & n6138 ) ;
  assign n6140 = n6119 | n6139 ;
  assign n6141 = x876 & n5883 ;
  assign n6142 = x710 & n5905 ;
  assign n6143 = n6141 | n6142 ;
  assign n6144 = x1037 & n5965 ;
  assign n6145 = x455 & n5892 ;
  assign n6146 = x296 & n5987 ;
  assign n6147 = ( ~n6144 & n6145 ) | ( ~n6144 & n6146 ) | ( n6145 & n6146 ) ;
  assign n6148 = x388 & n5890 ;
  assign n6149 = n6144 | n6148 ;
  assign n6150 = n6147 | n6149 ;
  assign n6151 = ~x803 & n5886 ;
  assign n6152 = ( ~n6143 & n6150 ) | ( ~n6143 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6153 = n6143 | n6152 ;
  assign n6154 = x436 & n5895 ;
  assign n6155 = x412 & n5879 ;
  assign n6156 = x748 & n5871 ;
  assign n6157 = ( ~n6154 & n6155 ) | ( ~n6154 & n6156 ) | ( n6155 & n6156 ) ;
  assign n6158 = n6154 | n6157 ;
  assign n6159 = x623 & n5903 ;
  assign n6160 = x730 & n5875 ;
  assign n6161 = x789 & n5867 ;
  assign n6162 = ( ~n6159 & n6160 ) | ( ~n6159 & n6161 ) | ( n6160 & n6161 ) ;
  assign n6163 = n6159 | n6162 ;
  assign n6164 = n6158 | n6163 ;
  assign n6165 = n6153 | n6164 ;
  assign n6166 = x1059 & n5965 ;
  assign n6167 = x386 & n5890 ;
  assign n6168 = x293 & n5987 ;
  assign n6169 = ( ~n6166 & n6167 ) | ( ~n6166 & n6168 ) | ( n6167 & n6168 ) ;
  assign n6170 = x361 & n5892 ;
  assign n6171 = n6166 | n6170 ;
  assign n6172 = n6169 | n6171 ;
  assign n6173 = x787 & n5867 ;
  assign n6174 = x746 & n5871 ;
  assign n6175 = ( ~n6172 & n6173 ) | ( ~n6172 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6176 = n6172 | n6175 ;
  assign n6177 = x881 & n5883 ;
  assign n6178 = x606 & n5903 ;
  assign n6179 = x434 & n5895 ;
  assign n6180 = ( ~n6177 & n6178 ) | ( ~n6177 & n6179 ) | ( n6178 & n6179 ) ;
  assign n6181 = x410 & n5879 ;
  assign n6182 = n6177 | n6181 ;
  assign n6183 = n6180 | n6182 ;
  assign n6184 = ~x812 & n5886 ;
  assign n6185 = x729 & n5875 ;
  assign n6186 = x643 & n5905 ;
  assign n6187 = ( ~n6184 & n6185 ) | ( ~n6184 & n6186 ) | ( n6185 & n6186 ) ;
  assign n6188 = n6184 | n6187 ;
  assign n6189 = n6183 | n6188 ;
  assign n6190 = n6176 | n6189 ;
  assign n6191 = x366 & n5890 ;
  assign n6192 = x1069 & n5965 ;
  assign n6193 = x344 & n5892 ;
  assign n6194 = ( ~n6191 & n6192 ) | ( ~n6191 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6195 = x259 & n5987 ;
  assign n6196 = n6191 | n6195 ;
  assign n6197 = n6194 | n6196 ;
  assign n6198 = x620 & n5903 ;
  assign n6199 = x416 & n5895 ;
  assign n6200 = ( ~n6197 & n6198 ) | ( ~n6197 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = n6197 | n6200 ;
  assign n6202 = ~x635 & n5905 ;
  assign n6203 = ~x704 & n5875 ;
  assign n6204 = ( ~n6197 & n6202 ) | ( ~n6197 & n6203 ) | ( n6202 & n6203 ) ;
  assign n6205 = ~x742 & n5871 ;
  assign n6206 = x335 & n5879 ;
  assign n6207 = x870 & n5883 ;
  assign n6208 = ( ~n6205 & n6206 ) | ( ~n6205 & n6207 ) | ( n6206 & n6207 ) ;
  assign n6209 = n6205 | n6208 ;
  assign n6210 = n6204 | n6209 ;
  assign n6211 = n6201 | n6210 ;
  assign n6212 = x346 & n5892 ;
  assign n6213 = x1067 & n5965 ;
  assign n6214 = x368 & n5890 ;
  assign n6215 = ( ~n6212 & n6213 ) | ( ~n6212 & n6214 ) | ( n6213 & n6214 ) ;
  assign n6216 = x260 & n5987 ;
  assign n6217 = n6212 | n6216 ;
  assign n6218 = n6215 | n6217 ;
  assign n6219 = ~x760 & n5871 ;
  assign n6220 = x613 & n5903 ;
  assign n6221 = ( ~n6218 & n6219 ) | ( ~n6218 & n6220 ) | ( n6219 & n6220 ) ;
  assign n6222 = n6218 | n6221 ;
  assign n6223 = x393 & n5879 ;
  assign n6224 = ~x632 & n5905 ;
  assign n6225 = ( ~n6218 & n6223 ) | ( ~n6218 & n6224 ) | ( n6223 & n6224 ) ;
  assign n6226 = ~x688 & n5875 ;
  assign n6227 = x418 & n5895 ;
  assign n6228 = x856 & n5883 ;
  assign n6229 = ( ~n6226 & n6227 ) | ( ~n6226 & n6228 ) | ( n6227 & n6228 ) ;
  assign n6230 = n6226 | n6229 ;
  assign n6231 = n6225 | n6230 ;
  assign n6232 = n6222 | n6231 ;
  assign n6233 = x450 & n5892 ;
  assign n6234 = x199 & x1036 ;
  assign n6235 = ~x199 & x255 ;
  assign n6236 = ( n5897 & n6234 ) | ( n5897 & n6235 ) | ( n6234 & n6235 ) ;
  assign n6237 = x810 | x1136 ;
  assign n6238 = ~x621 & x1136 ;
  assign n6239 = ( x1135 & n6237 ) | ( x1135 & ~n6238 ) | ( n6237 & ~n6238 ) ;
  assign n6240 = x791 | x1136 ;
  assign n6241 = ~x665 & x1136 ;
  assign n6242 = ( x1135 & ~n6240 ) | ( x1135 & n6241 ) | ( ~n6240 & n6241 ) ;
  assign n6243 = n6239 & ~n6242 ;
  assign n6244 = n5865 & n6243 ;
  assign n6245 = ( ~n6233 & n6236 ) | ( ~n6233 & n6244 ) | ( n6236 & n6244 ) ;
  assign n6246 = n6233 | n6245 ;
  assign n6247 = x438 & n5895 ;
  assign n6248 = x389 & n5890 ;
  assign n6249 = ( ~n6246 & n6247 ) | ( ~n6246 & n6248 ) | ( n6247 & n6248 ) ;
  assign n6250 = n6246 | n6249 ;
  assign n6251 = x874 & n5883 ;
  assign n6252 = x739 & n5871 ;
  assign n6253 = x690 & n5875 ;
  assign n6254 = ( ~n6251 & n6252 ) | ( ~n6251 & n6253 ) | ( n6252 & n6253 ) ;
  assign n6255 = x413 & n5879 ;
  assign n6256 = n6251 | n6255 ;
  assign n6257 = n6254 | n6256 ;
  assign n6258 = n6250 | n6257 ;
  assign n6259 = x680 & ~n5739 ;
  assign n6260 = x1100 & n5739 ;
  assign n6261 = ( ~x962 & n6259 ) | ( ~x962 & n6260 ) | ( n6259 & n6260 ) ;
  assign n6262 = x681 & ~n5739 ;
  assign n6263 = x1103 & n5739 ;
  assign n6264 = ( ~x962 & n6262 ) | ( ~x962 & n6263 ) | ( n6262 & n6263 ) ;
  assign n6265 = x367 & n5890 ;
  assign n6266 = x1039 & n5965 ;
  assign n6267 = x345 & n5892 ;
  assign n6268 = ( ~n6265 & n6266 ) | ( ~n6265 & n6267 ) | ( n6266 & n6267 ) ;
  assign n6269 = x251 & n5987 ;
  assign n6270 = n6265 | n6269 ;
  assign n6271 = n6268 | n6270 ;
  assign n6272 = ~x686 & n5875 ;
  assign n6273 = x610 & n5903 ;
  assign n6274 = ( ~n6271 & n6272 ) | ( ~n6271 & n6273 ) | ( n6272 & n6273 ) ;
  assign n6275 = n6271 | n6274 ;
  assign n6276 = x392 & n5879 ;
  assign n6277 = ~x757 & n5871 ;
  assign n6278 = ( ~n6271 & n6276 ) | ( ~n6271 & n6277 ) | ( n6276 & n6277 ) ;
  assign n6279 = x848 & n5883 ;
  assign n6280 = x417 & n5895 ;
  assign n6281 = ~x631 & n5905 ;
  assign n6282 = ( ~n6279 & n6280 ) | ( ~n6279 & n6281 ) | ( n6280 & n6281 ) ;
  assign n6283 = n6279 | n6282 ;
  assign n6284 = n6278 | n6283 ;
  assign n6285 = n6275 | n6284 ;
  assign n6286 = x953 & n5738 ;
  assign n6287 = x684 | n6286 ;
  assign n6288 = x1130 & n6286 ;
  assign n6289 = ( x962 & n6287 ) | ( x962 & ~n6288 ) | ( n6287 & ~n6288 ) ;
  assign n6290 = x1076 & n5965 ;
  assign n6291 = x382 & n5890 ;
  assign n6292 = x357 & n5892 ;
  assign n6293 = ( ~n6290 & n6291 ) | ( ~n6290 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6294 = n6290 | n6293 ;
  assign n6295 = n2621 & n5897 ;
  assign n6296 = x1067 & n6295 ;
  assign n6297 = ~x430 & n5895 ;
  assign n6298 = ( n5895 & n6296 ) | ( n5895 & ~n6297 ) | ( n6296 & ~n6297 ) ;
  assign n6299 = n6294 | n6298 ;
  assign n6300 = ~n2431 & n5897 ;
  assign n6301 = x1044 & n6300 ;
  assign n6302 = x657 & n5905 ;
  assign n6303 = ( n5905 & n6301 ) | ( n5905 & ~n6302 ) | ( n6301 & ~n6302 ) ;
  assign n6304 = x406 & n5879 ;
  assign n6305 = ~x728 & n5875 ;
  assign n6306 = ( ~n6303 & n6304 ) | ( ~n6303 & n6305 ) | ( n6304 & n6305 ) ;
  assign n6307 = n6303 | n6306 ;
  assign n6308 = x813 & n5886 ;
  assign n6309 = x860 & n5883 ;
  assign n6310 = ~x744 & n5871 ;
  assign n6311 = ( ~n6308 & n6309 ) | ( ~n6308 & n6310 ) | ( n6309 & n6310 ) ;
  assign n6312 = x652 & n5903 ;
  assign n6313 = n6308 | n6312 ;
  assign n6314 = n6311 | n6313 ;
  assign n6315 = ( ~n6299 & n6307 ) | ( ~n6299 & n6314 ) | ( n6307 & n6314 ) ;
  assign n6316 = n6299 | n6315 ;
  assign n6317 = x686 | n6286 ;
  assign n6318 = x1113 & n6286 ;
  assign n6319 = ( x962 & n6317 ) | ( x962 & ~n6318 ) | ( n6317 & ~n6318 ) ;
  assign n6320 = x687 & ~n6286 ;
  assign n6321 = x1127 & n6286 ;
  assign n6322 = ( ~x962 & n6320 ) | ( ~x962 & n6321 ) | ( n6320 & n6321 ) ;
  assign n6323 = x688 | n6286 ;
  assign n6324 = x1115 & n6286 ;
  assign n6325 = ( x962 & n6323 ) | ( x962 & ~n6324 ) | ( n6323 & ~n6324 ) ;
  assign n6326 = ~x752 & n5871 ;
  assign n6327 = x1036 & n6295 ;
  assign n6328 = x843 & n5883 ;
  assign n6329 = ( ~n6326 & n6327 ) | ( ~n6326 & n6328 ) | ( n6327 & n6328 ) ;
  assign n6330 = x401 & n5879 ;
  assign n6331 = n6326 | n6330 ;
  assign n6332 = n6329 | n6331 ;
  assign n6333 = x1079 & n5965 ;
  assign n6334 = x376 & n5890 ;
  assign n6335 = x351 & n5892 ;
  assign n6336 = ( ~n6333 & n6334 ) | ( ~n6333 & n6335 ) | ( n6334 & n6335 ) ;
  assign n6337 = n6333 | n6336 ;
  assign n6338 = x1049 & n6300 ;
  assign n6339 = x703 & n5875 ;
  assign n6340 = ( ~n6337 & n6338 ) | ( ~n6337 & n6339 ) | ( n6338 & n6339 ) ;
  assign n6341 = n6337 | n6340 ;
  assign n6342 = x798 & n5886 ;
  assign n6343 = ~x655 & n5905 ;
  assign n6344 = x426 & n5895 ;
  assign n6345 = ( ~n6342 & n6343 ) | ( ~n6342 & n6344 ) | ( n6343 & n6344 ) ;
  assign n6346 = x658 & n5903 ;
  assign n6347 = n6342 | n6346 ;
  assign n6348 = n6345 | n6347 ;
  assign n6349 = ( ~n6332 & n6341 ) | ( ~n6332 & n6348 ) | ( n6341 & n6348 ) ;
  assign n6350 = n6332 | n6349 ;
  assign n6351 = x690 & ~n6286 ;
  assign n6352 = x1108 & n6286 ;
  assign n6353 = ( ~x962 & n6351 ) | ( ~x962 & n6352 ) | ( n6351 & n6352 ) ;
  assign n6354 = x691 & ~n6286 ;
  assign n6355 = x1107 & n6286 ;
  assign n6356 = ( ~x962 & n6354 ) | ( ~x962 & n6355 ) | ( n6354 & n6355 ) ;
  assign n6357 = x844 & n5883 ;
  assign n6358 = x801 & n5886 ;
  assign n6359 = ~x770 & n5871 ;
  assign n6360 = ( ~n6357 & n6358 ) | ( ~n6357 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6361 = x656 & n5903 ;
  assign n6362 = n6357 | n6361 ;
  assign n6363 = n6360 | n6362 ;
  assign n6364 = ( ~x199 & n4068 ) | ( ~x199 & n4069 ) | ( n4068 & n4069 ) ;
  assign n6365 = x199 & x1078 ;
  assign n6366 = ( n5897 & n6364 ) | ( n5897 & n6365 ) | ( n6364 & n6365 ) ;
  assign n6367 = x352 & n5892 ;
  assign n6368 = x317 & n5890 ;
  assign n6369 = ( ~n6366 & n6367 ) | ( ~n6366 & n6368 ) | ( n6367 & n6368 ) ;
  assign n6370 = x427 | n6366 ;
  assign n6371 = ( n5895 & n6366 ) | ( n5895 & n6370 ) | ( n6366 & n6370 ) ;
  assign n6372 = n6369 | n6371 ;
  assign n6373 = ~x649 & n5905 ;
  assign n6374 = x402 & n5879 ;
  assign n6375 = x726 & n5875 ;
  assign n6376 = ( ~n6373 & n6374 ) | ( ~n6373 & n6375 ) | ( n6374 & n6375 ) ;
  assign n6377 = n6373 | n6376 ;
  assign n6378 = n6372 | n6377 ;
  assign n6379 = n6363 | n6378 ;
  assign n6380 = x693 | n5739 ;
  assign n6381 = x1129 & n5739 ;
  assign n6382 = ( x962 & n6380 ) | ( x962 & ~n6381 ) | ( n6380 & ~n6381 ) ;
  assign n6383 = x694 | n6286 ;
  assign n6384 = x1128 & n6286 ;
  assign n6385 = ( x962 & n6383 ) | ( x962 & ~n6384 ) | ( n6383 & ~n6384 ) ;
  assign n6386 = x695 | n5739 ;
  assign n6387 = x1111 & n5739 ;
  assign n6388 = ( x962 & n6386 ) | ( x962 & ~n6387 ) | ( n6386 & ~n6387 ) ;
  assign n6389 = x696 & ~n6286 ;
  assign n6390 = x1100 & n6286 ;
  assign n6391 = ( ~x962 & n6389 ) | ( ~x962 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6392 = x697 | n6286 ;
  assign n6393 = x1129 & n6286 ;
  assign n6394 = ( x962 & n6392 ) | ( x962 & ~n6393 ) | ( n6392 & ~n6393 ) ;
  assign n6395 = x698 | n6286 ;
  assign n6396 = x1116 & n6286 ;
  assign n6397 = ( x962 & n6395 ) | ( x962 & ~n6396 ) | ( n6395 & ~n6396 ) ;
  assign n6398 = x699 & ~n6286 ;
  assign n6399 = x1103 & n6286 ;
  assign n6400 = ( ~x962 & n6398 ) | ( ~x962 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6401 = x700 & ~n6286 ;
  assign n6402 = x1110 & n6286 ;
  assign n6403 = ( ~x962 & n6401 ) | ( ~x962 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6404 = x701 | n6286 ;
  assign n6405 = x1123 & n6286 ;
  assign n6406 = ( x962 & n6404 ) | ( x962 & ~n6405 ) | ( n6404 & ~n6405 ) ;
  assign n6407 = x702 | n6286 ;
  assign n6408 = x1117 & n6286 ;
  assign n6409 = ( x962 & n6407 ) | ( x962 & ~n6408 ) | ( n6407 & ~n6408 ) ;
  assign n6410 = x703 & ~n6286 ;
  assign n6411 = x1124 & n6286 ;
  assign n6412 = ( ~x962 & n6410 ) | ( ~x962 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6413 = x704 | n6286 ;
  assign n6414 = x1112 & n6286 ;
  assign n6415 = ( x962 & n6413 ) | ( x962 & ~n6414 ) | ( n6413 & ~n6414 ) ;
  assign n6416 = x705 & ~n6286 ;
  assign n6417 = x1125 & n6286 ;
  assign n6418 = ( ~x962 & n6416 ) | ( ~x962 & n6417 ) | ( n6416 & n6417 ) ;
  assign n6419 = x706 & ~n6286 ;
  assign n6420 = x1105 & n6286 ;
  assign n6421 = ( ~x962 & n6419 ) | ( ~x962 & n6420 ) | ( n6419 & n6420 ) ;
  assign n6422 = x1055 & n5965 ;
  assign n6423 = x347 & n5892 ;
  assign n6424 = x370 & n5890 ;
  assign n6425 = ( ~n6422 & n6423 ) | ( ~n6422 & n6424 ) | ( n6423 & n6424 ) ;
  assign n6426 = n6422 | n6425 ;
  assign n6427 = ~x753 & n5871 ;
  assign n6428 = x304 & n6300 ;
  assign n6429 = ( ~n6426 & n6427 ) | ( ~n6426 & n6428 ) | ( n6427 & n6428 ) ;
  assign n6430 = n6426 | n6429 ;
  assign n6431 = ~x702 & n5875 ;
  assign n6432 = x847 & n5883 ;
  assign n6433 = x627 & n5905 ;
  assign n6434 = ( ~n6431 & n6432 ) | ( ~n6431 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6435 = x395 & n5879 ;
  assign n6436 = n6431 | n6435 ;
  assign n6437 = n6434 | n6436 ;
  assign n6438 = x1048 & n6295 ;
  assign n6439 = x618 & n5903 ;
  assign n6440 = x420 & n5895 ;
  assign n6441 = ( ~n6438 & n6439 ) | ( ~n6438 & n6440 ) | ( n6439 & n6440 ) ;
  assign n6442 = n6438 | n6441 ;
  assign n6443 = n6437 | n6442 ;
  assign n6444 = n6430 | n6443 ;
  assign n6445 = x1058 & n5965 ;
  assign n6446 = x321 & n5892 ;
  assign n6447 = x442 & n5890 ;
  assign n6448 = ( ~n6445 & n6446 ) | ( ~n6445 & n6447 ) | ( n6446 & n6447 ) ;
  assign n6449 = n6445 | n6448 ;
  assign n6450 = x857 & n5883 ;
  assign n6451 = x305 & n6300 ;
  assign n6452 = ( ~n6449 & n6450 ) | ( ~n6449 & n6451 ) | ( n6450 & n6451 ) ;
  assign n6453 = n6449 | n6452 ;
  assign n6454 = ~x754 & n5871 ;
  assign n6455 = ~x709 & n5875 ;
  assign n6456 = x609 & n5903 ;
  assign n6457 = ( ~n6454 & n6455 ) | ( ~n6454 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = x328 & n5879 ;
  assign n6459 = n6454 | n6458 ;
  assign n6460 = n6457 | n6459 ;
  assign n6461 = x1084 & n6295 ;
  assign n6462 = x660 & n5905 ;
  assign n6463 = x459 & n5895 ;
  assign n6464 = ( ~n6461 & n6462 ) | ( ~n6461 & n6463 ) | ( n6462 & n6463 ) ;
  assign n6465 = n6461 | n6464 ;
  assign n6466 = n6460 | n6465 ;
  assign n6467 = n6453 | n6466 ;
  assign n6468 = x709 | n6286 ;
  assign n6469 = x1118 & n6286 ;
  assign n6470 = ( x962 & n6468 ) | ( x962 & ~n6469 ) | ( n6468 & ~n6469 ) ;
  assign n6471 = x710 & ~n5739 ;
  assign n6472 = x1106 & n5739 ;
  assign n6473 = ( ~x962 & n6471 ) | ( ~x962 & n6472 ) | ( n6471 & n6472 ) ;
  assign n6474 = x1087 & n5965 ;
  assign n6475 = x348 & n5892 ;
  assign n6476 = x373 & n5890 ;
  assign n6477 = ( ~n6474 & n6475 ) | ( ~n6474 & n6476 ) | ( n6475 & n6476 ) ;
  assign n6478 = n6474 | n6477 ;
  assign n6479 = x647 & n5905 ;
  assign n6480 = x306 & n6300 ;
  assign n6481 = ( ~n6478 & n6479 ) | ( ~n6478 & n6480 ) | ( n6479 & n6480 ) ;
  assign n6482 = n6478 | n6481 ;
  assign n6483 = x858 & n5883 ;
  assign n6484 = x630 & n5903 ;
  assign n6485 = x398 & n5879 ;
  assign n6486 = ( ~n6483 & n6484 ) | ( ~n6483 & n6485 ) | ( n6484 & n6485 ) ;
  assign n6487 = x423 & n5895 ;
  assign n6488 = n6483 | n6487 ;
  assign n6489 = n6486 | n6488 ;
  assign n6490 = ~x755 & n5871 ;
  assign n6491 = ~x725 & n5875 ;
  assign n6492 = x1059 & n6295 ;
  assign n6493 = ( ~n6490 & n6491 ) | ( ~n6490 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6494 = n6490 | n6493 ;
  assign n6495 = n6489 | n6494 ;
  assign n6496 = n6482 | n6495 ;
  assign n6497 = x374 & n5890 ;
  assign n6498 = x350 & n5892 ;
  assign n6499 = x1035 & n5965 ;
  assign n6500 = ( ~n6497 & n6498 ) | ( ~n6497 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6501 = n6497 | n6500 ;
  assign n6502 = x425 & n5895 ;
  assign n6503 = x842 & n5883 ;
  assign n6504 = ( ~n6501 & n6502 ) | ( ~n6501 & n6503 ) | ( n6502 & n6503 ) ;
  assign n6505 = n6501 | n6504 ;
  assign n6506 = x1044 & n6295 ;
  assign n6507 = x298 & n6300 ;
  assign n6508 = n6506 | n6507 ;
  assign n6509 = ~x751 & n5871 ;
  assign n6510 = x715 & n5905 ;
  assign n6511 = ( ~n6508 & n6509 ) | ( ~n6508 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6512 = n6508 | n6511 ;
  assign n6513 = ~x701 & n5875 ;
  assign n6514 = x400 & n5879 ;
  assign n6515 = x644 & n5903 ;
  assign n6516 = ( ~n6513 & n6514 ) | ( ~n6513 & n6515 ) | ( n6514 & n6515 ) ;
  assign n6517 = n6513 | n6516 ;
  assign n6518 = n6512 | n6517 ;
  assign n6519 = n6505 | n6518 ;
  assign n6520 = x1051 & n5965 ;
  assign n6521 = x371 & n5890 ;
  assign n6522 = x322 & n5892 ;
  assign n6523 = ( ~n6520 & n6521 ) | ( ~n6520 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6524 = n6520 | n6523 ;
  assign n6525 = x1072 & n6295 ;
  assign n6526 = x628 & n5905 ;
  assign n6527 = ( ~n6524 & n6525 ) | ( ~n6524 & n6526 ) | ( n6525 & n6526 ) ;
  assign n6528 = n6524 | n6527 ;
  assign n6529 = ~x734 & n5875 ;
  assign n6530 = x854 & n5883 ;
  assign n6531 = x396 & n5879 ;
  assign n6532 = ( ~n6529 & n6530 ) | ( ~n6529 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6533 = x309 & n6300 ;
  assign n6534 = n6529 | n6533 ;
  assign n6535 = n6532 | n6534 ;
  assign n6536 = ~x756 & n5871 ;
  assign n6537 = x629 & n5903 ;
  assign n6538 = x421 & n5895 ;
  assign n6539 = ( ~n6536 & n6537 ) | ( ~n6536 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6540 = n6536 | n6539 ;
  assign n6541 = n6535 | n6540 ;
  assign n6542 = n6528 | n6541 ;
  assign n6543 = x1057 & n5965 ;
  assign n6544 = x461 & n5892 ;
  assign n6545 = x439 & n5890 ;
  assign n6546 = ( ~n6543 & n6544 ) | ( ~n6543 & n6545 ) | ( n6544 & n6545 ) ;
  assign n6547 = n6543 | n6546 ;
  assign n6548 = ~x762 & n5871 ;
  assign n6549 = x1053 & n6300 ;
  assign n6550 = ( ~n6547 & n6548 ) | ( ~n6547 & n6549 ) | ( n6548 & n6549 ) ;
  assign n6551 = n6547 | n6550 ;
  assign n6552 = ~x693 & n5905 ;
  assign n6553 = x816 & n5886 ;
  assign n6554 = x326 & n5879 ;
  assign n6555 = ( ~n6552 & n6553 ) | ( ~n6552 & n6554 ) | ( n6553 & n6554 ) ;
  assign n6556 = x449 & n5895 ;
  assign n6557 = n6552 | n6556 ;
  assign n6558 = n6555 | n6557 ;
  assign n6559 = x1039 & n6295 ;
  assign n6560 = x867 & n5883 ;
  assign n6561 = x653 & n5903 ;
  assign n6562 = ( ~n6559 & n6560 ) | ( ~n6559 & n6561 ) | ( n6560 & n6561 ) ;
  assign n6563 = ~x697 & n5875 ;
  assign n6564 = n6559 | n6563 ;
  assign n6565 = n6562 | n6564 ;
  assign n6566 = n6558 | n6565 ;
  assign n6567 = n6551 | n6566 ;
  assign n6568 = x715 & ~n5739 ;
  assign n6569 = x1123 & n5739 ;
  assign n6570 = ( ~x962 & n6568 ) | ( ~x962 & n6569 ) | ( n6568 & n6569 ) ;
  assign n6571 = x626 & n5903 ;
  assign n6572 = x329 & n5879 ;
  assign n6573 = x641 & n5905 ;
  assign n6574 = ( ~n6571 & n6572 ) | ( ~n6571 & n6573 ) | ( n6572 & n6573 ) ;
  assign n6575 = n6571 | n6574 ;
  assign n6576 = x200 & x1053 ;
  assign n6577 = ~x200 & x307 ;
  assign n6578 = ( n5987 & n6576 ) | ( n5987 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6579 = x440 & n5890 ;
  assign n6580 = n6578 | n6579 ;
  assign n6581 = x349 & n5892 ;
  assign n6582 = x1043 & n5965 ;
  assign n6583 = ( ~n6580 & n6581 ) | ( ~n6580 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6584 = n6580 | n6583 ;
  assign n6585 = x454 & n5895 ;
  assign n6586 = ( ~n6575 & n6584 ) | ( ~n6575 & n6585 ) | ( n6584 & n6585 ) ;
  assign n6587 = n6575 | n6586 ;
  assign n6588 = ~x761 & n5871 ;
  assign n6589 = ~x738 & n5875 ;
  assign n6590 = x845 & n5883 ;
  assign n6591 = ( ~n6588 & n6589 ) | ( ~n6588 & n6590 ) | ( n6589 & n6590 ) ;
  assign n6592 = n6588 | n6591 ;
  assign n6593 = n6587 | n6592 ;
  assign n6594 = x1074 & n5965 ;
  assign n6595 = x462 & n5892 ;
  assign n6596 = x377 & n5890 ;
  assign n6597 = ( ~n6594 & n6595 ) | ( ~n6594 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6598 = n6594 | n6597 ;
  assign n6599 = x839 & n5883 ;
  assign n6600 = x1048 & n6300 ;
  assign n6601 = ( ~n6598 & n6599 ) | ( ~n6598 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6602 = n6598 | n6601 ;
  assign n6603 = x1070 & n6295 ;
  assign n6604 = x705 & n5875 ;
  assign n6605 = x645 & n5903 ;
  assign n6606 = ( ~n6603 & n6604 ) | ( ~n6603 & n6605 ) | ( n6604 & n6605 ) ;
  assign n6607 = x318 & n5879 ;
  assign n6608 = n6603 | n6607 ;
  assign n6609 = n6606 | n6608 ;
  assign n6610 = x800 & n5886 ;
  assign n6611 = ~x669 & n5905 ;
  assign n6612 = x448 & n5895 ;
  assign n6613 = ( ~n6610 & n6611 ) | ( ~n6610 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = ~x768 & n5871 ;
  assign n6615 = n6610 | n6614 ;
  assign n6616 = n6613 | n6615 ;
  assign n6617 = n6609 | n6616 ;
  assign n6618 = n6602 | n6617 ;
  assign n6619 = x1080 & n5965 ;
  assign n6620 = x369 & n5890 ;
  assign n6621 = n6619 | n6620 ;
  assign n6622 = x608 & n5903 ;
  assign n6623 = n6621 | n6622 ;
  assign n6624 = x315 & n5892 ;
  assign n6625 = x1049 & n6295 ;
  assign n6626 = ( ~n6623 & n6624 ) | ( ~n6623 & n6625 ) | ( n6624 & n6625 ) ;
  assign n6627 = n6623 | n6626 ;
  assign n6628 = ~x698 & n5875 ;
  assign n6629 = x853 & n5883 ;
  assign n6630 = x625 & n5905 ;
  assign n6631 = ( ~n6628 & n6629 ) | ( ~n6628 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6632 = x419 & n5895 ;
  assign n6633 = n6628 | n6632 ;
  assign n6634 = n6631 | n6633 ;
  assign n6635 = x394 & n5879 ;
  assign n6636 = x303 & n6300 ;
  assign n6637 = ~x767 & n5871 ;
  assign n6638 = ( ~n6635 & n6636 ) | ( ~n6635 & n6637 ) | ( n6636 & n6637 ) ;
  assign n6639 = n6635 | n6638 ;
  assign n6640 = n6634 | n6639 ;
  assign n6641 = n6627 | n6640 ;
  assign n6642 = x1063 & n5965 ;
  assign n6643 = x353 & n5892 ;
  assign n6644 = x378 & n5890 ;
  assign n6645 = ( ~n6642 & n6643 ) | ( ~n6642 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = n6642 | n6645 ;
  assign n6647 = ~x650 & n5905 ;
  assign n6648 = x1072 & n6300 ;
  assign n6649 = ( ~n6646 & n6647 ) | ( ~n6646 & n6648 ) | ( n6647 & n6648 ) ;
  assign n6650 = n6646 | n6649 ;
  assign n6651 = x636 & n5903 ;
  assign n6652 = x807 & n5886 ;
  assign n6653 = x325 & n5879 ;
  assign n6654 = ( ~n6651 & n6652 ) | ( ~n6651 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6655 = x451 & n5895 ;
  assign n6656 = n6651 | n6655 ;
  assign n6657 = n6654 | n6656 ;
  assign n6658 = x1062 & n6295 ;
  assign n6659 = ~x774 & n5871 ;
  assign n6660 = x687 & n5875 ;
  assign n6661 = ( ~n6658 & n6659 ) | ( ~n6658 & n6660 ) | ( n6659 & n6660 ) ;
  assign n6662 = x868 & n5883 ;
  assign n6663 = n6658 | n6662 ;
  assign n6664 = n6661 | n6663 ;
  assign n6665 = n6657 | n6664 ;
  assign n6666 = n6650 | n6665 ;
  assign n6667 = x1081 & n5965 ;
  assign n6668 = x381 & n5890 ;
  assign n6669 = x356 & n5892 ;
  assign n6670 = ( ~n6667 & n6668 ) | ( ~n6667 & n6669 ) | ( n6668 & n6669 ) ;
  assign n6671 = n6667 | n6670 ;
  assign n6672 = x794 & n5886 ;
  assign n6673 = x1040 & n6295 ;
  assign n6674 = ( ~n6671 & n6672 ) | ( ~n6671 & n6673 ) | ( n6672 & n6673 ) ;
  assign n6675 = n6671 | n6674 ;
  assign n6676 = x1037 & n6300 ;
  assign n6677 = ~x654 & n5905 ;
  assign n6678 = x445 & n5895 ;
  assign n6679 = ( ~n6676 & n6677 ) | ( ~n6676 & n6678 ) | ( n6677 & n6678 ) ;
  assign n6680 = x405 & n5879 ;
  assign n6681 = n6676 | n6680 ;
  assign n6682 = n6679 | n6681 ;
  assign n6683 = x880 & n5883 ;
  assign n6684 = ~x750 & n5871 ;
  assign n6685 = x651 & n5903 ;
  assign n6686 = ( ~n6683 & n6684 ) | ( ~n6683 & n6685 ) | ( n6684 & n6685 ) ;
  assign n6687 = ~x684 & n5875 ;
  assign n6688 = n6683 | n6687 ;
  assign n6689 = n6686 | n6688 ;
  assign n6690 = n6682 | n6689 ;
  assign n6691 = n6675 | n6690 ;
  assign n6692 = ~x769 & x794 ;
  assign n6693 = ( ~x747 & x807 ) | ( ~x747 & n6692 ) | ( x807 & n6692 ) ;
  assign n6694 = x769 & ~x794 ;
  assign n6695 = ( x747 & ~x807 ) | ( x747 & n6694 ) | ( ~x807 & n6694 ) ;
  assign n6696 = n6693 | n6695 ;
  assign n6697 = ~x771 & x800 ;
  assign n6698 = ( ~x721 & x813 ) | ( ~x721 & n6697 ) | ( x813 & n6697 ) ;
  assign n6699 = x771 & ~x800 ;
  assign n6700 = ( x721 & ~x813 ) | ( x721 & n6699 ) | ( ~x813 & n6699 ) ;
  assign n6701 = n6698 | n6700 ;
  assign n6702 = ~x765 & x798 ;
  assign n6703 = ( ~x731 & x795 ) | ( ~x731 & n6702 ) | ( x795 & n6702 ) ;
  assign n6704 = x765 & ~x798 ;
  assign n6705 = ( x731 & ~x795 ) | ( x731 & n6704 ) | ( ~x795 & n6704 ) ;
  assign n6706 = n6703 | n6705 ;
  assign n6707 = ( ~n6696 & n6701 ) | ( ~n6696 & n6706 ) | ( n6701 & n6706 ) ;
  assign n6708 = ~x775 & x816 ;
  assign n6709 = ( ~x773 & x801 ) | ( ~x773 & n6708 ) | ( x801 & n6708 ) ;
  assign n6710 = x775 & ~x816 ;
  assign n6711 = ( x773 & ~x801 ) | ( x773 & n6710 ) | ( ~x801 & n6710 ) ;
  assign n6712 = n6709 | n6711 ;
  assign n6713 = n6696 | n6712 ;
  assign n6714 = n6707 | n6713 ;
  assign n6715 = ~x945 & x988 ;
  assign n6716 = x773 & n6715 ;
  assign n6717 = x747 & n6716 ;
  assign n6718 = x731 & x775 ;
  assign n6719 = n6717 & n6718 ;
  assign n6720 = x769 & n6719 ;
  assign n6721 = x721 & ~n6720 ;
  assign n6722 = ~x721 & n6720 ;
  assign n6723 = ( n6714 & n6721 ) | ( n6714 & n6722 ) | ( n6721 & n6722 ) ;
  assign n6724 = x1059 & n6300 ;
  assign n6725 = x1069 & n6295 ;
  assign n6726 = n6724 | n6725 ;
  assign n6727 = ~x694 & n5875 ;
  assign n6728 = x795 & n5886 ;
  assign n6729 = ( ~n6726 & n6727 ) | ( ~n6726 & n6728 ) | ( n6727 & n6728 ) ;
  assign n6730 = n6726 | n6729 ;
  assign n6731 = x379 & n5890 ;
  assign n6732 = x354 & n5892 ;
  assign n6733 = x1045 & n5965 ;
  assign n6734 = ( ~n6731 & n6732 ) | ( ~n6731 & n6733 ) | ( n6732 & n6733 ) ;
  assign n6735 = n6731 | n6734 ;
  assign n6736 = ~x776 & n5871 ;
  assign n6737 = ~x732 & n5905 ;
  assign n6738 = ( ~n6735 & n6736 ) | ( ~n6735 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6739 = n6735 | n6738 ;
  assign n6740 = x851 & n5883 ;
  assign n6741 = x428 & n5895 ;
  assign n6742 = x403 & n5879 ;
  assign n6743 = ( ~n6740 & n6741 ) | ( ~n6740 & n6742 ) | ( n6741 & n6742 ) ;
  assign n6744 = x640 & n5903 ;
  assign n6745 = n6740 | n6744 ;
  assign n6746 = n6743 | n6745 ;
  assign n6747 = ( ~n6730 & n6739 ) | ( ~n6730 & n6746 ) | ( n6739 & n6746 ) ;
  assign n6748 = n6730 | n6747 ;
  assign n6749 = x723 | n6286 ;
  assign n6750 = x1111 & n6286 ;
  assign n6751 = ( x962 & n6749 ) | ( x962 & ~n6750 ) | ( n6749 & ~n6750 ) ;
  assign n6752 = x724 | n6286 ;
  assign n6753 = x1114 & n6286 ;
  assign n6754 = ( x962 & n6752 ) | ( x962 & ~n6753 ) | ( n6752 & ~n6753 ) ;
  assign n6755 = x725 | n6286 ;
  assign n6756 = x1120 & n6286 ;
  assign n6757 = ( x962 & n6755 ) | ( x962 & ~n6756 ) | ( n6755 & ~n6756 ) ;
  assign n6758 = x726 & ~n6286 ;
  assign n6759 = x1126 & n6286 ;
  assign n6760 = ( ~x962 & n6758 ) | ( ~x962 & n6759 ) | ( n6758 & n6759 ) ;
  assign n6761 = x727 & ~n6286 ;
  assign n6762 = x1102 & n6286 ;
  assign n6763 = ( ~x962 & n6761 ) | ( ~x962 & n6762 ) | ( n6761 & n6762 ) ;
  assign n6764 = x728 | n6286 ;
  assign n6765 = x1131 & n6286 ;
  assign n6766 = ( x962 & n6764 ) | ( x962 & ~n6765 ) | ( n6764 & ~n6765 ) ;
  assign n6767 = x729 & ~n6286 ;
  assign n6768 = x1104 & n6286 ;
  assign n6769 = ( ~x962 & n6767 ) | ( ~x962 & n6768 ) | ( n6767 & n6768 ) ;
  assign n6770 = x730 & ~n6286 ;
  assign n6771 = x1106 & n6286 ;
  assign n6772 = ( ~x962 & n6770 ) | ( ~x962 & n6771 ) | ( n6770 & n6771 ) ;
  assign n6773 = x731 & ~n6717 ;
  assign n6774 = ~x731 & n6717 ;
  assign n6775 = ( n6714 & n6773 ) | ( n6714 & n6774 ) | ( n6773 & n6774 ) ;
  assign n6776 = x732 | n5739 ;
  assign n6777 = x1128 & n5739 ;
  assign n6778 = ( x962 & n6776 ) | ( x962 & ~n6777 ) | ( n6776 & ~n6777 ) ;
  assign n6779 = x838 & n5883 ;
  assign n6780 = ~x737 & n5875 ;
  assign n6781 = x619 & n5903 ;
  assign n6782 = ( ~n6779 & n6780 ) | ( ~n6779 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6783 = ~x777 & n5871 ;
  assign n6784 = n6779 | n6783 ;
  assign n6785 = n6782 | n6784 ;
  assign n6786 = x375 & n5890 ;
  assign n6787 = x316 & n5892 ;
  assign n6788 = x1047 & n5965 ;
  assign n6789 = ( ~n6786 & n6787 ) | ( ~n6786 & n6788 ) | ( n6787 & n6788 ) ;
  assign n6790 = n6786 | n6789 ;
  assign n6791 = x424 & n5895 ;
  assign n6792 = x399 & n5879 ;
  assign n6793 = ( ~n6790 & n6791 ) | ( ~n6790 & n6792 ) | ( n6791 & n6792 ) ;
  assign n6794 = n6790 | n6793 ;
  assign n6795 = x648 & n5905 ;
  assign n6796 = x1037 & n6295 ;
  assign n6797 = x308 & n6300 ;
  assign n6798 = n6796 | n6797 ;
  assign n6799 = n6795 | n6798 ;
  assign n6800 = ( ~n6785 & n6794 ) | ( ~n6785 & n6799 ) | ( n6794 & n6799 ) ;
  assign n6801 = n6785 | n6800 ;
  assign n6802 = x734 | n6286 ;
  assign n6803 = x1119 & n6286 ;
  assign n6804 = ( x962 & n6802 ) | ( x962 & ~n6803 ) | ( n6802 & ~n6803 ) ;
  assign n6805 = x735 & ~n6286 ;
  assign n6806 = x1109 & n6286 ;
  assign n6807 = ( ~x962 & n6805 ) | ( ~x962 & n6806 ) | ( n6805 & n6806 ) ;
  assign n6808 = x736 & ~n6286 ;
  assign n6809 = x1101 & n6286 ;
  assign n6810 = ( ~x962 & n6808 ) | ( ~x962 & n6809 ) | ( n6808 & n6809 ) ;
  assign n6811 = x737 | n6286 ;
  assign n6812 = x1122 & n6286 ;
  assign n6813 = ( x962 & n6811 ) | ( x962 & ~n6812 ) | ( n6811 & ~n6812 ) ;
  assign n6814 = x738 | n6286 ;
  assign n6815 = x1121 & n6286 ;
  assign n6816 = ( x962 & n6814 ) | ( x962 & ~n6815 ) | ( n6814 & ~n6815 ) ;
  assign n6817 = ~x952 & n5649 ;
  assign n6818 = x739 | n6817 ;
  assign n6819 = ~x1108 & n6817 ;
  assign n6820 = ( x966 & n6818 ) | ( x966 & ~n6819 ) | ( n6818 & ~n6819 ) ;
  assign n6821 = x741 & ~n6817 ;
  assign n6822 = ~x1114 & n6817 ;
  assign n6823 = ( ~x966 & n6821 ) | ( ~x966 & n6822 ) | ( n6821 & n6822 ) ;
  assign n6824 = x742 & ~n6817 ;
  assign n6825 = ~x1112 & n6817 ;
  assign n6826 = ( ~x966 & n6824 ) | ( ~x966 & n6825 ) | ( n6824 & n6825 ) ;
  assign n6827 = x743 | n6817 ;
  assign n6828 = ~x1109 & n6817 ;
  assign n6829 = ( x966 & n6827 ) | ( x966 & ~n6828 ) | ( n6827 & ~n6828 ) ;
  assign n6830 = x744 & ~n6817 ;
  assign n6831 = ~x1131 & n6817 ;
  assign n6832 = ( ~x966 & n6830 ) | ( ~x966 & n6831 ) | ( n6830 & n6831 ) ;
  assign n6833 = x745 & ~n6817 ;
  assign n6834 = ~x1111 & n6817 ;
  assign n6835 = ( ~x966 & n6833 ) | ( ~x966 & n6834 ) | ( n6833 & n6834 ) ;
  assign n6836 = x746 | n6817 ;
  assign n6837 = ~x1104 & n6817 ;
  assign n6838 = ( x966 & n6836 ) | ( x966 & ~n6837 ) | ( n6836 & ~n6837 ) ;
  assign n6839 = ( x747 & n6714 ) | ( x747 & n6716 ) | ( n6714 & n6716 ) ;
  assign n6840 = ~n6717 & n6839 ;
  assign n6841 = x748 | n6817 ;
  assign n6842 = ~x1106 & n6817 ;
  assign n6843 = ( x966 & n6841 ) | ( x966 & ~n6842 ) | ( n6841 & ~n6842 ) ;
  assign n6844 = x749 | n6817 ;
  assign n6845 = ~x1105 & n6817 ;
  assign n6846 = ( x966 & n6844 ) | ( x966 & ~n6845 ) | ( n6844 & ~n6845 ) ;
  assign n6847 = x750 & ~n6817 ;
  assign n6848 = ~x1130 & n6817 ;
  assign n6849 = ( ~x966 & n6847 ) | ( ~x966 & n6848 ) | ( n6847 & n6848 ) ;
  assign n6850 = x751 & ~n6817 ;
  assign n6851 = ~x1123 & n6817 ;
  assign n6852 = ( ~x966 & n6850 ) | ( ~x966 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = x752 & ~n6817 ;
  assign n6854 = ~x1124 & n6817 ;
  assign n6855 = ( ~x966 & n6853 ) | ( ~x966 & n6854 ) | ( n6853 & n6854 ) ;
  assign n6856 = x753 & ~n6817 ;
  assign n6857 = ~x1117 & n6817 ;
  assign n6858 = ( ~x966 & n6856 ) | ( ~x966 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6859 = x754 & ~n6817 ;
  assign n6860 = ~x1118 & n6817 ;
  assign n6861 = ( ~x966 & n6859 ) | ( ~x966 & n6860 ) | ( n6859 & n6860 ) ;
  assign n6862 = x755 & ~n6817 ;
  assign n6863 = ~x1120 & n6817 ;
  assign n6864 = ( ~x966 & n6862 ) | ( ~x966 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6865 = x756 & ~n6817 ;
  assign n6866 = ~x1119 & n6817 ;
  assign n6867 = ( ~x966 & n6865 ) | ( ~x966 & n6866 ) | ( n6865 & n6866 ) ;
  assign n6868 = x757 & ~n6817 ;
  assign n6869 = ~x1113 & n6817 ;
  assign n6870 = ( ~x966 & n6868 ) | ( ~x966 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6871 = x758 | n6817 ;
  assign n6872 = ~x1101 & n6817 ;
  assign n6873 = ( x966 & n6871 ) | ( x966 & ~n6872 ) | ( n6871 & ~n6872 ) ;
  assign n6874 = x759 | n6817 ;
  assign n6875 = ~x1100 & n6817 ;
  assign n6876 = ( x966 & n6874 ) | ( x966 & ~n6875 ) | ( n6874 & ~n6875 ) ;
  assign n6877 = x760 & ~n6817 ;
  assign n6878 = ~x1115 & n6817 ;
  assign n6879 = ( ~x966 & n6877 ) | ( ~x966 & n6878 ) | ( n6877 & n6878 ) ;
  assign n6880 = x761 & ~n6817 ;
  assign n6881 = ~x1121 & n6817 ;
  assign n6882 = ( ~x966 & n6880 ) | ( ~x966 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6883 = x762 & ~n6817 ;
  assign n6884 = ~x1129 & n6817 ;
  assign n6885 = ( ~x966 & n6883 ) | ( ~x966 & n6884 ) | ( n6883 & n6884 ) ;
  assign n6886 = x763 | n6817 ;
  assign n6887 = ~x1103 & n6817 ;
  assign n6888 = ( x966 & n6886 ) | ( x966 & ~n6887 ) | ( n6886 & ~n6887 ) ;
  assign n6889 = x764 | n6817 ;
  assign n6890 = ~x1107 & n6817 ;
  assign n6891 = ( x966 & n6889 ) | ( x966 & ~n6890 ) | ( n6889 & ~n6890 ) ;
  assign n6892 = x794 | x800 ;
  assign n6893 = x721 | x731 ;
  assign n6894 = x765 | x773 ;
  assign n6895 = ( ~n6892 & n6893 ) | ( ~n6892 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6896 = x807 | x816 ;
  assign n6897 = n6892 | n6896 ;
  assign n6898 = n6895 | n6897 ;
  assign n6899 = ~n6714 & n6898 ;
  assign n6900 = x765 | x945 ;
  assign n6901 = x765 & x945 ;
  assign n6902 = ( n6899 & n6900 ) | ( n6899 & ~n6901 ) | ( n6900 & ~n6901 ) ;
  assign n6903 = x766 | n6817 ;
  assign n6904 = ~x1110 & n6817 ;
  assign n6905 = ( x966 & n6903 ) | ( x966 & ~n6904 ) | ( n6903 & ~n6904 ) ;
  assign n6906 = x767 & ~n6817 ;
  assign n6907 = ~x1116 & n6817 ;
  assign n6908 = ( ~x966 & n6906 ) | ( ~x966 & n6907 ) | ( n6906 & n6907 ) ;
  assign n6909 = x768 & ~n6817 ;
  assign n6910 = ~x1125 & n6817 ;
  assign n6911 = ( ~x966 & n6909 ) | ( ~x966 & n6910 ) | ( n6909 & n6910 ) ;
  assign n6912 = ( x769 & n6714 ) | ( x769 & n6719 ) | ( n6714 & n6719 ) ;
  assign n6913 = ~n6720 & n6912 ;
  assign n6914 = x770 & ~n6817 ;
  assign n6915 = ~x1126 & n6817 ;
  assign n6916 = ( ~x966 & n6914 ) | ( ~x966 & n6915 ) | ( n6914 & n6915 ) ;
  assign n6917 = x771 & x945 ;
  assign n6918 = ~x945 & x987 ;
  assign n6919 = ( ~n6899 & n6917 ) | ( ~n6899 & n6918 ) | ( n6917 & n6918 ) ;
  assign n6920 = x772 | n6817 ;
  assign n6921 = ~x1102 & n6817 ;
  assign n6922 = ( x966 & n6920 ) | ( x966 & ~n6921 ) | ( n6920 & ~n6921 ) ;
  assign n6923 = ( x773 & n6715 ) | ( x773 & ~n6899 ) | ( n6715 & ~n6899 ) ;
  assign n6924 = ~n6716 & n6923 ;
  assign n6925 = x774 & ~n6817 ;
  assign n6926 = ~x1127 & n6817 ;
  assign n6927 = ( ~x966 & n6925 ) | ( ~x966 & n6926 ) | ( n6925 & n6926 ) ;
  assign n6928 = x765 & ~x945 ;
  assign n6929 = x731 & x747 ;
  assign n6930 = x771 & x773 ;
  assign n6931 = ( ~n6928 & n6929 ) | ( ~n6928 & n6930 ) | ( n6929 & n6930 ) ;
  assign n6932 = n6928 & n6931 ;
  assign n6933 = x775 & ~n6932 ;
  assign n6934 = ~x775 & n6932 ;
  assign n6935 = ( n6714 & n6933 ) | ( n6714 & n6934 ) | ( n6933 & n6934 ) ;
  assign n6936 = x776 & ~n6817 ;
  assign n6937 = ~x1128 & n6817 ;
  assign n6938 = ( ~x966 & n6936 ) | ( ~x966 & n6937 ) | ( n6936 & n6937 ) ;
  assign n6939 = x777 & ~n6817 ;
  assign n6940 = ~x1122 & n6817 ;
  assign n6941 = ( ~x966 & n6939 ) | ( ~x966 & n6940 ) | ( n6939 & n6940 ) ;
  assign n6942 = x1046 | x1083 ;
  assign n6943 = ( ~x832 & x956 ) | ( ~x832 & x1085 ) | ( x956 & x1085 ) ;
  assign n6944 = ( x832 & n6942 ) | ( x832 & ~n6943 ) | ( n6942 & ~n6943 ) ;
  assign n6945 = x832 & ~n6944 ;
  assign n6946 = ~x968 & n6945 ;
  assign n6947 = ~x1100 & n6946 ;
  assign n6948 = x778 | n6946 ;
  assign n6949 = ~n6947 & n6948 ;
  assign n6950 = x779 & ~n5696 ;
  assign n6951 = x780 & ~n5627 ;
  assign n6952 = x781 & ~n6946 ;
  assign n6953 = x1101 & n6946 ;
  assign n6954 = n6952 | n6953 ;
  assign n6955 = n1683 & ~n5656 ;
  assign n6956 = n5626 & n6955 ;
  assign n6957 = x783 & ~n6946 ;
  assign n6958 = x1109 & n6946 ;
  assign n6959 = n6957 | n6958 ;
  assign n6960 = x784 & ~n6946 ;
  assign n6961 = x1110 & n6946 ;
  assign n6962 = n6960 | n6961 ;
  assign n6963 = x785 & ~n6946 ;
  assign n6964 = x1102 & n6946 ;
  assign n6965 = n6963 | n6964 ;
  assign n6966 = ~x786 & x954 ;
  assign n6967 = ( x24 & n1819 ) | ( x24 & ~n6966 ) | ( n1819 & ~n6966 ) ;
  assign n6968 = x787 & ~n6946 ;
  assign n6969 = x1104 & n6946 ;
  assign n6970 = n6968 | n6969 ;
  assign n6971 = x788 & ~n6946 ;
  assign n6972 = x1105 & n6946 ;
  assign n6973 = n6971 | n6972 ;
  assign n6974 = x789 & ~n6946 ;
  assign n6975 = x1106 & n6946 ;
  assign n6976 = n6974 | n6975 ;
  assign n6977 = x790 & ~n6946 ;
  assign n6978 = x1107 & n6946 ;
  assign n6979 = n6977 | n6978 ;
  assign n6980 = x791 & ~n6946 ;
  assign n6981 = x1108 & n6946 ;
  assign n6982 = n6980 | n6981 ;
  assign n6983 = x792 & ~n6946 ;
  assign n6984 = x1103 & n6946 ;
  assign n6985 = n6983 | n6984 ;
  assign n6986 = x968 & n6945 ;
  assign n6987 = ~x1130 & n6986 ;
  assign n6988 = x794 | n6986 ;
  assign n6989 = ~n6987 & n6988 ;
  assign n6990 = x795 & ~n6986 ;
  assign n6991 = x1128 & n6986 ;
  assign n6992 = n6990 | n6991 ;
  assign n6993 = ( x266 & x269 ) | ( x266 & x280 ) | ( x269 & x280 ) ;
  assign n6994 = x278 & x279 ;
  assign n6995 = ( x266 & n6993 ) | ( x266 & ~n6994 ) | ( n6993 & ~n6994 ) ;
  assign n6996 = x266 & ~n6995 ;
  assign n6997 = x264 | n6996 ;
  assign n6998 = ( x264 & n5847 ) | ( x264 & ~n6996 ) | ( n5847 & ~n6996 ) ;
  assign n6999 = ( ~n5848 & n6997 ) | ( ~n5848 & n6998 ) | ( n6997 & n6998 ) ;
  assign n7000 = x798 & ~n6986 ;
  assign n7001 = x1124 & n6986 ;
  assign n7002 = n7000 | n7001 ;
  assign n7003 = x799 | n6986 ;
  assign n7004 = x1107 & n6986 ;
  assign n7005 = n7003 & ~n7004 ;
  assign n7006 = x800 & ~n6986 ;
  assign n7007 = x1125 & n6986 ;
  assign n7008 = n7006 | n7007 ;
  assign n7009 = x801 & ~n6986 ;
  assign n7010 = x1126 & n6986 ;
  assign n7011 = n7009 | n7010 ;
  assign n7012 = x803 | n6986 ;
  assign n7013 = x1106 & n6986 ;
  assign n7014 = n7012 & ~n7013 ;
  assign n7015 = x804 & ~n6986 ;
  assign n7016 = x1109 & n6986 ;
  assign n7017 = n7015 | n7016 ;
  assign n7018 = n5844 & ~n5846 ;
  assign n7019 = ~x270 & n7018 ;
  assign n7020 = x270 & ~n7018 ;
  assign n7021 = n7019 | n7020 ;
  assign n7022 = x807 & ~n6986 ;
  assign n7023 = x1127 & n6986 ;
  assign n7024 = n7022 | n7023 ;
  assign n7025 = x808 & ~n6986 ;
  assign n7026 = x1101 & n6986 ;
  assign n7027 = n7025 | n7026 ;
  assign n7028 = x809 | n6986 ;
  assign n7029 = x1103 & n6986 ;
  assign n7030 = n7028 & ~n7029 ;
  assign n7031 = x810 & ~n6986 ;
  assign n7032 = x1108 & n6986 ;
  assign n7033 = n7031 | n7032 ;
  assign n7034 = x811 & ~n6986 ;
  assign n7035 = x1102 & n6986 ;
  assign n7036 = n7034 | n7035 ;
  assign n7037 = x812 | n6986 ;
  assign n7038 = x1104 & n6986 ;
  assign n7039 = n7037 & ~n7038 ;
  assign n7040 = x813 & ~n6986 ;
  assign n7041 = x1131 & n6986 ;
  assign n7042 = n7040 | n7041 ;
  assign n7043 = x814 | n6986 ;
  assign n7044 = x1105 & n6986 ;
  assign n7045 = n7043 & ~n7044 ;
  assign n7046 = x815 & ~n6986 ;
  assign n7047 = x1110 & n6986 ;
  assign n7048 = n7046 | n7047 ;
  assign n7049 = x816 & ~n6986 ;
  assign n7050 = x1129 & n6986 ;
  assign n7051 = n7049 | n7050 ;
  assign n7052 = x269 & ~n5843 ;
  assign n7053 = n5844 | n7052 ;
  assign n7054 = x265 & ~n5849 ;
  assign n7055 = n5850 | n7054 ;
  assign n7056 = x277 & n7019 ;
  assign n7057 = x277 | n7019 ;
  assign n7058 = ~n7056 & n7057 ;
  assign n7059 = x811 | x893 ;
  assign n7060 = n1463 & ~n2144 ;
  assign n7061 = ~x982 & x1092 ;
  assign n7062 = ( x1092 & n7060 ) | ( x1092 & n7061 ) | ( n7060 & n7061 ) ;
  assign n7063 = n1469 & n7062 ;
  assign n7064 = x123 & ~x222 ;
  assign n7065 = ~n1499 & n7064 ;
  assign n7066 = ( ~x1125 & x1126 ) | ( ~x1125 & x1130 ) | ( x1126 & x1130 ) ;
  assign n7067 = ( x1125 & x1126 ) | ( x1125 & x1130 ) | ( x1126 & x1130 ) ;
  assign n7068 = ( x1125 & n7066 ) | ( x1125 & ~n7067 ) | ( n7066 & ~n7067 ) ;
  assign n7069 = ( x1127 & ~x1131 ) | ( x1127 & n7068 ) | ( ~x1131 & n7068 ) ;
  assign n7070 = ( x1127 & x1131 ) | ( x1127 & ~n7068 ) | ( x1131 & ~n7068 ) ;
  assign n7071 = ( ~x1127 & n7069 ) | ( ~x1127 & n7070 ) | ( n7069 & n7070 ) ;
  assign n7072 = ( ~x1124 & x1128 ) | ( ~x1124 & x1129 ) | ( x1128 & x1129 ) ;
  assign n7073 = ( x1124 & x1128 ) | ( x1124 & x1129 ) | ( x1128 & x1129 ) ;
  assign n7074 = ( x1124 & n7072 ) | ( x1124 & ~n7073 ) | ( n7072 & ~n7073 ) ;
  assign n7075 = ( n7065 & ~n7071 ) | ( n7065 & n7074 ) | ( ~n7071 & n7074 ) ;
  assign n7076 = x825 & n7065 ;
  assign n7077 = n7071 & ~n7074 ;
  assign n7078 = ( n7075 & ~n7076 ) | ( n7075 & n7077 ) | ( ~n7076 & n7077 ) ;
  assign n7079 = ( ~x1117 & x1118 ) | ( ~x1117 & x1122 ) | ( x1118 & x1122 ) ;
  assign n7080 = ( x1117 & x1118 ) | ( x1117 & x1122 ) | ( x1118 & x1122 ) ;
  assign n7081 = ( x1117 & n7079 ) | ( x1117 & ~n7080 ) | ( n7079 & ~n7080 ) ;
  assign n7082 = ( x1119 & ~x1123 ) | ( x1119 & n7081 ) | ( ~x1123 & n7081 ) ;
  assign n7083 = ( x1119 & x1123 ) | ( x1119 & ~n7081 ) | ( x1123 & ~n7081 ) ;
  assign n7084 = ( ~x1119 & n7082 ) | ( ~x1119 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7085 = ( ~x1116 & x1120 ) | ( ~x1116 & x1121 ) | ( x1120 & x1121 ) ;
  assign n7086 = ( x1116 & x1120 ) | ( x1116 & x1121 ) | ( x1120 & x1121 ) ;
  assign n7087 = ( x1116 & n7085 ) | ( x1116 & ~n7086 ) | ( n7085 & ~n7086 ) ;
  assign n7088 = ( n7065 & ~n7084 ) | ( n7065 & n7087 ) | ( ~n7084 & n7087 ) ;
  assign n7089 = x826 & n7065 ;
  assign n7090 = n7084 & ~n7087 ;
  assign n7091 = ( n7088 & ~n7089 ) | ( n7088 & n7090 ) | ( ~n7089 & n7090 ) ;
  assign n7092 = ( ~x1101 & x1103 ) | ( ~x1101 & x1106 ) | ( x1103 & x1106 ) ;
  assign n7093 = ( x1101 & x1103 ) | ( x1101 & x1106 ) | ( x1103 & x1106 ) ;
  assign n7094 = ( x1101 & n7092 ) | ( x1101 & ~n7093 ) | ( n7092 & ~n7093 ) ;
  assign n7095 = ( x1102 & ~x1107 ) | ( x1102 & n7094 ) | ( ~x1107 & n7094 ) ;
  assign n7096 = ( x1102 & x1107 ) | ( x1102 & ~n7094 ) | ( x1107 & ~n7094 ) ;
  assign n7097 = ( ~x1102 & n7095 ) | ( ~x1102 & n7096 ) | ( n7095 & n7096 ) ;
  assign n7098 = ( ~x1100 & x1104 ) | ( ~x1100 & x1105 ) | ( x1104 & x1105 ) ;
  assign n7099 = ( x1100 & x1104 ) | ( x1100 & x1105 ) | ( x1104 & x1105 ) ;
  assign n7100 = ( x1100 & n7098 ) | ( x1100 & ~n7099 ) | ( n7098 & ~n7099 ) ;
  assign n7101 = ( n7065 & ~n7097 ) | ( n7065 & n7100 ) | ( ~n7097 & n7100 ) ;
  assign n7102 = x827 & n7065 ;
  assign n7103 = n7097 & ~n7100 ;
  assign n7104 = ( n7101 & ~n7102 ) | ( n7101 & n7103 ) | ( ~n7102 & n7103 ) ;
  assign n7105 = ( ~x1109 & x1111 ) | ( ~x1109 & x1114 ) | ( x1111 & x1114 ) ;
  assign n7106 = ( x1109 & x1111 ) | ( x1109 & x1114 ) | ( x1111 & x1114 ) ;
  assign n7107 = ( x1109 & n7105 ) | ( x1109 & ~n7106 ) | ( n7105 & ~n7106 ) ;
  assign n7108 = ( x1108 & ~x1115 ) | ( x1108 & n7107 ) | ( ~x1115 & n7107 ) ;
  assign n7109 = ( x1108 & x1115 ) | ( x1108 & ~n7107 ) | ( x1115 & ~n7107 ) ;
  assign n7110 = ( ~x1108 & n7108 ) | ( ~x1108 & n7109 ) | ( n7108 & n7109 ) ;
  assign n7111 = ( ~x1110 & x1112 ) | ( ~x1110 & x1113 ) | ( x1112 & x1113 ) ;
  assign n7112 = ( x1110 & x1112 ) | ( x1110 & x1113 ) | ( x1112 & x1113 ) ;
  assign n7113 = ( x1110 & n7111 ) | ( x1110 & ~n7112 ) | ( n7111 & ~n7112 ) ;
  assign n7114 = ( n7065 & ~n7110 ) | ( n7065 & n7113 ) | ( ~n7110 & n7113 ) ;
  assign n7115 = x828 & n7065 ;
  assign n7116 = n7110 & ~n7113 ;
  assign n7117 = ( n7114 & ~n7115 ) | ( n7114 & n7116 ) | ( ~n7115 & n7116 ) ;
  assign n7118 = ~n2144 & n3692 ;
  assign n7119 = ~x951 & x1092 ;
  assign n7120 = ( x1092 & n7118 ) | ( x1092 & n7119 ) | ( n7118 & n7119 ) ;
  assign n7121 = x281 & n6996 ;
  assign n7122 = x281 | n6996 ;
  assign n7123 = ~n7121 & n7122 ;
  assign n7124 = ~x832 & x1091 ;
  assign n7125 = n1843 & n7124 ;
  assign n7126 = x833 | n1841 ;
  assign n7127 = ~n1871 & n7126 ;
  assign n7128 = x946 & n1841 ;
  assign n7129 = x281 & x282 ;
  assign n7130 = ( ~x281 & x282 ) | ( ~x281 & n5844 ) | ( x282 & n5844 ) ;
  assign n7131 = x282 & n5844 ;
  assign n7132 = ( n7129 & n7130 ) | ( n7129 & ~n7131 ) | ( n7130 & ~n7131 ) ;
  assign n7133 = x837 & x955 ;
  assign n7134 = ~x955 & x1049 ;
  assign n7135 = n7133 | n7134 ;
  assign n7136 = x838 & x955 ;
  assign n7137 = ~x955 & x1047 ;
  assign n7138 = n7136 | n7137 ;
  assign n7139 = x839 & x955 ;
  assign n7140 = ~x955 & x1074 ;
  assign n7141 = n7139 | n7140 ;
  assign n7142 = x840 & ~n1841 ;
  assign n7143 = x1196 & n1841 ;
  assign n7144 = n7142 | n7143 ;
  assign n7145 = x842 & x955 ;
  assign n7146 = ~x955 & x1035 ;
  assign n7147 = n7145 | n7146 ;
  assign n7148 = x843 & x955 ;
  assign n7149 = ~x955 & x1079 ;
  assign n7150 = n7148 | n7149 ;
  assign n7151 = x844 & x955 ;
  assign n7152 = ~x955 & x1078 ;
  assign n7153 = n7151 | n7152 ;
  assign n7154 = x845 & x955 ;
  assign n7155 = ~x955 & x1043 ;
  assign n7156 = n7154 | n7155 ;
  assign n7157 = x846 & ~n4097 ;
  assign n7158 = ( x1134 & n4095 ) | ( x1134 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7159 = n7157 | n7158 ;
  assign n7160 = x847 & x955 ;
  assign n7161 = ~x955 & x1055 ;
  assign n7162 = n7160 | n7161 ;
  assign n7163 = x848 & x955 ;
  assign n7164 = ~x955 & x1039 ;
  assign n7165 = n7163 | n7164 ;
  assign n7166 = x849 & ~n1841 ;
  assign n7167 = x1198 & n1841 ;
  assign n7168 = n7166 | n7167 ;
  assign n7169 = x850 & x955 ;
  assign n7170 = ~x955 & x1048 ;
  assign n7171 = n7169 | n7170 ;
  assign n7172 = x851 & x955 ;
  assign n7173 = ~x955 & x1045 ;
  assign n7174 = n7172 | n7173 ;
  assign n7175 = x852 & x955 ;
  assign n7176 = ~x955 & x1062 ;
  assign n7177 = n7175 | n7176 ;
  assign n7178 = x853 & x955 ;
  assign n7179 = ~x955 & x1080 ;
  assign n7180 = n7178 | n7179 ;
  assign n7181 = x854 & x955 ;
  assign n7182 = ~x955 & x1051 ;
  assign n7183 = n7181 | n7182 ;
  assign n7184 = x855 & x955 ;
  assign n7185 = ~x955 & x1065 ;
  assign n7186 = n7184 | n7185 ;
  assign n7187 = x856 & x955 ;
  assign n7188 = ~x955 & x1067 ;
  assign n7189 = n7187 | n7188 ;
  assign n7190 = x857 & x955 ;
  assign n7191 = ~x955 & x1058 ;
  assign n7192 = n7190 | n7191 ;
  assign n7193 = x858 & x955 ;
  assign n7194 = ~x955 & x1087 ;
  assign n7195 = n7193 | n7194 ;
  assign n7196 = x859 & x955 ;
  assign n7197 = ~x955 & x1070 ;
  assign n7198 = n7196 | n7197 ;
  assign n7199 = x860 & x955 ;
  assign n7200 = ~x955 & x1076 ;
  assign n7201 = n7199 | n7200 ;
  assign n7202 = x861 & ~n4097 ;
  assign n7203 = ( x1141 & n4095 ) | ( x1141 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7204 = n7202 | n7203 ;
  assign n7205 = x862 & ~n4097 ;
  assign n7206 = ( x1139 & n4095 ) | ( x1139 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7207 = n7205 | n7206 ;
  assign n7208 = x863 & ~n1841 ;
  assign n7209 = x1199 & n1841 ;
  assign n7210 = n7208 | n7209 ;
  assign n7211 = x864 & ~n1841 ;
  assign n7212 = x1197 & n1841 ;
  assign n7213 = n7211 | n7212 ;
  assign n7214 = x865 & x955 ;
  assign n7215 = ~x955 & x1040 ;
  assign n7216 = n7214 | n7215 ;
  assign n7217 = x866 & x955 ;
  assign n7218 = ~x955 & x1053 ;
  assign n7219 = n7217 | n7218 ;
  assign n7220 = x867 & x955 ;
  assign n7221 = ~x955 & x1057 ;
  assign n7222 = n7220 | n7221 ;
  assign n7223 = x868 & x955 ;
  assign n7224 = ~x955 & x1063 ;
  assign n7225 = n7223 | n7224 ;
  assign n7226 = x869 & ~n4097 ;
  assign n7227 = ( x1140 & n4095 ) | ( x1140 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7228 = n7226 | n7227 ;
  assign n7229 = x870 & x955 ;
  assign n7230 = ~x955 & x1069 ;
  assign n7231 = n7229 | n7230 ;
  assign n7232 = x871 & x955 ;
  assign n7233 = ~x955 & x1072 ;
  assign n7234 = n7232 | n7233 ;
  assign n7235 = x872 & x955 ;
  assign n7236 = ~x955 & x1084 ;
  assign n7237 = n7235 | n7236 ;
  assign n7238 = x873 & x955 ;
  assign n7239 = ~x955 & x1044 ;
  assign n7240 = n7238 | n7239 ;
  assign n7241 = x874 & x955 ;
  assign n7242 = ~x955 & x1036 ;
  assign n7243 = n7241 | n7242 ;
  assign n7244 = x875 & ~n4097 ;
  assign n7245 = ( x1136 & n4095 ) | ( x1136 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7246 = n7244 | n7245 ;
  assign n7247 = x876 & x955 ;
  assign n7248 = ~x955 & x1037 ;
  assign n7249 = n7247 | n7248 ;
  assign n7250 = x877 & ~n4097 ;
  assign n7251 = ( x1138 & n4095 ) | ( x1138 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7252 = n7250 | n7251 ;
  assign n7253 = x878 & ~n4097 ;
  assign n7254 = ( x1137 & n4095 ) | ( x1137 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7255 = n7253 | n7254 ;
  assign n7256 = x879 & ~n4097 ;
  assign n7257 = ( x1135 & n4095 ) | ( x1135 & n4096 ) | ( n4095 & n4096 ) ;
  assign n7258 = n7256 | n7257 ;
  assign n7259 = x880 & x955 ;
  assign n7260 = ~x955 & x1081 ;
  assign n7261 = n7259 | n7260 ;
  assign n7262 = x881 & x955 ;
  assign n7263 = ~x955 & x1059 ;
  assign n7264 = n7262 | n7263 ;
  assign n7265 = ~x883 & n7065 ;
  assign n7266 = x1107 & ~n7065 ;
  assign n7267 = n7265 | n7266 ;
  assign n7268 = ~x884 & n7065 ;
  assign n7269 = x1124 & ~n7065 ;
  assign n7270 = n7268 | n7269 ;
  assign n7271 = ~x885 & n7065 ;
  assign n7272 = x1125 & ~n7065 ;
  assign n7273 = n7271 | n7272 ;
  assign n7274 = ~x886 & n7065 ;
  assign n7275 = x1109 & ~n7065 ;
  assign n7276 = n7274 | n7275 ;
  assign n7277 = ~x887 & n7065 ;
  assign n7278 = x1100 & ~n7065 ;
  assign n7279 = n7277 | n7278 ;
  assign n7280 = ~x888 & n7065 ;
  assign n7281 = x1120 & ~n7065 ;
  assign n7282 = n7280 | n7281 ;
  assign n7283 = ~x889 & n7065 ;
  assign n7284 = x1103 & ~n7065 ;
  assign n7285 = n7283 | n7284 ;
  assign n7286 = ~x890 & n7065 ;
  assign n7287 = x1126 & ~n7065 ;
  assign n7288 = n7286 | n7287 ;
  assign n7289 = ~x891 & n7065 ;
  assign n7290 = x1116 & ~n7065 ;
  assign n7291 = n7289 | n7290 ;
  assign n7292 = ~x892 & n7065 ;
  assign n7293 = x1101 & ~n7065 ;
  assign n7294 = n7292 | n7293 ;
  assign n7295 = ~x894 & n7065 ;
  assign n7296 = x1119 & ~n7065 ;
  assign n7297 = n7295 | n7296 ;
  assign n7298 = ~x895 & n7065 ;
  assign n7299 = x1113 & ~n7065 ;
  assign n7300 = n7298 | n7299 ;
  assign n7301 = ~x896 & n7065 ;
  assign n7302 = x1118 & ~n7065 ;
  assign n7303 = n7301 | n7302 ;
  assign n7304 = ~x898 & n7065 ;
  assign n7305 = x1129 & ~n7065 ;
  assign n7306 = n7304 | n7305 ;
  assign n7307 = ~x899 & n7065 ;
  assign n7308 = x1115 & ~n7065 ;
  assign n7309 = n7307 | n7308 ;
  assign n7310 = ~x900 & n7065 ;
  assign n7311 = x1110 & ~n7065 ;
  assign n7312 = n7310 | n7311 ;
  assign n7313 = ~x902 & n7065 ;
  assign n7314 = x1111 & ~n7065 ;
  assign n7315 = n7313 | n7314 ;
  assign n7316 = ~x903 & n7065 ;
  assign n7317 = x1121 & ~n7065 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = ~x904 & n7065 ;
  assign n7320 = x1127 & ~n7065 ;
  assign n7321 = n7319 | n7320 ;
  assign n7322 = ~x905 & n7065 ;
  assign n7323 = x1131 & ~n7065 ;
  assign n7324 = n7322 | n7323 ;
  assign n7325 = ~x906 & n7065 ;
  assign n7326 = x1128 & ~n7065 ;
  assign n7327 = n7325 | n7326 ;
  assign n7328 = ~x598 & x979 ;
  assign n7329 = x615 & n7328 ;
  assign n7330 = ~x782 & x907 ;
  assign n7331 = x624 | x979 ;
  assign n7332 = ~n7328 & n7331 ;
  assign n7333 = ( x604 & n7328 ) | ( x604 & ~n7332 ) | ( n7328 & ~n7332 ) ;
  assign n7334 = ( x782 & n7330 ) | ( x782 & n7333 ) | ( n7330 & n7333 ) ;
  assign n7335 = ( ~n7329 & n7330 ) | ( ~n7329 & n7334 ) | ( n7330 & n7334 ) ;
  assign n7336 = ~x908 & n7065 ;
  assign n7337 = x1122 & ~n7065 ;
  assign n7338 = n7336 | n7337 ;
  assign n7339 = ~x909 & n7065 ;
  assign n7340 = x1105 & ~n7065 ;
  assign n7341 = n7339 | n7340 ;
  assign n7342 = ~x910 & n7065 ;
  assign n7343 = x1117 & ~n7065 ;
  assign n7344 = n7342 | n7343 ;
  assign n7345 = ~x911 & n7065 ;
  assign n7346 = x1130 & ~n7065 ;
  assign n7347 = n7345 | n7346 ;
  assign n7348 = ~x912 & n7065 ;
  assign n7349 = x1114 & ~n7065 ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = ~x913 & n7065 ;
  assign n7352 = x1106 & ~n7065 ;
  assign n7353 = n7351 | n7352 ;
  assign n7354 = x280 & ~n5842 ;
  assign n7355 = n5843 | n7354 ;
  assign n7356 = ~x915 & n7065 ;
  assign n7357 = x1108 & ~n7065 ;
  assign n7358 = n7356 | n7357 ;
  assign n7359 = ~x916 & n7065 ;
  assign n7360 = x1123 & ~n7065 ;
  assign n7361 = n7359 | n7360 ;
  assign n7362 = ~x917 & n7065 ;
  assign n7363 = x1112 & ~n7065 ;
  assign n7364 = n7362 | n7363 ;
  assign n7365 = ~x918 & n7065 ;
  assign n7366 = x1104 & ~n7065 ;
  assign n7367 = n7365 | n7366 ;
  assign n7368 = ~x919 & n7065 ;
  assign n7369 = x1102 & ~n7065 ;
  assign n7370 = n7368 | n7369 ;
  assign n7371 = x920 & ~x1093 ;
  assign n7372 = x1093 & x1139 ;
  assign n7373 = n7371 | n7372 ;
  assign n7374 = x921 & ~x1093 ;
  assign n7375 = x1093 & x1140 ;
  assign n7376 = n7374 | n7375 ;
  assign n7377 = x922 & ~x1093 ;
  assign n7378 = x1093 & x1152 ;
  assign n7379 = n7377 | n7378 ;
  assign n7380 = x923 & ~x1093 ;
  assign n7381 = x1093 & x1154 ;
  assign n7382 = n7380 | n7381 ;
  assign n7383 = ~x300 & x301 ;
  assign n7384 = x311 & ~x312 ;
  assign n7385 = n7383 & n7384 ;
  assign n7386 = x925 & ~x1093 ;
  assign n7387 = x1093 & x1155 ;
  assign n7388 = n7386 | n7387 ;
  assign n7389 = x926 & ~x1093 ;
  assign n7390 = x1093 & x1157 ;
  assign n7391 = n7389 | n7390 ;
  assign n7392 = x927 & ~x1093 ;
  assign n7393 = x1093 & x1145 ;
  assign n7394 = n7392 | n7393 ;
  assign n7395 = x928 & ~x1093 ;
  assign n7396 = x1093 & x1136 ;
  assign n7397 = n7395 | n7396 ;
  assign n7398 = x929 & ~x1093 ;
  assign n7399 = x1093 & x1144 ;
  assign n7400 = n7398 | n7399 ;
  assign n7401 = x930 & ~x1093 ;
  assign n7402 = x1093 & x1134 ;
  assign n7403 = n7401 | n7402 ;
  assign n7404 = x931 & ~x1093 ;
  assign n7405 = x1093 & x1150 ;
  assign n7406 = n7404 | n7405 ;
  assign n7407 = x932 & ~x1093 ;
  assign n7408 = x1093 & x1142 ;
  assign n7409 = n7407 | n7408 ;
  assign n7410 = x933 & ~x1093 ;
  assign n7411 = x1093 & x1137 ;
  assign n7412 = n7410 | n7411 ;
  assign n7413 = x934 & ~x1093 ;
  assign n7414 = x1093 & x1147 ;
  assign n7415 = n7413 | n7414 ;
  assign n7416 = x935 & ~x1093 ;
  assign n7417 = x1093 & x1141 ;
  assign n7418 = n7416 | n7417 ;
  assign n7419 = x936 & ~x1093 ;
  assign n7420 = x1093 & x1149 ;
  assign n7421 = n7419 | n7420 ;
  assign n7422 = x937 & ~x1093 ;
  assign n7423 = x1093 & x1148 ;
  assign n7424 = n7422 | n7423 ;
  assign n7425 = x938 & ~x1093 ;
  assign n7426 = x1093 & x1135 ;
  assign n7427 = n7425 | n7426 ;
  assign n7428 = x939 & ~x1093 ;
  assign n7429 = x1093 & x1146 ;
  assign n7430 = n7428 | n7429 ;
  assign n7431 = x940 & ~x1093 ;
  assign n7432 = x1093 & x1138 ;
  assign n7433 = n7431 | n7432 ;
  assign n7434 = x941 & ~x1093 ;
  assign n7435 = x1093 & x1153 ;
  assign n7436 = n7434 | n7435 ;
  assign n7437 = x942 & ~x1093 ;
  assign n7438 = x1093 & x1156 ;
  assign n7439 = n7437 | n7438 ;
  assign n7440 = x943 & ~x1093 ;
  assign n7441 = x1093 & x1151 ;
  assign n7442 = n7440 | n7441 ;
  assign n7443 = x944 & ~x1093 ;
  assign n7444 = x1093 & x1143 ;
  assign n7445 = n7443 | n7444 ;
  assign n7446 = ~x782 & x947 ;
  assign n7447 = x782 | x947 ;
  assign n7448 = ( n7332 & n7446 ) | ( n7332 & n7447 ) | ( n7446 & n7447 ) ;
  assign n7449 = x266 | x992 ;
  assign n7450 = ~n5842 & n7449 ;
  assign n7451 = x949 & x954 ;
  assign n7452 = ( x313 & n4400 ) | ( x313 & ~n7451 ) | ( n4400 & ~n7451 ) ;
  assign n7453 = n1467 & n1841 ;
  assign n7454 = x957 & x1092 ;
  assign n7455 = x31 | n7454 ;
  assign n7456 = ~x782 & x960 ;
  assign n7457 = ~x230 & x961 ;
  assign n7458 = ~x782 & x963 ;
  assign n7459 = ~x230 & x967 ;
  assign n7460 = ~x230 & x969 ;
  assign n7461 = ~x782 & x970 ;
  assign n7462 = ~x230 & x971 ;
  assign n7463 = ~x782 & x972 ;
  assign n7464 = ~x230 & x974 ;
  assign n7465 = ~x782 & x975 ;
  assign n7466 = ~x230 & x977 ;
  assign n7467 = ~x782 & x978 ;
  assign n7468 = ~x598 & x615 ;
  assign n7469 = x604 | x624 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = n1516 ;
  assign y154 = n1531 ;
  assign y155 = n1540 ;
  assign y156 = ~n1551 ;
  assign y157 = ~n1562 ;
  assign y158 = n1573 ;
  assign y159 = n1584 ;
  assign y160 = n1595 ;
  assign y161 = n1606 ;
  assign y162 = n1617 ;
  assign y163 = n1628 ;
  assign y164 = n1639 ;
  assign y165 = n1650 ;
  assign y166 = ~1'b0 ;
  assign y167 = n1750 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n1792 ;
  assign y172 = ~n1798 ;
  assign y173 = ~n1802 ;
  assign y174 = ~n1805 ;
  assign y175 = ~n1808 ;
  assign y176 = ~n1811 ;
  assign y177 = ~n1814 ;
  assign y178 = ~n1817 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = n1750 ;
  assign y182 = n1821 ;
  assign y183 = n1828 ;
  assign y184 = ~n1833 ;
  assign y185 = ~n1835 ;
  assign y186 = ~n1837 ;
  assign y187 = ~n1839 ;
  assign y188 = x37 ;
  assign y189 = n2147 ;
  assign y190 = n2185 ;
  assign y191 = n2270 ;
  assign y192 = n2325 ;
  assign y193 = n2349 ;
  assign y194 = n2356 ;
  assign y195 = n1818 ;
  assign y196 = n2362 ;
  assign y197 = n2381 ;
  assign y198 = n2384 ;
  assign y199 = n2421 ;
  assign y200 = n2447 ;
  assign y201 = n2467 ;
  assign y202 = n2474 ;
  assign y203 = n2477 ;
  assign y204 = n2482 ;
  assign y205 = n2496 ;
  assign y206 = n2498 ;
  assign y207 = n2502 ;
  assign y208 = n2514 ;
  assign y209 = n2515 ;
  assign y210 = n2530 ;
  assign y211 = n2539 ;
  assign y212 = n2543 ;
  assign y213 = n2546 ;
  assign y214 = n2551 ;
  assign y215 = n2559 ;
  assign y216 = n2561 ;
  assign y217 = n2567 ;
  assign y218 = n2573 ;
  assign y219 = n2576 ;
  assign y220 = n2579 ;
  assign y221 = n2584 ;
  assign y222 = n2586 ;
  assign y223 = n2588 ;
  assign y224 = n2594 ;
  assign y225 = n2596 ;
  assign y226 = n2600 ;
  assign y227 = n2603 ;
  assign y228 = n2618 ;
  assign y229 = n2626 ;
  assign y230 = n2634 ;
  assign y231 = n2642 ;
  assign y232 = n2651 ;
  assign y233 = n2655 ;
  assign y234 = n2660 ;
  assign y235 = n2664 ;
  assign y236 = n2665 ;
  assign y237 = n2713 ;
  assign y238 = n2721 ;
  assign y239 = n2724 ;
  assign y240 = n2726 ;
  assign y241 = n2729 ;
  assign y242 = n2731 ;
  assign y243 = n2734 ;
  assign y244 = n2736 ;
  assign y245 = n2737 ;
  assign y246 = n2742 ;
  assign y247 = n2745 ;
  assign y248 = n2748 ;
  assign y249 = n2754 ;
  assign y250 = n2756 ;
  assign y251 = n2759 ;
  assign y252 = n2764 ;
  assign y253 = n2771 ;
  assign y254 = n2776 ;
  assign y255 = n2783 ;
  assign y256 = n2786 ;
  assign y257 = n2793 ;
  assign y258 = n2797 ;
  assign y259 = n2803 ;
  assign y260 = n2805 ;
  assign y261 = n2807 ;
  assign y262 = n2813 ;
  assign y263 = x117 ;
  assign y264 = n2816 ;
  assign y265 = n2817 ;
  assign y266 = n2822 ;
  assign y267 = n2663 ;
  assign y268 = n2829 ;
  assign y269 = n2833 ;
  assign y270 = ~n2834 ;
  assign y271 = n2838 ;
  assign y272 = n2841 ;
  assign y273 = n2845 ;
  assign y274 = n2848 ;
  assign y275 = n1827 ;
  assign y276 = n2894 ;
  assign y277 = n2908 ;
  assign y278 = n2917 ;
  assign y279 = n2968 ;
  assign y280 = n1878 ;
  assign y281 = ~n2984 ;
  assign y282 = n3007 ;
  assign y283 = n3030 ;
  assign y284 = n3040 ;
  assign y285 = x131 ;
  assign y286 = n3046 ;
  assign y287 = n3057 ;
  assign y288 = n2905 ;
  assign y289 = n3083 ;
  assign y290 = n3095 ;
  assign y291 = n3105 ;
  assign y292 = n3115 ;
  assign y293 = n3123 ;
  assign y294 = n3130 ;
  assign y295 = n3136 ;
  assign y296 = n3141 ;
  assign y297 = ~n3224 ;
  assign y298 = ~n3230 ;
  assign y299 = n3235 ;
  assign y300 = ~n3240 ;
  assign y301 = n3245 ;
  assign y302 = ~n3250 ;
  assign y303 = n3258 ;
  assign y304 = ~n3263 ;
  assign y305 = ~n3268 ;
  assign y306 = ~n3273 ;
  assign y307 = ~n3278 ;
  assign y308 = ~n3283 ;
  assign y309 = n3288 ;
  assign y310 = ~n3293 ;
  assign y311 = ~n3298 ;
  assign y312 = ~n3303 ;
  assign y313 = ~n3308 ;
  assign y314 = ~n3313 ;
  assign y315 = ~n3318 ;
  assign y316 = ~n3323 ;
  assign y317 = ~n3328 ;
  assign y318 = n3333 ;
  assign y319 = ~n3338 ;
  assign y320 = ~n3343 ;
  assign y321 = ~n3348 ;
  assign y322 = ~n3353 ;
  assign y323 = n3358 ;
  assign y324 = ~n3363 ;
  assign y325 = ~n3368 ;
  assign y326 = ~n3373 ;
  assign y327 = ~n3378 ;
  assign y328 = ~n3383 ;
  assign y329 = ~n3388 ;
  assign y330 = ~n3393 ;
  assign y331 = n3398 ;
  assign y332 = ~n3403 ;
  assign y333 = ~n3408 ;
  assign y334 = ~n3413 ;
  assign y335 = ~n3418 ;
  assign y336 = ~n3423 ;
  assign y337 = ~n3428 ;
  assign y338 = ~n3433 ;
  assign y339 = ~n3438 ;
  assign y340 = ~n3443 ;
  assign y341 = ~n3448 ;
  assign y342 = ~n3453 ;
  assign y343 = ~n3458 ;
  assign y344 = ~n3463 ;
  assign y345 = ~n3468 ;
  assign y346 = n3473 ;
  assign y347 = ~n3478 ;
  assign y348 = ~n3483 ;
  assign y349 = ~n3488 ;
  assign y350 = ~n3493 ;
  assign y351 = ~n3498 ;
  assign y352 = n3504 ;
  assign y353 = n3509 ;
  assign y354 = ~n3514 ;
  assign y355 = n3522 ;
  assign y356 = n3527 ;
  assign y357 = n3532 ;
  assign y358 = ~n3550 ;
  assign y359 = ~n3556 ;
  assign y360 = ~n3562 ;
  assign y361 = ~n3574 ;
  assign y362 = ~n3579 ;
  assign y363 = ~n3585 ;
  assign y364 = ~n3590 ;
  assign y365 = ~n3595 ;
  assign y366 = ~n3600 ;
  assign y367 = n3607 ;
  assign y368 = n3612 ;
  assign y369 = ~n3617 ;
  assign y370 = ~n3622 ;
  assign y371 = ~n3627 ;
  assign y372 = n3632 ;
  assign y373 = n3637 ;
  assign y374 = ~n3642 ;
  assign y375 = ~n3647 ;
  assign y376 = n3652 ;
  assign y377 = ~n3657 ;
  assign y378 = n3662 ;
  assign y379 = n3667 ;
  assign y380 = n3672 ;
  assign y381 = n3677 ;
  assign y382 = n1496 ;
  assign y383 = n3683 ;
  assign y384 = ~n3689 ;
  assign y385 = n3697 ;
  assign y386 = x232 ;
  assign y387 = n3156 ;
  assign y388 = x236 ;
  assign y389 = n3700 ;
  assign y390 = ~n3780 ;
  assign y391 = n3806 ;
  assign y392 = n3834 ;
  assign y393 = n3680 ;
  assign y394 = ~n3872 ;
  assign y395 = n3885 ;
  assign y396 = n3894 ;
  assign y397 = n3916 ;
  assign y398 = n3926 ;
  assign y399 = n3945 ;
  assign y400 = ~n3975 ;
  assign y401 = n3984 ;
  assign y402 = n3996 ;
  assign y403 = n4006 ;
  assign y404 = n4011 ;
  assign y405 = n4021 ;
  assign y406 = n4026 ;
  assign y407 = n4029 ;
  assign y408 = n4037 ;
  assign y409 = n4041 ;
  assign y410 = n4049 ;
  assign y411 = n4057 ;
  assign y412 = n4062 ;
  assign y413 = n4067 ;
  assign y414 = n4073 ;
  assign y415 = n4078 ;
  assign y416 = n4083 ;
  assign y417 = n4088 ;
  assign y418 = n4093 ;
  assign y419 = ~n4100 ;
  assign y420 = ~n4108 ;
  assign y421 = ~n4119 ;
  assign y422 = ~n4128 ;
  assign y423 = n4137 ;
  assign y424 = n4145 ;
  assign y425 = n4153 ;
  assign y426 = ~n4162 ;
  assign y427 = ~n4171 ;
  assign y428 = n4179 ;
  assign y429 = n4187 ;
  assign y430 = n4195 ;
  assign y431 = ~n4204 ;
  assign y432 = n4212 ;
  assign y433 = n4220 ;
  assign y434 = ~n4229 ;
  assign y435 = n4238 ;
  assign y436 = n4247 ;
  assign y437 = ~n4256 ;
  assign y438 = ~n4265 ;
  assign y439 = ~n4274 ;
  assign y440 = n4282 ;
  assign y441 = ~n4286 ;
  assign y442 = n4300 ;
  assign y443 = n4304 ;
  assign y444 = ~n4306 ;
  assign y445 = n4309 ;
  assign y446 = n4314 ;
  assign y447 = n4317 ;
  assign y448 = n4320 ;
  assign y449 = n4323 ;
  assign y450 = n4326 ;
  assign y451 = n4329 ;
  assign y452 = n4332 ;
  assign y453 = n4335 ;
  assign y454 = n4338 ;
  assign y455 = n4341 ;
  assign y456 = n4343 ;
  assign y457 = n4348 ;
  assign y458 = ~n4352 ;
  assign y459 = ~n4360 ;
  assign y460 = n4363 ;
  assign y461 = n4366 ;
  assign y462 = n4369 ;
  assign y463 = n4372 ;
  assign y464 = n4375 ;
  assign y465 = n4378 ;
  assign y466 = n4381 ;
  assign y467 = ~n4389 ;
  assign y468 = ~n4393 ;
  assign y469 = n4396 ;
  assign y470 = n4402 ;
  assign y471 = ~n4404 ;
  assign y472 = n4408 ;
  assign y473 = n4411 ;
  assign y474 = n4415 ;
  assign y475 = n4419 ;
  assign y476 = n4422 ;
  assign y477 = n4425 ;
  assign y478 = n4428 ;
  assign y479 = n4431 ;
  assign y480 = n4434 ;
  assign y481 = n4437 ;
  assign y482 = n4440 ;
  assign y483 = n4443 ;
  assign y484 = n4446 ;
  assign y485 = n4449 ;
  assign y486 = n4452 ;
  assign y487 = n4455 ;
  assign y488 = n4457 ;
  assign y489 = n4466 ;
  assign y490 = n4469 ;
  assign y491 = n4472 ;
  assign y492 = n4475 ;
  assign y493 = n4478 ;
  assign y494 = n4481 ;
  assign y495 = n4484 ;
  assign y496 = n4487 ;
  assign y497 = ~n4490 ;
  assign y498 = n4492 ;
  assign y499 = n4495 ;
  assign y500 = n4498 ;
  assign y501 = n4501 ;
  assign y502 = n4504 ;
  assign y503 = n4507 ;
  assign y504 = n4510 ;
  assign y505 = n4513 ;
  assign y506 = n4516 ;
  assign y507 = n4519 ;
  assign y508 = n4522 ;
  assign y509 = n4525 ;
  assign y510 = n4528 ;
  assign y511 = n4531 ;
  assign y512 = n4534 ;
  assign y513 = n4537 ;
  assign y514 = n4540 ;
  assign y515 = n4543 ;
  assign y516 = n4546 ;
  assign y517 = n4549 ;
  assign y518 = n4552 ;
  assign y519 = n4555 ;
  assign y520 = n4558 ;
  assign y521 = n4561 ;
  assign y522 = n4564 ;
  assign y523 = n4567 ;
  assign y524 = n4570 ;
  assign y525 = n4573 ;
  assign y526 = n4576 ;
  assign y527 = n4579 ;
  assign y528 = n4582 ;
  assign y529 = n4585 ;
  assign y530 = n4588 ;
  assign y531 = n4591 ;
  assign y532 = n4594 ;
  assign y533 = n4597 ;
  assign y534 = n4600 ;
  assign y535 = n4603 ;
  assign y536 = n4606 ;
  assign y537 = n4609 ;
  assign y538 = n4612 ;
  assign y539 = n4615 ;
  assign y540 = n4618 ;
  assign y541 = n4621 ;
  assign y542 = n4624 ;
  assign y543 = n4627 ;
  assign y544 = n4630 ;
  assign y545 = n4633 ;
  assign y546 = n4636 ;
  assign y547 = n4639 ;
  assign y548 = n4642 ;
  assign y549 = n4645 ;
  assign y550 = n4648 ;
  assign y551 = n4651 ;
  assign y552 = n4654 ;
  assign y553 = n4657 ;
  assign y554 = n4660 ;
  assign y555 = n4663 ;
  assign y556 = n4666 ;
  assign y557 = n4669 ;
  assign y558 = n4672 ;
  assign y559 = n4675 ;
  assign y560 = n4678 ;
  assign y561 = n4681 ;
  assign y562 = n4684 ;
  assign y563 = n4687 ;
  assign y564 = n4690 ;
  assign y565 = n4693 ;
  assign y566 = n4696 ;
  assign y567 = n4699 ;
  assign y568 = n4702 ;
  assign y569 = n4705 ;
  assign y570 = n4708 ;
  assign y571 = n4712 ;
  assign y572 = n4715 ;
  assign y573 = n4718 ;
  assign y574 = n4721 ;
  assign y575 = n4724 ;
  assign y576 = n4727 ;
  assign y577 = n4730 ;
  assign y578 = n4733 ;
  assign y579 = n4736 ;
  assign y580 = n4739 ;
  assign y581 = n4742 ;
  assign y582 = n4745 ;
  assign y583 = n4748 ;
  assign y584 = n4751 ;
  assign y585 = n4754 ;
  assign y586 = n4757 ;
  assign y587 = n4760 ;
  assign y588 = n4763 ;
  assign y589 = n4766 ;
  assign y590 = n4769 ;
  assign y591 = n4772 ;
  assign y592 = n4775 ;
  assign y593 = n4778 ;
  assign y594 = n4781 ;
  assign y595 = n4784 ;
  assign y596 = n4787 ;
  assign y597 = n4790 ;
  assign y598 = n4793 ;
  assign y599 = n4796 ;
  assign y600 = n4799 ;
  assign y601 = n4802 ;
  assign y602 = n4805 ;
  assign y603 = n4808 ;
  assign y604 = n4811 ;
  assign y605 = n4814 ;
  assign y606 = n4817 ;
  assign y607 = n4820 ;
  assign y608 = n4823 ;
  assign y609 = n4826 ;
  assign y610 = n4829 ;
  assign y611 = n4832 ;
  assign y612 = n4835 ;
  assign y613 = n4838 ;
  assign y614 = n4861 ;
  assign y615 = n4864 ;
  assign y616 = n4867 ;
  assign y617 = n4870 ;
  assign y618 = n4873 ;
  assign y619 = n4876 ;
  assign y620 = n4879 ;
  assign y621 = n4882 ;
  assign y622 = n4887 ;
  assign y623 = n4892 ;
  assign y624 = n4898 ;
  assign y625 = n4901 ;
  assign y626 = n4906 ;
  assign y627 = n4911 ;
  assign y628 = n4916 ;
  assign y629 = n4921 ;
  assign y630 = n4926 ;
  assign y631 = n4931 ;
  assign y632 = n4936 ;
  assign y633 = n4939 ;
  assign y634 = ~n4399 ;
  assign y635 = n4940 ;
  assign y636 = x583 ;
  assign y637 = n4287 ;
  assign y638 = n4943 ;
  assign y639 = n4946 ;
  assign y640 = n4949 ;
  assign y641 = n4952 ;
  assign y642 = n4955 ;
  assign y643 = n4958 ;
  assign y644 = n4961 ;
  assign y645 = ~n4964 ;
  assign y646 = n4967 ;
  assign y647 = n4970 ;
  assign y648 = n4973 ;
  assign y649 = n4976 ;
  assign y650 = n4979 ;
  assign y651 = ~n4982 ;
  assign y652 = n4985 ;
  assign y653 = n4988 ;
  assign y654 = ~n4991 ;
  assign y655 = n4994 ;
  assign y656 = n4997 ;
  assign y657 = n5000 ;
  assign y658 = n5003 ;
  assign y659 = n5006 ;
  assign y660 = n5009 ;
  assign y661 = n5012 ;
  assign y662 = n5015 ;
  assign y663 = n5018 ;
  assign y664 = n5021 ;
  assign y665 = n5024 ;
  assign y666 = n5027 ;
  assign y667 = n5030 ;
  assign y668 = n5033 ;
  assign y669 = n5036 ;
  assign y670 = n5039 ;
  assign y671 = n5042 ;
  assign y672 = n5045 ;
  assign y673 = n5048 ;
  assign y674 = n5051 ;
  assign y675 = n5054 ;
  assign y676 = ~n5057 ;
  assign y677 = n5060 ;
  assign y678 = n5063 ;
  assign y679 = n5066 ;
  assign y680 = n5069 ;
  assign y681 = ~n5072 ;
  assign y682 = n5075 ;
  assign y683 = n5078 ;
  assign y684 = n5081 ;
  assign y685 = n5084 ;
  assign y686 = n5087 ;
  assign y687 = n5090 ;
  assign y688 = n5093 ;
  assign y689 = n5096 ;
  assign y690 = n5099 ;
  assign y691 = ~n5102 ;
  assign y692 = n5105 ;
  assign y693 = n5108 ;
  assign y694 = n5111 ;
  assign y695 = n5114 ;
  assign y696 = n5117 ;
  assign y697 = n5120 ;
  assign y698 = n5123 ;
  assign y699 = n5126 ;
  assign y700 = n5129 ;
  assign y701 = n5132 ;
  assign y702 = n5135 ;
  assign y703 = n5138 ;
  assign y704 = n5141 ;
  assign y705 = n5144 ;
  assign y706 = n5147 ;
  assign y707 = ~n5150 ;
  assign y708 = n5153 ;
  assign y709 = n5156 ;
  assign y710 = n5159 ;
  assign y711 = n5162 ;
  assign y712 = n5165 ;
  assign y713 = n5168 ;
  assign y714 = n5171 ;
  assign y715 = n5174 ;
  assign y716 = n5177 ;
  assign y717 = n5180 ;
  assign y718 = n5183 ;
  assign y719 = n5186 ;
  assign y720 = n5189 ;
  assign y721 = n5192 ;
  assign y722 = n5195 ;
  assign y723 = n5198 ;
  assign y724 = n5205 ;
  assign y725 = n5208 ;
  assign y726 = ~n5211 ;
  assign y727 = n5214 ;
  assign y728 = n5217 ;
  assign y729 = n5220 ;
  assign y730 = n5223 ;
  assign y731 = n5226 ;
  assign y732 = n5229 ;
  assign y733 = n5232 ;
  assign y734 = n5235 ;
  assign y735 = n5238 ;
  assign y736 = n5241 ;
  assign y737 = n5244 ;
  assign y738 = n5247 ;
  assign y739 = n5250 ;
  assign y740 = n1732 ;
  assign y741 = n5253 ;
  assign y742 = n5256 ;
  assign y743 = n5259 ;
  assign y744 = n5262 ;
  assign y745 = n5266 ;
  assign y746 = n5283 ;
  assign y747 = ~n5286 ;
  assign y748 = n5289 ;
  assign y749 = n5292 ;
  assign y750 = n5607 ;
  assign y751 = n5612 ;
  assign y752 = n5616 ;
  assign y753 = n5622 ;
  assign y754 = n5625 ;
  assign y755 = n5631 ;
  assign y756 = n5635 ;
  assign y757 = n5637 ;
  assign y758 = n5640 ;
  assign y759 = n5643 ;
  assign y760 = n5654 ;
  assign y761 = n5661 ;
  assign y762 = ~n5664 ;
  assign y763 = n5670 ;
  assign y764 = n5673 ;
  assign y765 = n5676 ;
  assign y766 = n5679 ;
  assign y767 = n5682 ;
  assign y768 = n5685 ;
  assign y769 = n5688 ;
  assign y770 = n5691 ;
  assign y771 = n5695 ;
  assign y772 = ~n5700 ;
  assign y773 = n5705 ;
  assign y774 = n5710 ;
  assign y775 = n5713 ;
  assign y776 = n5716 ;
  assign y777 = n5719 ;
  assign y778 = n5722 ;
  assign y779 = n5725 ;
  assign y780 = n5728 ;
  assign y781 = n5734 ;
  assign y782 = n5742 ;
  assign y783 = n5745 ;
  assign y784 = n5748 ;
  assign y785 = n5751 ;
  assign y786 = n5754 ;
  assign y787 = n5757 ;
  assign y788 = ~n5760 ;
  assign y789 = ~n5763 ;
  assign y790 = n5766 ;
  assign y791 = n5769 ;
  assign y792 = ~n5772 ;
  assign y793 = n5775 ;
  assign y794 = n5778 ;
  assign y795 = n5781 ;
  assign y796 = n5784 ;
  assign y797 = n5787 ;
  assign y798 = n5790 ;
  assign y799 = n5793 ;
  assign y800 = n5796 ;
  assign y801 = n5799 ;
  assign y802 = n5802 ;
  assign y803 = ~n5805 ;
  assign y804 = n5808 ;
  assign y805 = n5811 ;
  assign y806 = ~n5814 ;
  assign y807 = ~n5817 ;
  assign y808 = n5820 ;
  assign y809 = n5823 ;
  assign y810 = n5826 ;
  assign y811 = ~n5829 ;
  assign y812 = ~n5832 ;
  assign y813 = n5835 ;
  assign y814 = ~n5838 ;
  assign y815 = n5841 ;
  assign y816 = ~n5853 ;
  assign y817 = n5856 ;
  assign y818 = n5859 ;
  assign y819 = n5862 ;
  assign y820 = n5909 ;
  assign y821 = n5935 ;
  assign y822 = n5938 ;
  assign y823 = n5964 ;
  assign y824 = n5992 ;
  assign y825 = n6018 ;
  assign y826 = ~n6021 ;
  assign y827 = n6042 ;
  assign y828 = n6063 ;
  assign y829 = n6089 ;
  assign y830 = n6114 ;
  assign y831 = n6140 ;
  assign y832 = n6165 ;
  assign y833 = n6190 ;
  assign y834 = n6211 ;
  assign y835 = n6232 ;
  assign y836 = n6258 ;
  assign y837 = n6261 ;
  assign y838 = n6264 ;
  assign y839 = n6285 ;
  assign y840 = n1470 ;
  assign y841 = ~n6289 ;
  assign y842 = n6316 ;
  assign y843 = ~n6319 ;
  assign y844 = n6322 ;
  assign y845 = ~n6325 ;
  assign y846 = n6350 ;
  assign y847 = n6353 ;
  assign y848 = n6356 ;
  assign y849 = n6379 ;
  assign y850 = ~n6382 ;
  assign y851 = ~n6385 ;
  assign y852 = ~n6388 ;
  assign y853 = n6391 ;
  assign y854 = ~n6394 ;
  assign y855 = ~n6397 ;
  assign y856 = n6400 ;
  assign y857 = n6403 ;
  assign y858 = ~n6406 ;
  assign y859 = ~n6409 ;
  assign y860 = n6412 ;
  assign y861 = ~n6415 ;
  assign y862 = n6418 ;
  assign y863 = n6421 ;
  assign y864 = n6444 ;
  assign y865 = n6467 ;
  assign y866 = ~n6470 ;
  assign y867 = n6473 ;
  assign y868 = n6496 ;
  assign y869 = n6519 ;
  assign y870 = n6542 ;
  assign y871 = n6567 ;
  assign y872 = n6570 ;
  assign y873 = n6593 ;
  assign y874 = n6618 ;
  assign y875 = n6641 ;
  assign y876 = n6666 ;
  assign y877 = n6691 ;
  assign y878 = n6723 ;
  assign y879 = n6748 ;
  assign y880 = ~n6751 ;
  assign y881 = ~n6754 ;
  assign y882 = ~n6757 ;
  assign y883 = n6760 ;
  assign y884 = n6763 ;
  assign y885 = ~n6766 ;
  assign y886 = n6769 ;
  assign y887 = n6772 ;
  assign y888 = n6775 ;
  assign y889 = ~n6778 ;
  assign y890 = n6801 ;
  assign y891 = ~n6804 ;
  assign y892 = n6807 ;
  assign y893 = n6810 ;
  assign y894 = ~n6813 ;
  assign y895 = ~n6816 ;
  assign y896 = n6820 ;
  assign y897 = n5650 ;
  assign y898 = ~n6823 ;
  assign y899 = ~n6826 ;
  assign y900 = n6829 ;
  assign y901 = ~n6832 ;
  assign y902 = ~n6835 ;
  assign y903 = n6838 ;
  assign y904 = n6840 ;
  assign y905 = n6843 ;
  assign y906 = n6846 ;
  assign y907 = ~n6849 ;
  assign y908 = ~n6852 ;
  assign y909 = ~n6855 ;
  assign y910 = ~n6858 ;
  assign y911 = ~n6861 ;
  assign y912 = ~n6864 ;
  assign y913 = ~n6867 ;
  assign y914 = ~n6870 ;
  assign y915 = n6873 ;
  assign y916 = n6876 ;
  assign y917 = ~n6879 ;
  assign y918 = ~n6882 ;
  assign y919 = ~n6885 ;
  assign y920 = n6888 ;
  assign y921 = n6891 ;
  assign y922 = ~n6902 ;
  assign y923 = n6905 ;
  assign y924 = ~n6908 ;
  assign y925 = ~n6911 ;
  assign y926 = n6913 ;
  assign y927 = ~n6916 ;
  assign y928 = n6919 ;
  assign y929 = n6922 ;
  assign y930 = n6924 ;
  assign y931 = ~n6927 ;
  assign y932 = n6935 ;
  assign y933 = ~n6938 ;
  assign y934 = ~n6941 ;
  assign y935 = n6949 ;
  assign y936 = ~n6950 ;
  assign y937 = ~n6951 ;
  assign y938 = n6954 ;
  assign y939 = ~n6956 ;
  assign y940 = n6959 ;
  assign y941 = n6962 ;
  assign y942 = n6965 ;
  assign y943 = ~n6967 ;
  assign y944 = n6970 ;
  assign y945 = n6973 ;
  assign y946 = n6976 ;
  assign y947 = n6979 ;
  assign y948 = n6982 ;
  assign y949 = n6985 ;
  assign y950 = ~n1691 ;
  assign y951 = n6989 ;
  assign y952 = n6992 ;
  assign y953 = ~n6999 ;
  assign y954 = n5739 ;
  assign y955 = n7002 ;
  assign y956 = ~n7005 ;
  assign y957 = n7008 ;
  assign y958 = n7011 ;
  assign y959 = n5851 ;
  assign y960 = ~n7014 ;
  assign y961 = n7017 ;
  assign y962 = ~n7021 ;
  assign y963 = n6899 ;
  assign y964 = n7024 ;
  assign y965 = n7027 ;
  assign y966 = ~n7030 ;
  assign y967 = n7033 ;
  assign y968 = n7036 ;
  assign y969 = ~n7039 ;
  assign y970 = n7042 ;
  assign y971 = ~n7045 ;
  assign y972 = n7048 ;
  assign y973 = n7051 ;
  assign y974 = ~n7053 ;
  assign y975 = n2914 ;
  assign y976 = ~n7055 ;
  assign y977 = ~n7058 ;
  assign y978 = ~n6714 ;
  assign y979 = ~n7059 ;
  assign y980 = n6286 ;
  assign y981 = n7063 ;
  assign y982 = n7078 ;
  assign y983 = n7091 ;
  assign y984 = n7104 ;
  assign y985 = n7117 ;
  assign y986 = n7120 ;
  assign y987 = ~n7123 ;
  assign y988 = n6817 ;
  assign y989 = n7125 ;
  assign y990 = n7127 ;
  assign y991 = n7128 ;
  assign y992 = ~n7132 ;
  assign y993 = n7135 ;
  assign y994 = n7138 ;
  assign y995 = n7141 ;
  assign y996 = n7144 ;
  assign y997 = ~n2193 ;
  assign y998 = n7147 ;
  assign y999 = n7150 ;
  assign y1000 = n7153 ;
  assign y1001 = n7156 ;
  assign y1002 = n7159 ;
  assign y1003 = n7162 ;
  assign y1004 = n7165 ;
  assign y1005 = n7168 ;
  assign y1006 = n7171 ;
  assign y1007 = n7174 ;
  assign y1008 = n7177 ;
  assign y1009 = n7180 ;
  assign y1010 = n7183 ;
  assign y1011 = n7186 ;
  assign y1012 = n7189 ;
  assign y1013 = n7192 ;
  assign y1014 = n7195 ;
  assign y1015 = n7198 ;
  assign y1016 = n7201 ;
  assign y1017 = n7204 ;
  assign y1018 = n7207 ;
  assign y1019 = n7210 ;
  assign y1020 = n7213 ;
  assign y1021 = n7216 ;
  assign y1022 = n7219 ;
  assign y1023 = n7222 ;
  assign y1024 = n7225 ;
  assign y1025 = n7228 ;
  assign y1026 = n7231 ;
  assign y1027 = n7234 ;
  assign y1028 = n7237 ;
  assign y1029 = n7240 ;
  assign y1030 = n7243 ;
  assign y1031 = n7246 ;
  assign y1032 = n7249 ;
  assign y1033 = n7252 ;
  assign y1034 = n7255 ;
  assign y1035 = n7258 ;
  assign y1036 = n7261 ;
  assign y1037 = n7264 ;
  assign y1038 = n1380 ;
  assign y1039 = n7267 ;
  assign y1040 = n7270 ;
  assign y1041 = n7273 ;
  assign y1042 = n7276 ;
  assign y1043 = n7279 ;
  assign y1044 = n7282 ;
  assign y1045 = n7285 ;
  assign y1046 = n7288 ;
  assign y1047 = n7291 ;
  assign y1048 = n7294 ;
  assign y1049 = n1211 ;
  assign y1050 = n7297 ;
  assign y1051 = n7300 ;
  assign y1052 = n7303 ;
  assign y1053 = x67 ;
  assign y1054 = n7306 ;
  assign y1055 = n7309 ;
  assign y1056 = n7312 ;
  assign y1057 = n1726 ;
  assign y1058 = n7315 ;
  assign y1059 = n7318 ;
  assign y1060 = n7321 ;
  assign y1061 = n7324 ;
  assign y1062 = n7327 ;
  assign y1063 = n7335 ;
  assign y1064 = n7338 ;
  assign y1065 = n7341 ;
  assign y1066 = n7344 ;
  assign y1067 = n7347 ;
  assign y1068 = n7350 ;
  assign y1069 = n7353 ;
  assign y1070 = ~n7355 ;
  assign y1071 = n7358 ;
  assign y1072 = n7361 ;
  assign y1073 = n7364 ;
  assign y1074 = n7367 ;
  assign y1075 = n7370 ;
  assign y1076 = n7373 ;
  assign y1077 = n7376 ;
  assign y1078 = n7379 ;
  assign y1079 = n7382 ;
  assign y1080 = n7385 ;
  assign y1081 = n7388 ;
  assign y1082 = n7391 ;
  assign y1083 = n7394 ;
  assign y1084 = n7397 ;
  assign y1085 = n7400 ;
  assign y1086 = n7403 ;
  assign y1087 = n7406 ;
  assign y1088 = n7409 ;
  assign y1089 = n7412 ;
  assign y1090 = n7415 ;
  assign y1091 = n7418 ;
  assign y1092 = n7421 ;
  assign y1093 = n7424 ;
  assign y1094 = n7427 ;
  assign y1095 = n7430 ;
  assign y1096 = n7433 ;
  assign y1097 = n7436 ;
  assign y1098 = n7439 ;
  assign y1099 = n7442 ;
  assign y1100 = n7445 ;
  assign y1101 = n1660 ;
  assign y1102 = n5199 ;
  assign y1103 = n7448 ;
  assign y1104 = n7450 ;
  assign y1105 = ~n7452 ;
  assign y1106 = n7453 ;
  assign y1107 = n1465 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n7455 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n7456 ;
  assign y1116 = n7457 ;
  assign y1117 = x1014 ;
  assign y1118 = n7458 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n7459 ;
  assign y1123 = x1135 ;
  assign y1124 = n7460 ;
  assign y1125 = n7461 ;
  assign y1126 = n7462 ;
  assign y1127 = n7463 ;
  assign y1128 = n7464 ;
  assign y1129 = n7465 ;
  assign y1130 = ~x278 ;
  assign y1131 = n7466 ;
  assign y1132 = n7467 ;
  assign y1133 = ~n7468 ;
  assign y1134 = x1064 ;
  assign y1135 = n1689 ;
  assign y1136 = x299 ;
  assign y1137 = n7469 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
