module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 ;
  assign n129 = x0 & x64 ;
  assign n130 = x0 & ~x65 ;
  assign n131 = x1 & x64 ;
  assign n132 = ( x0 & n130 ) | ( x0 & n131 ) | ( n130 & n131 ) ;
  assign n133 = ( x0 & ~n130 ) | ( x0 & n131 ) | ( ~n130 & n131 ) ;
  assign n134 = ( n130 & ~n132 ) | ( n130 & n133 ) | ( ~n132 & n133 ) ;
  assign n135 = ~x1 & x2 ;
  assign n136 = ~x0 & n135 ;
  assign n137 = x64 & n136 ;
  assign n138 = ~x64 & x65 ;
  assign n139 = x66 | n138 ;
  assign n140 = x0 & ~n139 ;
  assign n141 = x1 & x65 ;
  assign n142 = x0 | n141 ;
  assign n143 = ( n137 & ~n140 ) | ( n137 & n142 ) | ( ~n140 & n142 ) ;
  assign n144 = x1 & x2 ;
  assign n145 = ( x1 & n135 ) | ( x1 & ~n144 ) | ( n135 & ~n144 ) ;
  assign n146 = x0 & n145 ;
  assign n147 = x0 & ~n146 ;
  assign n148 = x65 & x66 ;
  assign n149 = ~x64 & n148 ;
  assign n150 = n147 | n149 ;
  assign n151 = x66 & ~n146 ;
  assign n152 = n150 & ~n151 ;
  assign n153 = n143 & ~n152 ;
  assign n154 = n129 | n134 ;
  assign n155 = x2 & n154 ;
  assign n156 = n153 & n155 ;
  assign n157 = n153 | n155 ;
  assign n158 = ~n156 & n157 ;
  assign n159 = x2 & x3 ;
  assign n160 = ~x2 & x3 ;
  assign n161 = ( x2 & ~n159 ) | ( x2 & n160 ) | ( ~n159 & n160 ) ;
  assign n162 = x64 & n161 ;
  assign n163 = x2 & ~n157 ;
  assign n164 = n162 | n163 ;
  assign n165 = x64 & x65 ;
  assign n166 = ( x65 & x66 ) | ( x65 & n165 ) | ( x66 & n165 ) ;
  assign n167 = ( x66 & x67 ) | ( x66 & n166 ) | ( x67 & n166 ) ;
  assign n168 = ( ~x66 & x67 ) | ( ~x66 & n166 ) | ( x67 & n166 ) ;
  assign n169 = ( x66 & ~n167 ) | ( x66 & n168 ) | ( ~n167 & n168 ) ;
  assign n170 = x0 & n169 ;
  assign n171 = ( x1 & x2 ) | ( x1 & n170 ) | ( x2 & n170 ) ;
  assign n172 = ~x0 & x1 ;
  assign n173 = x66 & n172 ;
  assign n174 = x0 & n135 ;
  assign n175 = ( ~x65 & n135 ) | ( ~x65 & n174 ) | ( n135 & n174 ) ;
  assign n176 = n173 | n175 ;
  assign n177 = x67 & n147 ;
  assign n178 = n176 | n177 ;
  assign n179 = ~n171 & n178 ;
  assign n180 = n171 & ~n178 ;
  assign n181 = n179 | n180 ;
  assign n182 = n164 | n181 ;
  assign n183 = n164 & n181 ;
  assign n184 = n182 & ~n183 ;
  assign n185 = x66 & n136 ;
  assign n186 = x67 & n172 ;
  assign n187 = ( x0 & x68 ) | ( x0 & n146 ) | ( x68 & n146 ) ;
  assign n188 = ~x67 & n148 ;
  assign n189 = ~x68 & n188 ;
  assign n190 = ~n166 & n168 ;
  assign n191 = ( x68 & n188 ) | ( x68 & n190 ) | ( n188 & n190 ) ;
  assign n192 = x68 | n190 ;
  assign n193 = ( n189 & ~n191 ) | ( n189 & n192 ) | ( ~n191 & n192 ) ;
  assign n194 = n146 & ~n193 ;
  assign n195 = ( n186 & n187 ) | ( n186 & ~n194 ) | ( n187 & ~n194 ) ;
  assign n196 = ( x2 & ~n185 ) | ( x2 & n195 ) | ( ~n185 & n195 ) ;
  assign n197 = ( x2 & n185 ) | ( x2 & n195 ) | ( n185 & n195 ) ;
  assign n198 = n196 & ~n197 ;
  assign n199 = ~x2 & x4 ;
  assign n200 = x3 & x4 ;
  assign n201 = ( n159 & n199 ) | ( n159 & ~n200 ) | ( n199 & ~n200 ) ;
  assign n202 = x65 & ~n201 ;
  assign n203 = x4 | x5 ;
  assign n204 = x4 & x5 ;
  assign n205 = ( n161 & ~n203 ) | ( n161 & n204 ) | ( ~n203 & n204 ) ;
  assign n206 = n161 & ~n205 ;
  assign n207 = ( n201 & ~n202 ) | ( n201 & n206 ) | ( ~n202 & n206 ) ;
  assign n208 = ( x65 & n138 ) | ( x65 & n205 ) | ( n138 & n205 ) ;
  assign n209 = n161 & n208 ;
  assign n210 = x64 | n209 ;
  assign n211 = ( n207 & n209 ) | ( n207 & n210 ) | ( n209 & n210 ) ;
  assign n212 = n162 | n211 ;
  assign n213 = ( x5 & n162 ) | ( x5 & ~n211 ) | ( n162 & ~n211 ) ;
  assign n214 = x5 & ~n211 ;
  assign n215 = ( n212 & ~n213 ) | ( n212 & n214 ) | ( ~n213 & n214 ) ;
  assign n216 = ( n183 & ~n198 ) | ( n183 & n215 ) | ( ~n198 & n215 ) ;
  assign n217 = ( n183 & n198 ) | ( n183 & n215 ) | ( n198 & n215 ) ;
  assign n218 = ( n198 & n216 ) | ( n198 & ~n217 ) | ( n216 & ~n217 ) ;
  assign n219 = ~x3 & x5 ;
  assign n220 = ( x2 & x5 ) | ( x2 & n201 ) | ( x5 & n201 ) ;
  assign n221 = ( n159 & n219 ) | ( n159 & ~n220 ) | ( n219 & ~n220 ) ;
  assign n222 = x64 & n221 ;
  assign n223 = x66 & ~n205 ;
  assign n224 = ( x66 & n222 ) | ( x66 & ~n223 ) | ( n222 & ~n223 ) ;
  assign n225 = n139 & ~n149 ;
  assign n226 = ( x66 & ~n148 ) | ( x66 & n225 ) | ( ~n148 & n225 ) ;
  assign n227 = n206 & n226 ;
  assign n228 = ( x65 & n207 ) | ( x65 & n227 ) | ( n207 & n227 ) ;
  assign n229 = n224 | n228 ;
  assign n230 = ~x5 & n229 ;
  assign n231 = ( x5 & n212 ) | ( x5 & n229 ) | ( n212 & n229 ) ;
  assign n232 = n212 & n229 ;
  assign n233 = ( n230 & n231 ) | ( n230 & ~n232 ) | ( n231 & ~n232 ) ;
  assign n234 = x67 & x68 ;
  assign n235 = ( x68 & n148 ) | ( x68 & n234 ) | ( n148 & n234 ) ;
  assign n236 = ~x69 & n235 ;
  assign n237 = ( x68 & n167 ) | ( x68 & ~n189 ) | ( n167 & ~n189 ) ;
  assign n238 = ( x69 & n235 ) | ( x69 & ~n237 ) | ( n235 & ~n237 ) ;
  assign n239 = ~x69 & n237 ;
  assign n240 = ( ~n236 & n238 ) | ( ~n236 & n239 ) | ( n238 & n239 ) ;
  assign n241 = x0 & n240 ;
  assign n242 = ( x1 & x2 ) | ( x1 & n241 ) | ( x2 & n241 ) ;
  assign n243 = x68 & n172 ;
  assign n244 = ( ~x67 & n135 ) | ( ~x67 & n174 ) | ( n135 & n174 ) ;
  assign n245 = n243 | n244 ;
  assign n246 = x69 & n147 ;
  assign n247 = n245 | n246 ;
  assign n248 = n242 | n247 ;
  assign n249 = n242 & n247 ;
  assign n250 = n248 & ~n249 ;
  assign n251 = ( n217 & n233 ) | ( n217 & n250 ) | ( n233 & n250 ) ;
  assign n252 = ( ~n217 & n233 ) | ( ~n217 & n250 ) | ( n233 & n250 ) ;
  assign n253 = ( n217 & ~n251 ) | ( n217 & n252 ) | ( ~n251 & n252 ) ;
  assign n254 = x67 & n205 ;
  assign n255 = n169 & n206 ;
  assign n256 = n254 | n255 ;
  assign n257 = x66 & n201 ;
  assign n258 = x65 & n221 ;
  assign n259 = n257 | n258 ;
  assign n260 = n256 | n259 ;
  assign n261 = x5 & ~n212 ;
  assign n262 = ~n229 & n261 ;
  assign n263 = x5 | x6 ;
  assign n264 = x5 & x6 ;
  assign n265 = n263 & ~n264 ;
  assign n266 = x64 & n265 ;
  assign n267 = x5 | n266 ;
  assign n268 = n260 & n267 ;
  assign n269 = ~x6 & x64 ;
  assign n270 = ( n260 & n267 ) | ( n260 & ~n269 ) | ( n267 & ~n269 ) ;
  assign n271 = ( n262 & ~n268 ) | ( n262 & n270 ) | ( ~n268 & n270 ) ;
  assign n272 = ( ~n262 & n269 ) | ( ~n262 & n271 ) | ( n269 & n271 ) ;
  assign n273 = ( n260 & n271 ) | ( n260 & n272 ) | ( n271 & n272 ) ;
  assign n274 = ( ~x70 & n235 ) | ( ~x70 & n238 ) | ( n235 & n238 ) ;
  assign n275 = ( x70 & n235 ) | ( x70 & n238 ) | ( n235 & n238 ) ;
  assign n276 = ( x70 & n274 ) | ( x70 & ~n275 ) | ( n274 & ~n275 ) ;
  assign n277 = x0 & n276 ;
  assign n278 = ( x1 & x2 ) | ( x1 & n277 ) | ( x2 & n277 ) ;
  assign n279 = x69 & n172 ;
  assign n280 = ( ~x68 & n135 ) | ( ~x68 & n174 ) | ( n135 & n174 ) ;
  assign n281 = n279 | n280 ;
  assign n282 = x70 & n147 ;
  assign n283 = n281 | n282 ;
  assign n284 = n278 | n283 ;
  assign n285 = n278 & n283 ;
  assign n286 = n284 & ~n285 ;
  assign n287 = ( n251 & n273 ) | ( n251 & n286 ) | ( n273 & n286 ) ;
  assign n288 = ( ~n251 & n273 ) | ( ~n251 & n286 ) | ( n273 & n286 ) ;
  assign n289 = ( n251 & ~n287 ) | ( n251 & n288 ) | ( ~n287 & n288 ) ;
  assign n290 = n262 | n266 ;
  assign n291 = ( n267 & n268 ) | ( n267 & ~n290 ) | ( n268 & ~n290 ) ;
  assign n292 = x68 & n205 ;
  assign n293 = x66 & n221 ;
  assign n294 = n292 | n293 ;
  assign n295 = n193 & n206 ;
  assign n296 = n294 | n295 ;
  assign n297 = x67 & n201 ;
  assign n298 = n296 | n297 ;
  assign n299 = ~x7 & x8 ;
  assign n300 = x7 & ~x8 ;
  assign n301 = ( n265 & n299 ) | ( n265 & n300 ) | ( n299 & n300 ) ;
  assign n302 = ( x64 & n138 ) | ( x64 & ~n165 ) | ( n138 & ~n165 ) ;
  assign n303 = n301 & n302 ;
  assign n304 = ~x5 & x7 ;
  assign n305 = x6 & x7 ;
  assign n306 = ( n264 & n304 ) | ( n264 & ~n305 ) | ( n304 & ~n305 ) ;
  assign n307 = x64 & n306 ;
  assign n308 = n303 | n307 ;
  assign n309 = n265 & ~n301 ;
  assign n310 = x65 & n309 ;
  assign n311 = n308 | n310 ;
  assign n312 = n266 | n311 ;
  assign n313 = ( x8 & n266 ) | ( x8 & ~n311 ) | ( n266 & ~n311 ) ;
  assign n314 = x8 & ~n311 ;
  assign n315 = ( n312 & ~n313 ) | ( n312 & n314 ) | ( ~n313 & n314 ) ;
  assign n316 = ( n291 & n298 ) | ( n291 & n315 ) | ( n298 & n315 ) ;
  assign n317 = ( ~n291 & n298 ) | ( ~n291 & n315 ) | ( n298 & n315 ) ;
  assign n318 = ( n291 & ~n316 ) | ( n291 & n317 ) | ( ~n316 & n317 ) ;
  assign n319 = ( x69 & n237 ) | ( x69 & n275 ) | ( n237 & n275 ) ;
  assign n320 = ( x70 & ~x71 ) | ( x70 & n319 ) | ( ~x71 & n319 ) ;
  assign n321 = ( x70 & x71 ) | ( x70 & ~n319 ) | ( x71 & ~n319 ) ;
  assign n322 = ( ~x70 & n320 ) | ( ~x70 & n321 ) | ( n320 & n321 ) ;
  assign n323 = x0 & n322 ;
  assign n324 = ( x1 & x2 ) | ( x1 & n323 ) | ( x2 & n323 ) ;
  assign n325 = x70 & n172 ;
  assign n326 = ( ~x69 & n135 ) | ( ~x69 & n174 ) | ( n135 & n174 ) ;
  assign n327 = n325 | n326 ;
  assign n328 = x71 & n147 ;
  assign n329 = n327 | n328 ;
  assign n330 = n324 | n329 ;
  assign n331 = n324 & n329 ;
  assign n332 = n330 & ~n331 ;
  assign n333 = ( n287 & n318 ) | ( n287 & n332 ) | ( n318 & n332 ) ;
  assign n334 = ( ~n287 & n318 ) | ( ~n287 & n332 ) | ( n318 & n332 ) ;
  assign n335 = ( n287 & ~n333 ) | ( n287 & n334 ) | ( ~n333 & n334 ) ;
  assign n336 = ( n260 & n298 ) | ( n260 & n315 ) | ( n298 & n315 ) ;
  assign n337 = x5 & n260 ;
  assign n338 = x5 & ~n298 ;
  assign n339 = ( n336 & ~n337 ) | ( n336 & n338 ) | ( ~n337 & n338 ) ;
  assign n340 = n290 & n339 ;
  assign n341 = ( ~n318 & n339 ) | ( ~n318 & n340 ) | ( n339 & n340 ) ;
  assign n342 = n206 & n240 ;
  assign n343 = x5 & n342 ;
  assign n344 = x69 & n205 ;
  assign n345 = x68 & n201 ;
  assign n346 = n344 | n345 ;
  assign n347 = x67 & n221 ;
  assign n348 = n346 | n347 ;
  assign n349 = ( ~x5 & n342 ) | ( ~x5 & n348 ) | ( n342 & n348 ) ;
  assign n350 = x5 & ~n348 ;
  assign n351 = ( ~n343 & n349 ) | ( ~n343 & n350 ) | ( n349 & n350 ) ;
  assign n352 = x66 & n309 ;
  assign n353 = x65 & n306 ;
  assign n354 = n352 | n353 ;
  assign n355 = n226 & n301 ;
  assign n356 = n354 | n355 ;
  assign n357 = n264 & n300 ;
  assign n358 = ~n263 & n299 ;
  assign n359 = n357 | n358 ;
  assign n360 = x64 & n359 ;
  assign n361 = n356 | n360 ;
  assign n362 = ~x8 & n361 ;
  assign n363 = ( x8 & n312 ) | ( x8 & n361 ) | ( n312 & n361 ) ;
  assign n364 = n312 & n361 ;
  assign n365 = ( n362 & n363 ) | ( n362 & ~n364 ) | ( n363 & ~n364 ) ;
  assign n366 = ( n341 & n351 ) | ( n341 & n365 ) | ( n351 & n365 ) ;
  assign n367 = ( ~n341 & n351 ) | ( ~n341 & n365 ) | ( n351 & n365 ) ;
  assign n368 = ( n341 & ~n366 ) | ( n341 & n367 ) | ( ~n366 & n367 ) ;
  assign n369 = ( ~x70 & x72 ) | ( ~x70 & n319 ) | ( x72 & n319 ) ;
  assign n370 = ( x70 & x71 ) | ( x70 & n369 ) | ( x71 & n369 ) ;
  assign n371 = ( x70 & x72 ) | ( x70 & ~n321 ) | ( x72 & ~n321 ) ;
  assign n372 = ( x71 & ~n370 ) | ( x71 & n371 ) | ( ~n370 & n371 ) ;
  assign n373 = x0 & n372 ;
  assign n374 = ( x1 & x2 ) | ( x1 & n373 ) | ( x2 & n373 ) ;
  assign n375 = x71 & n172 ;
  assign n376 = x72 | n375 ;
  assign n377 = ( n147 & n375 ) | ( n147 & n376 ) | ( n375 & n376 ) ;
  assign n378 = ( ~x70 & n135 ) | ( ~x70 & n174 ) | ( n135 & n174 ) ;
  assign n379 = n377 | n378 ;
  assign n380 = n374 | n379 ;
  assign n381 = n374 & n379 ;
  assign n382 = n380 & ~n381 ;
  assign n383 = ( n333 & n368 ) | ( n333 & n382 ) | ( n368 & n382 ) ;
  assign n384 = ( ~n333 & n368 ) | ( ~n333 & n382 ) | ( n368 & n382 ) ;
  assign n385 = ( n333 & ~n383 ) | ( n333 & n384 ) | ( ~n383 & n384 ) ;
  assign n386 = ( x72 & x73 ) | ( x72 & n370 ) | ( x73 & n370 ) ;
  assign n387 = ( x72 & x73 ) | ( x72 & ~n370 ) | ( x73 & ~n370 ) ;
  assign n388 = ( n370 & ~n386 ) | ( n370 & n387 ) | ( ~n386 & n387 ) ;
  assign n389 = x0 & n388 ;
  assign n390 = ( x1 & x2 ) | ( x1 & n389 ) | ( x2 & n389 ) ;
  assign n391 = x73 & n147 ;
  assign n392 = ~x71 & n136 ;
  assign n393 = x72 & n172 ;
  assign n394 = n174 | n393 ;
  assign n395 = n392 | n394 ;
  assign n396 = n391 | n395 ;
  assign n397 = n390 | n396 ;
  assign n398 = n390 & n396 ;
  assign n399 = n397 & ~n398 ;
  assign n400 = n312 | n361 ;
  assign n401 = x8 & n400 ;
  assign n402 = x66 & n306 ;
  assign n403 = n169 & n301 ;
  assign n404 = x67 & n309 ;
  assign n405 = x65 & ~n359 ;
  assign n406 = ( x65 & n404 ) | ( x65 & ~n405 ) | ( n404 & ~n405 ) ;
  assign n407 = n403 | n406 ;
  assign n408 = n402 | n407 ;
  assign n409 = x8 | x9 ;
  assign n410 = x8 & x9 ;
  assign n411 = n409 & ~n410 ;
  assign n412 = x64 & n411 ;
  assign n413 = ( n401 & ~n408 ) | ( n401 & n412 ) | ( ~n408 & n412 ) ;
  assign n414 = x8 & ~n408 ;
  assign n415 = ( ~n401 & n408 ) | ( ~n401 & n414 ) | ( n408 & n414 ) ;
  assign n416 = ( n412 & n414 ) | ( n412 & n415 ) | ( n414 & n415 ) ;
  assign n417 = ( n413 & n415 ) | ( n413 & ~n416 ) | ( n415 & ~n416 ) ;
  assign n418 = n206 & n276 ;
  assign n419 = x5 & n418 ;
  assign n420 = x70 & n205 ;
  assign n421 = x69 & n201 ;
  assign n422 = n420 | n421 ;
  assign n423 = x68 & n221 ;
  assign n424 = n422 | n423 ;
  assign n425 = ( ~x5 & n418 ) | ( ~x5 & n424 ) | ( n418 & n424 ) ;
  assign n426 = x5 & ~n424 ;
  assign n427 = ( ~n419 & n425 ) | ( ~n419 & n426 ) | ( n425 & n426 ) ;
  assign n428 = ( n366 & ~n417 ) | ( n366 & n427 ) | ( ~n417 & n427 ) ;
  assign n429 = ( n366 & n417 ) | ( n366 & n427 ) | ( n417 & n427 ) ;
  assign n430 = ( n417 & n428 ) | ( n417 & ~n429 ) | ( n428 & ~n429 ) ;
  assign n431 = ( n383 & n399 ) | ( n383 & n430 ) | ( n399 & n430 ) ;
  assign n432 = ( ~n383 & n399 ) | ( ~n383 & n430 ) | ( n399 & n430 ) ;
  assign n433 = ( n383 & ~n431 ) | ( n383 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = ( ~x72 & x74 ) | ( ~x72 & n387 ) | ( x74 & n387 ) ;
  assign n435 = ( x72 & x74 ) | ( x72 & n387 ) | ( x74 & n387 ) ;
  assign n436 = ( x72 & n434 ) | ( x72 & ~n435 ) | ( n434 & ~n435 ) ;
  assign n437 = x0 & n436 ;
  assign n438 = ( x1 & x2 ) | ( x1 & n437 ) | ( x2 & n437 ) ;
  assign n439 = x73 & n172 ;
  assign n440 = x74 | n439 ;
  assign n441 = ( n147 & n439 ) | ( n147 & n440 ) | ( n439 & n440 ) ;
  assign n442 = ( ~x72 & n135 ) | ( ~x72 & n174 ) | ( n135 & n174 ) ;
  assign n443 = n441 | n442 ;
  assign n444 = n438 | n443 ;
  assign n445 = n438 & n443 ;
  assign n446 = n444 & ~n445 ;
  assign n447 = ~x10 & x11 ;
  assign n448 = x10 & ~x11 ;
  assign n449 = ( n411 & n447 ) | ( n411 & n448 ) | ( n447 & n448 ) ;
  assign n450 = n302 & n449 ;
  assign n451 = ~x8 & x10 ;
  assign n452 = x9 & x10 ;
  assign n453 = ( n410 & n451 ) | ( n410 & ~n452 ) | ( n451 & ~n452 ) ;
  assign n454 = x64 & n453 ;
  assign n455 = n450 | n454 ;
  assign n456 = n411 & ~n449 ;
  assign n457 = x65 & n456 ;
  assign n458 = n455 | n457 ;
  assign n459 = n412 | n458 ;
  assign n460 = ( x11 & n412 ) | ( x11 & ~n458 ) | ( n412 & ~n458 ) ;
  assign n461 = x11 & ~n458 ;
  assign n462 = ( n459 & ~n460 ) | ( n459 & n461 ) | ( ~n460 & n461 ) ;
  assign n463 = x68 & n309 ;
  assign n464 = x8 & n463 ;
  assign n465 = x67 & n306 ;
  assign n466 = x66 & n359 ;
  assign n467 = n465 | n466 ;
  assign n468 = n193 & n301 ;
  assign n469 = n467 | n468 ;
  assign n470 = ( ~x8 & n463 ) | ( ~x8 & n469 ) | ( n463 & n469 ) ;
  assign n471 = x8 & ~n469 ;
  assign n472 = ( ~n464 & n470 ) | ( ~n464 & n471 ) | ( n470 & n471 ) ;
  assign n473 = ( n416 & ~n462 ) | ( n416 & n472 ) | ( ~n462 & n472 ) ;
  assign n474 = ( n416 & n462 ) | ( n416 & n472 ) | ( n462 & n472 ) ;
  assign n475 = ( n462 & n473 ) | ( n462 & ~n474 ) | ( n473 & ~n474 ) ;
  assign n476 = n206 & n322 ;
  assign n477 = x5 & n476 ;
  assign n478 = x71 & n205 ;
  assign n479 = x70 & n201 ;
  assign n480 = n478 | n479 ;
  assign n481 = x69 & n221 ;
  assign n482 = n480 | n481 ;
  assign n483 = ( ~x5 & n476 ) | ( ~x5 & n482 ) | ( n476 & n482 ) ;
  assign n484 = x5 & ~n482 ;
  assign n485 = ( ~n477 & n483 ) | ( ~n477 & n484 ) | ( n483 & n484 ) ;
  assign n486 = ( n429 & ~n475 ) | ( n429 & n485 ) | ( ~n475 & n485 ) ;
  assign n487 = ( n429 & n475 ) | ( n429 & n485 ) | ( n475 & n485 ) ;
  assign n488 = ( n475 & n486 ) | ( n475 & ~n487 ) | ( n486 & ~n487 ) ;
  assign n489 = ( ~n431 & n446 ) | ( ~n431 & n488 ) | ( n446 & n488 ) ;
  assign n490 = ( n431 & n446 ) | ( n431 & n488 ) | ( n446 & n488 ) ;
  assign n491 = ( n431 & n489 ) | ( n431 & ~n490 ) | ( n489 & ~n490 ) ;
  assign n492 = x74 & ~x75 ;
  assign n493 = x72 & ~x73 ;
  assign n494 = ( x73 & x74 ) | ( x73 & ~n493 ) | ( x74 & ~n493 ) ;
  assign n495 = x72 & ~x74 ;
  assign n496 = ( x73 & n493 ) | ( x73 & ~n495 ) | ( n493 & ~n495 ) ;
  assign n497 = ( x75 & n494 ) | ( x75 & ~n496 ) | ( n494 & ~n496 ) ;
  assign n498 = x73 & ~n497 ;
  assign n499 = x74 & n493 ;
  assign n500 = ( ~n492 & n498 ) | ( ~n492 & n499 ) | ( n498 & n499 ) ;
  assign n501 = n370 & n500 ;
  assign n502 = ( x73 & x74 ) | ( x73 & ~x75 ) | ( x74 & ~x75 ) ;
  assign n503 = ( x74 & n386 ) | ( x74 & n494 ) | ( n386 & n494 ) ;
  assign n504 = ~n502 & n503 ;
  assign n505 = ~n370 & n492 ;
  assign n506 = ( n497 & ~n498 ) | ( n497 & n505 ) | ( ~n498 & n505 ) ;
  assign n507 = n501 | n506 ;
  assign n508 = ( n501 & ~n504 ) | ( n501 & n507 ) | ( ~n504 & n507 ) ;
  assign n509 = x0 & n508 ;
  assign n510 = ( x1 & x2 ) | ( x1 & n509 ) | ( x2 & n509 ) ;
  assign n511 = x74 & n172 ;
  assign n512 = x75 | n511 ;
  assign n513 = ( n147 & n511 ) | ( n147 & n512 ) | ( n511 & n512 ) ;
  assign n514 = ( ~x73 & n135 ) | ( ~x73 & n174 ) | ( n135 & n174 ) ;
  assign n515 = n513 | n514 ;
  assign n516 = n510 | n515 ;
  assign n517 = n510 & n515 ;
  assign n518 = n516 & ~n517 ;
  assign n519 = n206 & n372 ;
  assign n520 = x5 & n519 ;
  assign n521 = x72 & n205 ;
  assign n522 = x71 & n201 ;
  assign n523 = n521 | n522 ;
  assign n524 = x70 & n221 ;
  assign n525 = n523 | n524 ;
  assign n526 = ( ~x5 & n519 ) | ( ~x5 & n525 ) | ( n519 & n525 ) ;
  assign n527 = x5 & ~n525 ;
  assign n528 = ( ~n520 & n526 ) | ( ~n520 & n527 ) | ( n526 & n527 ) ;
  assign n529 = x65 & n453 ;
  assign n530 = n226 & n449 ;
  assign n531 = n529 | n530 ;
  assign n532 = x66 & n456 ;
  assign n533 = n531 | n532 ;
  assign n534 = n410 & n448 ;
  assign n535 = ~n409 & n447 ;
  assign n536 = n534 | n535 ;
  assign n537 = x64 & n536 ;
  assign n538 = n533 | n537 ;
  assign n539 = ~x11 & n538 ;
  assign n540 = ( x11 & n459 ) | ( x11 & n538 ) | ( n459 & n538 ) ;
  assign n541 = n459 & n538 ;
  assign n542 = ( n539 & n540 ) | ( n539 & ~n541 ) | ( n540 & ~n541 ) ;
  assign n543 = n240 & n301 ;
  assign n544 = x8 & n543 ;
  assign n545 = x69 & n309 ;
  assign n546 = x68 & n306 ;
  assign n547 = n545 | n546 ;
  assign n548 = x67 & n359 ;
  assign n549 = n547 | n548 ;
  assign n550 = ( ~x8 & n543 ) | ( ~x8 & n549 ) | ( n543 & n549 ) ;
  assign n551 = x8 & ~n549 ;
  assign n552 = ( ~n544 & n550 ) | ( ~n544 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( n474 & n542 ) | ( n474 & n552 ) | ( n542 & n552 ) ;
  assign n554 = ( ~n474 & n542 ) | ( ~n474 & n552 ) | ( n542 & n552 ) ;
  assign n555 = ( n474 & ~n553 ) | ( n474 & n554 ) | ( ~n553 & n554 ) ;
  assign n556 = ( n487 & ~n528 ) | ( n487 & n555 ) | ( ~n528 & n555 ) ;
  assign n557 = ( n487 & n528 ) | ( n487 & n555 ) | ( n528 & n555 ) ;
  assign n558 = ( n528 & n556 ) | ( n528 & ~n557 ) | ( n556 & ~n557 ) ;
  assign n559 = ( n490 & n518 ) | ( n490 & n558 ) | ( n518 & n558 ) ;
  assign n560 = ( ~n490 & n518 ) | ( ~n490 & n558 ) | ( n518 & n558 ) ;
  assign n561 = ( n490 & ~n559 ) | ( n490 & n560 ) | ( ~n559 & n560 ) ;
  assign n562 = ( x75 & n503 ) | ( x75 & ~n507 ) | ( n503 & ~n507 ) ;
  assign n563 = ( x75 & x76 ) | ( x75 & n562 ) | ( x76 & n562 ) ;
  assign n564 = ( ~x75 & x76 ) | ( ~x75 & n562 ) | ( x76 & n562 ) ;
  assign n565 = ( x75 & ~n563 ) | ( x75 & n564 ) | ( ~n563 & n564 ) ;
  assign n566 = x0 & n565 ;
  assign n567 = ( x1 & x2 ) | ( x1 & n566 ) | ( x2 & n566 ) ;
  assign n568 = x76 & n147 ;
  assign n569 = x75 & n172 ;
  assign n570 = n174 | n569 ;
  assign n571 = ~x74 & n136 ;
  assign n572 = n570 | n571 ;
  assign n573 = n568 | n572 ;
  assign n574 = n567 | n573 ;
  assign n575 = n567 & n573 ;
  assign n576 = n574 & ~n575 ;
  assign n577 = n276 & n301 ;
  assign n578 = x8 & n577 ;
  assign n579 = x70 & n309 ;
  assign n580 = x69 & n306 ;
  assign n581 = n579 | n580 ;
  assign n582 = x68 & n359 ;
  assign n583 = n581 | n582 ;
  assign n584 = ( ~x8 & n577 ) | ( ~x8 & n583 ) | ( n577 & n583 ) ;
  assign n585 = x8 & ~n583 ;
  assign n586 = ( ~n578 & n584 ) | ( ~n578 & n585 ) | ( n584 & n585 ) ;
  assign n587 = n459 | n538 ;
  assign n588 = x11 & n587 ;
  assign n589 = x66 & n453 ;
  assign n590 = n169 & n449 ;
  assign n591 = x67 & n456 ;
  assign n592 = x65 & ~n536 ;
  assign n593 = ( x65 & n591 ) | ( x65 & ~n592 ) | ( n591 & ~n592 ) ;
  assign n594 = n590 | n593 ;
  assign n595 = n589 | n594 ;
  assign n596 = x11 | x12 ;
  assign n597 = x11 & x12 ;
  assign n598 = n596 & ~n597 ;
  assign n599 = x64 & n598 ;
  assign n600 = ( n588 & ~n595 ) | ( n588 & n599 ) | ( ~n595 & n599 ) ;
  assign n601 = x11 & ~n595 ;
  assign n602 = ( ~n588 & n595 ) | ( ~n588 & n601 ) | ( n595 & n601 ) ;
  assign n603 = ( n599 & n601 ) | ( n599 & n602 ) | ( n601 & n602 ) ;
  assign n604 = ( n600 & n602 ) | ( n600 & ~n603 ) | ( n602 & ~n603 ) ;
  assign n605 = ( n553 & n586 ) | ( n553 & n604 ) | ( n586 & n604 ) ;
  assign n606 = ( ~n553 & n586 ) | ( ~n553 & n604 ) | ( n586 & n604 ) ;
  assign n607 = ( n553 & ~n605 ) | ( n553 & n606 ) | ( ~n605 & n606 ) ;
  assign n608 = n206 & n388 ;
  assign n609 = x5 & n608 ;
  assign n610 = x73 & n205 ;
  assign n611 = x72 & n201 ;
  assign n612 = n610 | n611 ;
  assign n613 = x71 & n221 ;
  assign n614 = n612 | n613 ;
  assign n615 = ( ~x5 & n608 ) | ( ~x5 & n614 ) | ( n608 & n614 ) ;
  assign n616 = x5 & ~n614 ;
  assign n617 = ( ~n609 & n615 ) | ( ~n609 & n616 ) | ( n615 & n616 ) ;
  assign n618 = ( n557 & ~n607 ) | ( n557 & n617 ) | ( ~n607 & n617 ) ;
  assign n619 = ( n557 & n607 ) | ( n557 & n617 ) | ( n607 & n617 ) ;
  assign n620 = ( n607 & n618 ) | ( n607 & ~n619 ) | ( n618 & ~n619 ) ;
  assign n621 = ( n559 & n576 ) | ( n559 & n620 ) | ( n576 & n620 ) ;
  assign n622 = ( ~n559 & n576 ) | ( ~n559 & n620 ) | ( n576 & n620 ) ;
  assign n623 = ( n559 & ~n621 ) | ( n559 & n622 ) | ( ~n621 & n622 ) ;
  assign n624 = ( x76 & x77 ) | ( x76 & n563 ) | ( x77 & n563 ) ;
  assign n625 = ( x76 & x77 ) | ( x76 & ~n563 ) | ( x77 & ~n563 ) ;
  assign n626 = ( n563 & ~n624 ) | ( n563 & n625 ) | ( ~n624 & n625 ) ;
  assign n627 = x0 & n626 ;
  assign n628 = ( x1 & x2 ) | ( x1 & n627 ) | ( x2 & n627 ) ;
  assign n629 = x76 & n172 ;
  assign n630 = ( ~x75 & n135 ) | ( ~x75 & n174 ) | ( n135 & n174 ) ;
  assign n631 = n629 | n630 ;
  assign n632 = x77 & n147 ;
  assign n633 = n631 | n632 ;
  assign n634 = n628 | n633 ;
  assign n635 = n628 & n633 ;
  assign n636 = n634 & ~n635 ;
  assign n637 = x67 & n453 ;
  assign n638 = x11 & n637 ;
  assign n639 = x68 & n456 ;
  assign n640 = x66 & n536 ;
  assign n641 = n639 | n640 ;
  assign n642 = n193 & n449 ;
  assign n643 = n641 | n642 ;
  assign n644 = ( ~x11 & n637 ) | ( ~x11 & n643 ) | ( n637 & n643 ) ;
  assign n645 = x11 & ~n643 ;
  assign n646 = ( ~n638 & n644 ) | ( ~n638 & n645 ) | ( n644 & n645 ) ;
  assign n647 = ~x13 & x14 ;
  assign n648 = x13 & ~x14 ;
  assign n649 = ( n598 & n647 ) | ( n598 & n648 ) | ( n647 & n648 ) ;
  assign n650 = n302 & n649 ;
  assign n651 = ~x11 & x13 ;
  assign n652 = x12 & x13 ;
  assign n653 = ( n597 & n651 ) | ( n597 & ~n652 ) | ( n651 & ~n652 ) ;
  assign n654 = x64 & n653 ;
  assign n655 = n650 | n654 ;
  assign n656 = n598 & ~n649 ;
  assign n657 = x65 & n656 ;
  assign n658 = n655 | n657 ;
  assign n659 = n599 | n658 ;
  assign n660 = ( x14 & n599 ) | ( x14 & ~n658 ) | ( n599 & ~n658 ) ;
  assign n661 = x14 & ~n658 ;
  assign n662 = ( n659 & ~n660 ) | ( n659 & n661 ) | ( ~n660 & n661 ) ;
  assign n663 = ( ~n603 & n646 ) | ( ~n603 & n662 ) | ( n646 & n662 ) ;
  assign n664 = ( n603 & n646 ) | ( n603 & n662 ) | ( n646 & n662 ) ;
  assign n665 = ( n603 & n663 ) | ( n603 & ~n664 ) | ( n663 & ~n664 ) ;
  assign n666 = n301 & n322 ;
  assign n667 = x8 & n666 ;
  assign n668 = x71 & n309 ;
  assign n669 = x70 & n306 ;
  assign n670 = n668 | n669 ;
  assign n671 = x69 & n359 ;
  assign n672 = n670 | n671 ;
  assign n673 = ( ~x8 & n666 ) | ( ~x8 & n672 ) | ( n666 & n672 ) ;
  assign n674 = x8 & ~n672 ;
  assign n675 = ( ~n667 & n673 ) | ( ~n667 & n674 ) | ( n673 & n674 ) ;
  assign n676 = ( n605 & ~n665 ) | ( n605 & n675 ) | ( ~n665 & n675 ) ;
  assign n677 = ( n605 & n665 ) | ( n605 & n675 ) | ( n665 & n675 ) ;
  assign n678 = ( n665 & n676 ) | ( n665 & ~n677 ) | ( n676 & ~n677 ) ;
  assign n679 = n206 & n436 ;
  assign n680 = x5 & n679 ;
  assign n681 = x74 & n205 ;
  assign n682 = x73 & n201 ;
  assign n683 = n681 | n682 ;
  assign n684 = x72 & n221 ;
  assign n685 = n683 | n684 ;
  assign n686 = ( ~x5 & n679 ) | ( ~x5 & n685 ) | ( n679 & n685 ) ;
  assign n687 = x5 & ~n685 ;
  assign n688 = ( ~n680 & n686 ) | ( ~n680 & n687 ) | ( n686 & n687 ) ;
  assign n689 = ( n619 & ~n678 ) | ( n619 & n688 ) | ( ~n678 & n688 ) ;
  assign n690 = ( n619 & n678 ) | ( n619 & n688 ) | ( n678 & n688 ) ;
  assign n691 = ( n678 & n689 ) | ( n678 & ~n690 ) | ( n689 & ~n690 ) ;
  assign n692 = ( ~n621 & n636 ) | ( ~n621 & n691 ) | ( n636 & n691 ) ;
  assign n693 = ( n621 & n636 ) | ( n621 & n691 ) | ( n636 & n691 ) ;
  assign n694 = ( n621 & n692 ) | ( n621 & ~n693 ) | ( n692 & ~n693 ) ;
  assign n695 = ( x76 & x78 ) | ( x76 & ~n625 ) | ( x78 & ~n625 ) ;
  assign n696 = ( x77 & x78 ) | ( x77 & n624 ) | ( x78 & n624 ) ;
  assign n697 = ( x77 & n695 ) | ( x77 & ~n696 ) | ( n695 & ~n696 ) ;
  assign n698 = x0 & n697 ;
  assign n699 = ( x1 & x2 ) | ( x1 & n698 ) | ( x2 & n698 ) ;
  assign n700 = x77 & n172 ;
  assign n701 = x78 | n700 ;
  assign n702 = ( n147 & n700 ) | ( n147 & n701 ) | ( n700 & n701 ) ;
  assign n703 = ( ~x76 & n135 ) | ( ~x76 & n174 ) | ( n135 & n174 ) ;
  assign n704 = n702 | n703 ;
  assign n705 = n699 | n704 ;
  assign n706 = n699 & n704 ;
  assign n707 = n705 & ~n706 ;
  assign n708 = n206 & n508 ;
  assign n709 = x5 & n708 ;
  assign n710 = x75 & n205 ;
  assign n711 = x74 & n201 ;
  assign n712 = n710 | n711 ;
  assign n713 = x73 & n221 ;
  assign n714 = n712 | n713 ;
  assign n715 = ( ~x5 & n708 ) | ( ~x5 & n714 ) | ( n708 & n714 ) ;
  assign n716 = x5 & ~n714 ;
  assign n717 = ( ~n709 & n715 ) | ( ~n709 & n716 ) | ( n715 & n716 ) ;
  assign n718 = n301 & n372 ;
  assign n719 = x8 & n718 ;
  assign n720 = x72 & n309 ;
  assign n721 = x71 & n306 ;
  assign n722 = n720 | n721 ;
  assign n723 = x70 & n359 ;
  assign n724 = n722 | n723 ;
  assign n725 = ( ~x8 & n718 ) | ( ~x8 & n724 ) | ( n718 & n724 ) ;
  assign n726 = x8 & ~n724 ;
  assign n727 = ( ~n719 & n725 ) | ( ~n719 & n726 ) | ( n725 & n726 ) ;
  assign n728 = n240 & n449 ;
  assign n729 = x11 & n728 ;
  assign n730 = x69 & n456 ;
  assign n731 = x68 & n453 ;
  assign n732 = n730 | n731 ;
  assign n733 = x67 & n536 ;
  assign n734 = n732 | n733 ;
  assign n735 = ( ~x11 & n728 ) | ( ~x11 & n734 ) | ( n728 & n734 ) ;
  assign n736 = x11 & ~n734 ;
  assign n737 = ( ~n729 & n735 ) | ( ~n729 & n736 ) | ( n735 & n736 ) ;
  assign n738 = x66 & n656 ;
  assign n739 = n226 & n649 ;
  assign n740 = n738 | n739 ;
  assign n741 = x65 & n653 ;
  assign n742 = n597 & n648 ;
  assign n743 = ~n596 & n647 ;
  assign n744 = n742 | n743 ;
  assign n745 = x64 & ~n744 ;
  assign n746 = ( x64 & n741 ) | ( x64 & ~n745 ) | ( n741 & ~n745 ) ;
  assign n747 = n740 | n746 ;
  assign n748 = ~x14 & n747 ;
  assign n749 = ( x14 & n659 ) | ( x14 & n747 ) | ( n659 & n747 ) ;
  assign n750 = n659 & n747 ;
  assign n751 = ( n748 & n749 ) | ( n748 & ~n750 ) | ( n749 & ~n750 ) ;
  assign n752 = ( n664 & ~n737 ) | ( n664 & n751 ) | ( ~n737 & n751 ) ;
  assign n753 = ( n664 & n737 ) | ( n664 & n751 ) | ( n737 & n751 ) ;
  assign n754 = ( n737 & n752 ) | ( n737 & ~n753 ) | ( n752 & ~n753 ) ;
  assign n755 = ( ~n677 & n727 ) | ( ~n677 & n754 ) | ( n727 & n754 ) ;
  assign n756 = ( n677 & n727 ) | ( n677 & n754 ) | ( n727 & n754 ) ;
  assign n757 = ( n677 & n755 ) | ( n677 & ~n756 ) | ( n755 & ~n756 ) ;
  assign n758 = ( n690 & ~n717 ) | ( n690 & n757 ) | ( ~n717 & n757 ) ;
  assign n759 = ( n690 & n717 ) | ( n690 & n757 ) | ( n717 & n757 ) ;
  assign n760 = ( n717 & n758 ) | ( n717 & ~n759 ) | ( n758 & ~n759 ) ;
  assign n761 = ( n693 & n707 ) | ( n693 & n760 ) | ( n707 & n760 ) ;
  assign n762 = ( ~n693 & n707 ) | ( ~n693 & n760 ) | ( n707 & n760 ) ;
  assign n763 = ( n693 & ~n761 ) | ( n693 & n762 ) | ( ~n761 & n762 ) ;
  assign n764 = n206 & n565 ;
  assign n765 = x5 & n764 ;
  assign n766 = x76 & n205 ;
  assign n767 = x75 & n201 ;
  assign n768 = n766 | n767 ;
  assign n769 = x74 & n221 ;
  assign n770 = n768 | n769 ;
  assign n771 = ( ~x5 & n764 ) | ( ~x5 & n770 ) | ( n764 & n770 ) ;
  assign n772 = x5 & ~n770 ;
  assign n773 = ( ~n765 & n771 ) | ( ~n765 & n772 ) | ( n771 & n772 ) ;
  assign n774 = n276 & n449 ;
  assign n775 = x11 & n774 ;
  assign n776 = x70 & n456 ;
  assign n777 = x69 & n453 ;
  assign n778 = n776 | n777 ;
  assign n779 = x68 & n536 ;
  assign n780 = n778 | n779 ;
  assign n781 = ( ~x11 & n774 ) | ( ~x11 & n780 ) | ( n774 & n780 ) ;
  assign n782 = x11 & ~n780 ;
  assign n783 = ( ~n775 & n781 ) | ( ~n775 & n782 ) | ( n781 & n782 ) ;
  assign n784 = x14 & n747 ;
  assign n785 = ( x14 & n659 ) | ( x14 & n784 ) | ( n659 & n784 ) ;
  assign n786 = x66 & n653 ;
  assign n787 = n169 & n649 ;
  assign n788 = x67 & n656 ;
  assign n789 = x65 & ~n744 ;
  assign n790 = ( x65 & n788 ) | ( x65 & ~n789 ) | ( n788 & ~n789 ) ;
  assign n791 = n787 | n790 ;
  assign n792 = n786 | n791 ;
  assign n793 = x14 & x15 ;
  assign n794 = x14 | x15 ;
  assign n795 = ~n793 & n794 ;
  assign n796 = x64 & n795 ;
  assign n797 = ( n785 & ~n792 ) | ( n785 & n796 ) | ( ~n792 & n796 ) ;
  assign n798 = x14 & ~n792 ;
  assign n799 = ( ~n785 & n792 ) | ( ~n785 & n798 ) | ( n792 & n798 ) ;
  assign n800 = ( n796 & n798 ) | ( n796 & n799 ) | ( n798 & n799 ) ;
  assign n801 = ( n797 & n799 ) | ( n797 & ~n800 ) | ( n799 & ~n800 ) ;
  assign n802 = ( n753 & n783 ) | ( n753 & n801 ) | ( n783 & n801 ) ;
  assign n803 = ( ~n753 & n783 ) | ( ~n753 & n801 ) | ( n783 & n801 ) ;
  assign n804 = ( n753 & ~n802 ) | ( n753 & n803 ) | ( ~n802 & n803 ) ;
  assign n805 = n301 & n388 ;
  assign n806 = x8 & n805 ;
  assign n807 = x73 & n309 ;
  assign n808 = x72 & n306 ;
  assign n809 = n807 | n808 ;
  assign n810 = x71 & n359 ;
  assign n811 = n809 | n810 ;
  assign n812 = ( ~x8 & n805 ) | ( ~x8 & n811 ) | ( n805 & n811 ) ;
  assign n813 = x8 & ~n811 ;
  assign n814 = ( ~n806 & n812 ) | ( ~n806 & n813 ) | ( n812 & n813 ) ;
  assign n815 = ( n756 & ~n804 ) | ( n756 & n814 ) | ( ~n804 & n814 ) ;
  assign n816 = ( n756 & n804 ) | ( n756 & n814 ) | ( n804 & n814 ) ;
  assign n817 = ( n804 & n815 ) | ( n804 & ~n816 ) | ( n815 & ~n816 ) ;
  assign n818 = ( n759 & n773 ) | ( n759 & n817 ) | ( n773 & n817 ) ;
  assign n819 = ( ~n759 & n773 ) | ( ~n759 & n817 ) | ( n773 & n817 ) ;
  assign n820 = ( n759 & ~n818 ) | ( n759 & n819 ) | ( ~n818 & n819 ) ;
  assign n821 = ( ~x78 & x79 ) | ( ~x78 & n696 ) | ( x79 & n696 ) ;
  assign n822 = ( x78 & x79 ) | ( x78 & n696 ) | ( x79 & n696 ) ;
  assign n823 = ( x78 & n821 ) | ( x78 & ~n822 ) | ( n821 & ~n822 ) ;
  assign n824 = x0 & n823 ;
  assign n825 = ( x1 & x2 ) | ( x1 & n824 ) | ( x2 & n824 ) ;
  assign n826 = x79 & n147 ;
  assign n827 = ~x77 & n136 ;
  assign n828 = x78 & n172 ;
  assign n829 = n174 | n828 ;
  assign n830 = n827 | n829 ;
  assign n831 = n826 | n830 ;
  assign n832 = n825 | n831 ;
  assign n833 = n825 & n831 ;
  assign n834 = n832 & ~n833 ;
  assign n835 = ( n761 & ~n820 ) | ( n761 & n834 ) | ( ~n820 & n834 ) ;
  assign n836 = ( n761 & n820 ) | ( n761 & n834 ) | ( n820 & n834 ) ;
  assign n837 = ( n820 & n835 ) | ( n820 & ~n836 ) | ( n835 & ~n836 ) ;
  assign n838 = ( x79 & x80 ) | ( x79 & n822 ) | ( x80 & n822 ) ;
  assign n839 = ( x79 & x80 ) | ( x79 & ~n822 ) | ( x80 & ~n822 ) ;
  assign n840 = ( n822 & ~n838 ) | ( n822 & n839 ) | ( ~n838 & n839 ) ;
  assign n841 = x0 & n840 ;
  assign n842 = ( x1 & x2 ) | ( x1 & n841 ) | ( x2 & n841 ) ;
  assign n843 = x79 & n172 ;
  assign n844 = ( ~x78 & n135 ) | ( ~x78 & n174 ) | ( n135 & n174 ) ;
  assign n845 = n843 | n844 ;
  assign n846 = x80 & n147 ;
  assign n847 = n845 | n846 ;
  assign n848 = n842 | n847 ;
  assign n849 = n842 & n847 ;
  assign n850 = n848 & ~n849 ;
  assign n851 = n322 & n449 ;
  assign n852 = x11 & n851 ;
  assign n853 = x71 & n456 ;
  assign n854 = x70 & n453 ;
  assign n855 = n853 | n854 ;
  assign n856 = x69 & n536 ;
  assign n857 = n855 | n856 ;
  assign n858 = ( ~x11 & n851 ) | ( ~x11 & n857 ) | ( n851 & n857 ) ;
  assign n859 = x11 & ~n857 ;
  assign n860 = ( ~n852 & n858 ) | ( ~n852 & n859 ) | ( n858 & n859 ) ;
  assign n861 = x68 & n656 ;
  assign n862 = x14 & n861 ;
  assign n863 = x67 & n653 ;
  assign n864 = x66 & n744 ;
  assign n865 = n863 | n864 ;
  assign n866 = n193 & n649 ;
  assign n867 = n865 | n866 ;
  assign n868 = ( ~x14 & n861 ) | ( ~x14 & n867 ) | ( n861 & n867 ) ;
  assign n869 = x14 & ~n867 ;
  assign n870 = ( ~n862 & n868 ) | ( ~n862 & n869 ) | ( n868 & n869 ) ;
  assign n871 = x16 & x17 ;
  assign n872 = x16 | x17 ;
  assign n873 = ~n871 & n872 ;
  assign n874 = n795 & n873 ;
  assign n875 = n302 & n874 ;
  assign n876 = ~x14 & x16 ;
  assign n877 = x15 & x16 ;
  assign n878 = ( n793 & n876 ) | ( n793 & ~n877 ) | ( n876 & ~n877 ) ;
  assign n879 = x64 & n878 ;
  assign n880 = n875 | n879 ;
  assign n881 = ( n795 & n871 ) | ( n795 & ~n872 ) | ( n871 & ~n872 ) ;
  assign n882 = x65 & n881 ;
  assign n883 = n880 | n882 ;
  assign n884 = n796 | n883 ;
  assign n885 = ( x17 & n796 ) | ( x17 & ~n883 ) | ( n796 & ~n883 ) ;
  assign n886 = x17 & ~n883 ;
  assign n887 = ( n884 & ~n885 ) | ( n884 & n886 ) | ( ~n885 & n886 ) ;
  assign n888 = ( n800 & ~n870 ) | ( n800 & n887 ) | ( ~n870 & n887 ) ;
  assign n889 = ( n800 & n870 ) | ( n800 & n887 ) | ( n870 & n887 ) ;
  assign n890 = ( n870 & n888 ) | ( n870 & ~n889 ) | ( n888 & ~n889 ) ;
  assign n891 = ( n802 & n860 ) | ( n802 & n890 ) | ( n860 & n890 ) ;
  assign n892 = ( ~n802 & n860 ) | ( ~n802 & n890 ) | ( n860 & n890 ) ;
  assign n893 = ( n802 & ~n891 ) | ( n802 & n892 ) | ( ~n891 & n892 ) ;
  assign n894 = n301 & n436 ;
  assign n895 = x8 & n894 ;
  assign n896 = x74 & n309 ;
  assign n897 = x73 & n306 ;
  assign n898 = n896 | n897 ;
  assign n899 = x72 & n359 ;
  assign n900 = n898 | n899 ;
  assign n901 = ( ~x8 & n894 ) | ( ~x8 & n900 ) | ( n894 & n900 ) ;
  assign n902 = x8 & ~n900 ;
  assign n903 = ( ~n895 & n901 ) | ( ~n895 & n902 ) | ( n901 & n902 ) ;
  assign n904 = ( n816 & ~n893 ) | ( n816 & n903 ) | ( ~n893 & n903 ) ;
  assign n905 = ( n816 & n893 ) | ( n816 & n903 ) | ( n893 & n903 ) ;
  assign n906 = ( n893 & n904 ) | ( n893 & ~n905 ) | ( n904 & ~n905 ) ;
  assign n907 = n206 & n626 ;
  assign n908 = x5 & n907 ;
  assign n909 = x77 & n205 ;
  assign n910 = x76 & n201 ;
  assign n911 = n909 | n910 ;
  assign n912 = x75 & n221 ;
  assign n913 = n911 | n912 ;
  assign n914 = ( ~x5 & n907 ) | ( ~x5 & n913 ) | ( n907 & n913 ) ;
  assign n915 = x5 & ~n913 ;
  assign n916 = ( ~n908 & n914 ) | ( ~n908 & n915 ) | ( n914 & n915 ) ;
  assign n917 = ( n818 & ~n906 ) | ( n818 & n916 ) | ( ~n906 & n916 ) ;
  assign n918 = ( n818 & n906 ) | ( n818 & n916 ) | ( n906 & n916 ) ;
  assign n919 = ( n906 & n917 ) | ( n906 & ~n918 ) | ( n917 & ~n918 ) ;
  assign n920 = ( n836 & n850 ) | ( n836 & n919 ) | ( n850 & n919 ) ;
  assign n921 = ( ~n836 & n850 ) | ( ~n836 & n919 ) | ( n850 & n919 ) ;
  assign n922 = ( n836 & ~n920 ) | ( n836 & n921 ) | ( ~n920 & n921 ) ;
  assign n923 = n206 & n697 ;
  assign n924 = x5 & n923 ;
  assign n925 = x78 & n205 ;
  assign n926 = x77 & n201 ;
  assign n927 = n925 | n926 ;
  assign n928 = x76 & n221 ;
  assign n929 = n927 | n928 ;
  assign n930 = ( ~x5 & n923 ) | ( ~x5 & n929 ) | ( n923 & n929 ) ;
  assign n931 = x5 & ~n929 ;
  assign n932 = ( ~n924 & n930 ) | ( ~n924 & n931 ) | ( n930 & n931 ) ;
  assign n933 = n301 & n508 ;
  assign n934 = x8 & n933 ;
  assign n935 = x75 & n309 ;
  assign n936 = x74 & n306 ;
  assign n937 = n935 | n936 ;
  assign n938 = x73 & n359 ;
  assign n939 = n937 | n938 ;
  assign n940 = ( ~x8 & n933 ) | ( ~x8 & n939 ) | ( n933 & n939 ) ;
  assign n941 = x8 & ~n939 ;
  assign n942 = ( ~n934 & n940 ) | ( ~n934 & n941 ) | ( n940 & n941 ) ;
  assign n943 = n372 & n449 ;
  assign n944 = x11 & n943 ;
  assign n945 = x72 & n456 ;
  assign n946 = x71 & n453 ;
  assign n947 = n945 | n946 ;
  assign n948 = x70 & n536 ;
  assign n949 = n947 | n948 ;
  assign n950 = ( ~x11 & n943 ) | ( ~x11 & n949 ) | ( n943 & n949 ) ;
  assign n951 = x11 & ~n949 ;
  assign n952 = ( ~n944 & n950 ) | ( ~n944 & n951 ) | ( n950 & n951 ) ;
  assign n953 = x65 & n878 ;
  assign n954 = n226 & n874 ;
  assign n955 = n953 | n954 ;
  assign n956 = x66 & n881 ;
  assign n957 = n955 | n956 ;
  assign n958 = ~n795 & n873 ;
  assign n959 = ~n878 & n958 ;
  assign n960 = x64 & n959 ;
  assign n961 = n957 | n960 ;
  assign n962 = ~x17 & n961 ;
  assign n963 = ( x17 & n884 ) | ( x17 & n961 ) | ( n884 & n961 ) ;
  assign n964 = n884 & n961 ;
  assign n965 = ( n962 & n963 ) | ( n962 & ~n964 ) | ( n963 & ~n964 ) ;
  assign n966 = n240 & n649 ;
  assign n967 = x14 & n966 ;
  assign n968 = x69 & n656 ;
  assign n969 = x68 & n653 ;
  assign n970 = n968 | n969 ;
  assign n971 = x67 & n744 ;
  assign n972 = n970 | n971 ;
  assign n973 = ( ~x14 & n966 ) | ( ~x14 & n972 ) | ( n966 & n972 ) ;
  assign n974 = x14 & ~n972 ;
  assign n975 = ( ~n967 & n973 ) | ( ~n967 & n974 ) | ( n973 & n974 ) ;
  assign n976 = ( n889 & n965 ) | ( n889 & n975 ) | ( n965 & n975 ) ;
  assign n977 = ( ~n889 & n965 ) | ( ~n889 & n975 ) | ( n965 & n975 ) ;
  assign n978 = ( n889 & ~n976 ) | ( n889 & n977 ) | ( ~n976 & n977 ) ;
  assign n979 = ( n891 & ~n952 ) | ( n891 & n978 ) | ( ~n952 & n978 ) ;
  assign n980 = ( n891 & n952 ) | ( n891 & n978 ) | ( n952 & n978 ) ;
  assign n981 = ( n952 & n979 ) | ( n952 & ~n980 ) | ( n979 & ~n980 ) ;
  assign n982 = ( n905 & n942 ) | ( n905 & n981 ) | ( n942 & n981 ) ;
  assign n983 = ( ~n905 & n942 ) | ( ~n905 & n981 ) | ( n942 & n981 ) ;
  assign n984 = ( n905 & ~n982 ) | ( n905 & n983 ) | ( ~n982 & n983 ) ;
  assign n985 = ( n918 & n932 ) | ( n918 & n984 ) | ( n932 & n984 ) ;
  assign n986 = ( ~n918 & n932 ) | ( ~n918 & n984 ) | ( n932 & n984 ) ;
  assign n987 = ( n918 & ~n985 ) | ( n918 & n986 ) | ( ~n985 & n986 ) ;
  assign n988 = ( x80 & x81 ) | ( x80 & n838 ) | ( x81 & n838 ) ;
  assign n989 = ( x79 & x81 ) | ( x79 & ~n839 ) | ( x81 & ~n839 ) ;
  assign n990 = ( x80 & ~n988 ) | ( x80 & n989 ) | ( ~n988 & n989 ) ;
  assign n991 = x0 & n990 ;
  assign n992 = ( x1 & x2 ) | ( x1 & n991 ) | ( x2 & n991 ) ;
  assign n993 = x80 & n172 ;
  assign n994 = x81 | n993 ;
  assign n995 = ( n147 & n993 ) | ( n147 & n994 ) | ( n993 & n994 ) ;
  assign n996 = ( ~x79 & n135 ) | ( ~x79 & n174 ) | ( n135 & n174 ) ;
  assign n997 = n995 | n996 ;
  assign n998 = n992 | n997 ;
  assign n999 = n992 & n997 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ( n920 & ~n987 ) | ( n920 & n1000 ) | ( ~n987 & n1000 ) ;
  assign n1002 = ( n920 & n987 ) | ( n920 & n1000 ) | ( n987 & n1000 ) ;
  assign n1003 = ( n987 & n1001 ) | ( n987 & ~n1002 ) | ( n1001 & ~n1002 ) ;
  assign n1004 = ( ~x81 & x82 ) | ( ~x81 & n988 ) | ( x82 & n988 ) ;
  assign n1005 = ( x81 & x82 ) | ( x81 & n988 ) | ( x82 & n988 ) ;
  assign n1006 = ( x81 & n1004 ) | ( x81 & ~n1005 ) | ( n1004 & ~n1005 ) ;
  assign n1007 = x0 & n1006 ;
  assign n1008 = ( x1 & x2 ) | ( x1 & n1007 ) | ( x2 & n1007 ) ;
  assign n1009 = x82 & n147 ;
  assign n1010 = x81 & n172 ;
  assign n1011 = n174 | n1010 ;
  assign n1012 = ~x80 & n136 ;
  assign n1013 = n1011 | n1012 ;
  assign n1014 = n1009 | n1013 ;
  assign n1015 = n1008 | n1014 ;
  assign n1016 = n1008 & n1014 ;
  assign n1017 = n1015 & ~n1016 ;
  assign n1018 = n206 & n823 ;
  assign n1019 = x5 & n1018 ;
  assign n1020 = x79 & n205 ;
  assign n1021 = x78 & n201 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = x77 & n221 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = ( ~x5 & n1018 ) | ( ~x5 & n1024 ) | ( n1018 & n1024 ) ;
  assign n1026 = x5 & ~n1024 ;
  assign n1027 = ( ~n1019 & n1025 ) | ( ~n1019 & n1026 ) | ( n1025 & n1026 ) ;
  assign n1028 = n301 & n565 ;
  assign n1029 = x8 & n1028 ;
  assign n1030 = x76 & n309 ;
  assign n1031 = x75 & n306 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = x74 & n359 ;
  assign n1034 = n1032 | n1033 ;
  assign n1035 = ( ~x8 & n1028 ) | ( ~x8 & n1034 ) | ( n1028 & n1034 ) ;
  assign n1036 = x8 & ~n1034 ;
  assign n1037 = ( ~n1029 & n1035 ) | ( ~n1029 & n1036 ) | ( n1035 & n1036 ) ;
  assign n1038 = n388 & n449 ;
  assign n1039 = x11 & n1038 ;
  assign n1040 = x73 & n456 ;
  assign n1041 = x72 & n453 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = x71 & n536 ;
  assign n1044 = n1042 | n1043 ;
  assign n1045 = ( ~x11 & n1038 ) | ( ~x11 & n1044 ) | ( n1038 & n1044 ) ;
  assign n1046 = x11 & ~n1044 ;
  assign n1047 = ( ~n1039 & n1045 ) | ( ~n1039 & n1046 ) | ( n1045 & n1046 ) ;
  assign n1048 = n276 & n649 ;
  assign n1049 = x14 & n1048 ;
  assign n1050 = x70 & n656 ;
  assign n1051 = x69 & n653 ;
  assign n1052 = n1050 | n1051 ;
  assign n1053 = x68 & n744 ;
  assign n1054 = n1052 | n1053 ;
  assign n1055 = ( ~x14 & n1048 ) | ( ~x14 & n1054 ) | ( n1048 & n1054 ) ;
  assign n1056 = x14 & ~n1054 ;
  assign n1057 = ( ~n1049 & n1055 ) | ( ~n1049 & n1056 ) | ( n1055 & n1056 ) ;
  assign n1058 = n884 | n961 ;
  assign n1059 = x17 & n1058 ;
  assign n1060 = x67 & n881 ;
  assign n1061 = x66 & n878 ;
  assign n1062 = n1060 | n1061 ;
  assign n1063 = x65 & n959 ;
  assign n1064 = n1062 | n1063 ;
  assign n1065 = n169 & n874 ;
  assign n1066 = n1064 | n1065 ;
  assign n1067 = x17 | x18 ;
  assign n1068 = x17 & x18 ;
  assign n1069 = n1067 & ~n1068 ;
  assign n1070 = x64 & n1069 ;
  assign n1071 = ( n1059 & ~n1066 ) | ( n1059 & n1070 ) | ( ~n1066 & n1070 ) ;
  assign n1072 = x17 & ~n1066 ;
  assign n1073 = ( ~n1059 & n1066 ) | ( ~n1059 & n1072 ) | ( n1066 & n1072 ) ;
  assign n1074 = ( n1070 & n1072 ) | ( n1070 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1075 = ( n1071 & n1073 ) | ( n1071 & ~n1074 ) | ( n1073 & ~n1074 ) ;
  assign n1076 = ( n976 & n1057 ) | ( n976 & n1075 ) | ( n1057 & n1075 ) ;
  assign n1077 = ( ~n976 & n1057 ) | ( ~n976 & n1075 ) | ( n1057 & n1075 ) ;
  assign n1078 = ( n976 & ~n1076 ) | ( n976 & n1077 ) | ( ~n1076 & n1077 ) ;
  assign n1079 = ( n980 & ~n1047 ) | ( n980 & n1078 ) | ( ~n1047 & n1078 ) ;
  assign n1080 = ( n980 & n1047 ) | ( n980 & n1078 ) | ( n1047 & n1078 ) ;
  assign n1081 = ( n1047 & n1079 ) | ( n1047 & ~n1080 ) | ( n1079 & ~n1080 ) ;
  assign n1082 = ( n982 & n1037 ) | ( n982 & n1081 ) | ( n1037 & n1081 ) ;
  assign n1083 = ( ~n982 & n1037 ) | ( ~n982 & n1081 ) | ( n1037 & n1081 ) ;
  assign n1084 = ( n982 & ~n1082 ) | ( n982 & n1083 ) | ( ~n1082 & n1083 ) ;
  assign n1085 = ( n985 & ~n1027 ) | ( n985 & n1084 ) | ( ~n1027 & n1084 ) ;
  assign n1086 = ( n985 & n1027 ) | ( n985 & n1084 ) | ( n1027 & n1084 ) ;
  assign n1087 = ( n1027 & n1085 ) | ( n1027 & ~n1086 ) | ( n1085 & ~n1086 ) ;
  assign n1088 = ( n1002 & n1017 ) | ( n1002 & n1087 ) | ( n1017 & n1087 ) ;
  assign n1089 = ( ~n1002 & n1017 ) | ( ~n1002 & n1087 ) | ( n1017 & n1087 ) ;
  assign n1090 = ( n1002 & ~n1088 ) | ( n1002 & n1089 ) | ( ~n1088 & n1089 ) ;
  assign n1091 = ( ~x82 & x83 ) | ( ~x82 & n1005 ) | ( x83 & n1005 ) ;
  assign n1092 = ( x82 & x83 ) | ( x82 & n1005 ) | ( x83 & n1005 ) ;
  assign n1093 = ( x82 & n1091 ) | ( x82 & ~n1092 ) | ( n1091 & ~n1092 ) ;
  assign n1094 = x0 & n1093 ;
  assign n1095 = ( x1 & x2 ) | ( x1 & n1094 ) | ( x2 & n1094 ) ;
  assign n1096 = x82 & n172 ;
  assign n1097 = ( ~x81 & n135 ) | ( ~x81 & n174 ) | ( n135 & n174 ) ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = x83 & n147 ;
  assign n1100 = n1098 | n1099 ;
  assign n1101 = n1095 | n1100 ;
  assign n1102 = n1095 & n1100 ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = n206 & n840 ;
  assign n1105 = x5 & n1104 ;
  assign n1106 = x80 & n205 ;
  assign n1107 = x79 & n201 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = x78 & n221 ;
  assign n1110 = n1108 | n1109 ;
  assign n1111 = ( ~x5 & n1104 ) | ( ~x5 & n1110 ) | ( n1104 & n1110 ) ;
  assign n1112 = x5 & ~n1110 ;
  assign n1113 = ( ~n1105 & n1111 ) | ( ~n1105 & n1112 ) | ( n1111 & n1112 ) ;
  assign n1114 = n301 & n626 ;
  assign n1115 = x8 & n1114 ;
  assign n1116 = x77 & n309 ;
  assign n1117 = x76 & n306 ;
  assign n1118 = n1116 | n1117 ;
  assign n1119 = x75 & n359 ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = ( ~x8 & n1114 ) | ( ~x8 & n1120 ) | ( n1114 & n1120 ) ;
  assign n1122 = x8 & ~n1120 ;
  assign n1123 = ( ~n1115 & n1121 ) | ( ~n1115 & n1122 ) | ( n1121 & n1122 ) ;
  assign n1124 = n436 & n449 ;
  assign n1125 = x11 & n1124 ;
  assign n1126 = x74 & n456 ;
  assign n1127 = x73 & n453 ;
  assign n1128 = n1126 | n1127 ;
  assign n1129 = x72 & n536 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = ( ~x11 & n1124 ) | ( ~x11 & n1130 ) | ( n1124 & n1130 ) ;
  assign n1132 = x11 & ~n1130 ;
  assign n1133 = ( ~n1125 & n1131 ) | ( ~n1125 & n1132 ) | ( n1131 & n1132 ) ;
  assign n1134 = n193 & n874 ;
  assign n1135 = x17 & n1134 ;
  assign n1136 = x68 & n881 ;
  assign n1137 = x67 & n878 ;
  assign n1138 = n1136 | n1137 ;
  assign n1139 = x66 & n959 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = ( ~x17 & n1134 ) | ( ~x17 & n1140 ) | ( n1134 & n1140 ) ;
  assign n1142 = x17 & ~n1140 ;
  assign n1143 = ( ~n1135 & n1141 ) | ( ~n1135 & n1142 ) | ( n1141 & n1142 ) ;
  assign n1144 = ~x19 & x20 ;
  assign n1145 = x19 & ~x20 ;
  assign n1146 = ( n1069 & n1144 ) | ( n1069 & n1145 ) | ( n1144 & n1145 ) ;
  assign n1147 = n302 & n1146 ;
  assign n1148 = ~x17 & x19 ;
  assign n1149 = x18 & x19 ;
  assign n1150 = ( n1068 & n1148 ) | ( n1068 & ~n1149 ) | ( n1148 & ~n1149 ) ;
  assign n1151 = x64 & n1150 ;
  assign n1152 = n1147 | n1151 ;
  assign n1153 = n1069 & ~n1146 ;
  assign n1154 = x65 & n1153 ;
  assign n1155 = n1152 | n1154 ;
  assign n1156 = n1070 | n1155 ;
  assign n1157 = ( x20 & n1070 ) | ( x20 & ~n1155 ) | ( n1070 & ~n1155 ) ;
  assign n1158 = x20 & ~n1155 ;
  assign n1159 = ( n1156 & ~n1157 ) | ( n1156 & n1158 ) | ( ~n1157 & n1158 ) ;
  assign n1160 = ( ~n1074 & n1143 ) | ( ~n1074 & n1159 ) | ( n1143 & n1159 ) ;
  assign n1161 = ( n1074 & n1143 ) | ( n1074 & n1159 ) | ( n1143 & n1159 ) ;
  assign n1162 = ( n1074 & n1160 ) | ( n1074 & ~n1161 ) | ( n1160 & ~n1161 ) ;
  assign n1163 = n322 & n649 ;
  assign n1164 = x14 & n1163 ;
  assign n1165 = x71 & n656 ;
  assign n1166 = x70 & n653 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = x69 & n744 ;
  assign n1169 = n1167 | n1168 ;
  assign n1170 = ( ~x14 & n1163 ) | ( ~x14 & n1169 ) | ( n1163 & n1169 ) ;
  assign n1171 = x14 & ~n1169 ;
  assign n1172 = ( ~n1164 & n1170 ) | ( ~n1164 & n1171 ) | ( n1170 & n1171 ) ;
  assign n1173 = ( n1076 & n1162 ) | ( n1076 & n1172 ) | ( n1162 & n1172 ) ;
  assign n1174 = ( ~n1076 & n1162 ) | ( ~n1076 & n1172 ) | ( n1162 & n1172 ) ;
  assign n1175 = ( n1076 & ~n1173 ) | ( n1076 & n1174 ) | ( ~n1173 & n1174 ) ;
  assign n1176 = ( n1080 & ~n1133 ) | ( n1080 & n1175 ) | ( ~n1133 & n1175 ) ;
  assign n1177 = ( n1080 & n1133 ) | ( n1080 & n1175 ) | ( n1133 & n1175 ) ;
  assign n1178 = ( n1133 & n1176 ) | ( n1133 & ~n1177 ) | ( n1176 & ~n1177 ) ;
  assign n1179 = ( ~n1082 & n1123 ) | ( ~n1082 & n1178 ) | ( n1123 & n1178 ) ;
  assign n1180 = ( n1082 & n1123 ) | ( n1082 & n1178 ) | ( n1123 & n1178 ) ;
  assign n1181 = ( n1082 & n1179 ) | ( n1082 & ~n1180 ) | ( n1179 & ~n1180 ) ;
  assign n1182 = ( n1086 & ~n1113 ) | ( n1086 & n1181 ) | ( ~n1113 & n1181 ) ;
  assign n1183 = ( n1086 & n1113 ) | ( n1086 & n1181 ) | ( n1113 & n1181 ) ;
  assign n1184 = ( n1113 & n1182 ) | ( n1113 & ~n1183 ) | ( n1182 & ~n1183 ) ;
  assign n1185 = ( n1088 & n1103 ) | ( n1088 & n1184 ) | ( n1103 & n1184 ) ;
  assign n1186 = ( ~n1088 & n1103 ) | ( ~n1088 & n1184 ) | ( n1103 & n1184 ) ;
  assign n1187 = ( n1088 & ~n1185 ) | ( n1088 & n1186 ) | ( ~n1185 & n1186 ) ;
  assign n1188 = ( ~x83 & x84 ) | ( ~x83 & n1092 ) | ( x84 & n1092 ) ;
  assign n1189 = ( x83 & x84 ) | ( x83 & n1092 ) | ( x84 & n1092 ) ;
  assign n1190 = ( x83 & n1188 ) | ( x83 & ~n1189 ) | ( n1188 & ~n1189 ) ;
  assign n1191 = x0 & n1190 ;
  assign n1192 = ( x1 & x2 ) | ( x1 & n1191 ) | ( x2 & n1191 ) ;
  assign n1193 = x83 & n172 ;
  assign n1194 = ( ~x82 & n135 ) | ( ~x82 & n174 ) | ( n135 & n174 ) ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = x84 & n147 ;
  assign n1197 = n1195 | n1196 ;
  assign n1198 = n1192 | n1197 ;
  assign n1199 = n1192 & n1197 ;
  assign n1200 = n1198 & ~n1199 ;
  assign n1201 = n301 & n697 ;
  assign n1202 = x8 & n1201 ;
  assign n1203 = x78 & n309 ;
  assign n1204 = x77 & n306 ;
  assign n1205 = n1203 | n1204 ;
  assign n1206 = x76 & n359 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = ( ~x8 & n1201 ) | ( ~x8 & n1207 ) | ( n1201 & n1207 ) ;
  assign n1209 = x8 & ~n1207 ;
  assign n1210 = ( ~n1202 & n1208 ) | ( ~n1202 & n1209 ) | ( n1208 & n1209 ) ;
  assign n1211 = x66 & n1153 ;
  assign n1212 = x65 & n1150 ;
  assign n1213 = n1211 | n1212 ;
  assign n1214 = n226 & n1146 ;
  assign n1215 = n1068 & n1145 ;
  assign n1216 = ~n1067 & n1144 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = x64 & ~n1217 ;
  assign n1219 = ( x64 & n1214 ) | ( x64 & ~n1218 ) | ( n1214 & ~n1218 ) ;
  assign n1220 = n1213 | n1219 ;
  assign n1221 = ~x20 & n1220 ;
  assign n1222 = ( x20 & n1156 ) | ( x20 & n1220 ) | ( n1156 & n1220 ) ;
  assign n1223 = n1156 & n1220 ;
  assign n1224 = ( n1221 & n1222 ) | ( n1221 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1225 = n240 & n874 ;
  assign n1226 = x17 & n1225 ;
  assign n1227 = x69 & n881 ;
  assign n1228 = x68 & n878 ;
  assign n1229 = n1227 | n1228 ;
  assign n1230 = x67 & n959 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = ( ~x17 & n1225 ) | ( ~x17 & n1231 ) | ( n1225 & n1231 ) ;
  assign n1233 = x17 & ~n1231 ;
  assign n1234 = ( ~n1226 & n1232 ) | ( ~n1226 & n1233 ) | ( n1232 & n1233 ) ;
  assign n1235 = ( n1161 & n1224 ) | ( n1161 & n1234 ) | ( n1224 & n1234 ) ;
  assign n1236 = ( ~n1161 & n1224 ) | ( ~n1161 & n1234 ) | ( n1224 & n1234 ) ;
  assign n1237 = ( n1161 & ~n1235 ) | ( n1161 & n1236 ) | ( ~n1235 & n1236 ) ;
  assign n1238 = n372 & n649 ;
  assign n1239 = x14 & n1238 ;
  assign n1240 = x72 & n656 ;
  assign n1241 = x71 & n653 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = x70 & n744 ;
  assign n1244 = n1242 | n1243 ;
  assign n1245 = ( ~x14 & n1238 ) | ( ~x14 & n1244 ) | ( n1238 & n1244 ) ;
  assign n1246 = x14 & ~n1244 ;
  assign n1247 = ( ~n1239 & n1245 ) | ( ~n1239 & n1246 ) | ( n1245 & n1246 ) ;
  assign n1248 = ( n1173 & ~n1237 ) | ( n1173 & n1247 ) | ( ~n1237 & n1247 ) ;
  assign n1249 = ( n1173 & n1237 ) | ( n1173 & n1247 ) | ( n1237 & n1247 ) ;
  assign n1250 = ( n1237 & n1248 ) | ( n1237 & ~n1249 ) | ( n1248 & ~n1249 ) ;
  assign n1251 = n449 & n508 ;
  assign n1252 = x11 & n1251 ;
  assign n1253 = x75 & n456 ;
  assign n1254 = x74 & n453 ;
  assign n1255 = n1253 | n1254 ;
  assign n1256 = x73 & n536 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = ( ~x11 & n1251 ) | ( ~x11 & n1257 ) | ( n1251 & n1257 ) ;
  assign n1259 = x11 & ~n1257 ;
  assign n1260 = ( ~n1252 & n1258 ) | ( ~n1252 & n1259 ) | ( n1258 & n1259 ) ;
  assign n1261 = ( n1177 & ~n1250 ) | ( n1177 & n1260 ) | ( ~n1250 & n1260 ) ;
  assign n1262 = ( n1177 & n1250 ) | ( n1177 & n1260 ) | ( n1250 & n1260 ) ;
  assign n1263 = ( n1250 & n1261 ) | ( n1250 & ~n1262 ) | ( n1261 & ~n1262 ) ;
  assign n1264 = ( n1180 & n1210 ) | ( n1180 & n1263 ) | ( n1210 & n1263 ) ;
  assign n1265 = ( ~n1180 & n1210 ) | ( ~n1180 & n1263 ) | ( n1210 & n1263 ) ;
  assign n1266 = ( n1180 & ~n1264 ) | ( n1180 & n1265 ) | ( ~n1264 & n1265 ) ;
  assign n1267 = n206 & n990 ;
  assign n1268 = x5 & n1267 ;
  assign n1269 = x81 & n205 ;
  assign n1270 = x80 & n201 ;
  assign n1271 = n1269 | n1270 ;
  assign n1272 = x79 & n221 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = ( ~x5 & n1267 ) | ( ~x5 & n1273 ) | ( n1267 & n1273 ) ;
  assign n1275 = x5 & ~n1273 ;
  assign n1276 = ( ~n1268 & n1274 ) | ( ~n1268 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1277 = ( n1183 & ~n1266 ) | ( n1183 & n1276 ) | ( ~n1266 & n1276 ) ;
  assign n1278 = ( n1183 & n1266 ) | ( n1183 & n1276 ) | ( n1266 & n1276 ) ;
  assign n1279 = ( n1266 & n1277 ) | ( n1266 & ~n1278 ) | ( n1277 & ~n1278 ) ;
  assign n1280 = ( n1185 & n1200 ) | ( n1185 & n1279 ) | ( n1200 & n1279 ) ;
  assign n1281 = ( ~n1185 & n1200 ) | ( ~n1185 & n1279 ) | ( n1200 & n1279 ) ;
  assign n1282 = ( n1185 & ~n1280 ) | ( n1185 & n1281 ) | ( ~n1280 & n1281 ) ;
  assign n1283 = n449 & n565 ;
  assign n1284 = x11 & n1283 ;
  assign n1285 = x76 & n456 ;
  assign n1286 = x75 & n453 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = x74 & n536 ;
  assign n1289 = n1287 | n1288 ;
  assign n1290 = ( ~x11 & n1283 ) | ( ~x11 & n1289 ) | ( n1283 & n1289 ) ;
  assign n1291 = x11 & ~n1289 ;
  assign n1292 = ( ~n1284 & n1290 ) | ( ~n1284 & n1291 ) | ( n1290 & n1291 ) ;
  assign n1293 = n276 & n874 ;
  assign n1294 = x17 & n1293 ;
  assign n1295 = x70 & n881 ;
  assign n1296 = x69 & n878 ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = x68 & n959 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = ( ~x17 & n1293 ) | ( ~x17 & n1299 ) | ( n1293 & n1299 ) ;
  assign n1301 = x17 & ~n1299 ;
  assign n1302 = ( ~n1294 & n1300 ) | ( ~n1294 & n1301 ) | ( n1300 & n1301 ) ;
  assign n1303 = n1156 | n1220 ;
  assign n1304 = x20 & n1303 ;
  assign n1305 = x67 & n1153 ;
  assign n1306 = x66 & n1150 ;
  assign n1307 = x65 & n1217 ;
  assign n1308 = n1306 | n1307 ;
  assign n1309 = n1305 | n1308 ;
  assign n1310 = n169 & n1146 ;
  assign n1311 = n1309 | n1310 ;
  assign n1312 = x20 | x21 ;
  assign n1313 = x20 & x21 ;
  assign n1314 = n1312 & ~n1313 ;
  assign n1315 = x64 & n1314 ;
  assign n1316 = ( n1304 & ~n1311 ) | ( n1304 & n1315 ) | ( ~n1311 & n1315 ) ;
  assign n1317 = x20 & ~n1311 ;
  assign n1318 = ( ~n1304 & n1311 ) | ( ~n1304 & n1317 ) | ( n1311 & n1317 ) ;
  assign n1319 = ( n1315 & n1317 ) | ( n1315 & n1318 ) | ( n1317 & n1318 ) ;
  assign n1320 = ( n1316 & n1318 ) | ( n1316 & ~n1319 ) | ( n1318 & ~n1319 ) ;
  assign n1321 = ( n1235 & n1302 ) | ( n1235 & n1320 ) | ( n1302 & n1320 ) ;
  assign n1322 = ( ~n1235 & n1302 ) | ( ~n1235 & n1320 ) | ( n1302 & n1320 ) ;
  assign n1323 = ( n1235 & ~n1321 ) | ( n1235 & n1322 ) | ( ~n1321 & n1322 ) ;
  assign n1324 = n388 & n649 ;
  assign n1325 = x14 & n1324 ;
  assign n1326 = x73 & n656 ;
  assign n1327 = x72 & n653 ;
  assign n1328 = n1326 | n1327 ;
  assign n1329 = x71 & n744 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = ( ~x14 & n1324 ) | ( ~x14 & n1330 ) | ( n1324 & n1330 ) ;
  assign n1332 = x14 & ~n1330 ;
  assign n1333 = ( ~n1325 & n1331 ) | ( ~n1325 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ( n1249 & ~n1323 ) | ( n1249 & n1333 ) | ( ~n1323 & n1333 ) ;
  assign n1335 = ( n1249 & n1323 ) | ( n1249 & n1333 ) | ( n1323 & n1333 ) ;
  assign n1336 = ( n1323 & n1334 ) | ( n1323 & ~n1335 ) | ( n1334 & ~n1335 ) ;
  assign n1337 = ( n1262 & n1292 ) | ( n1262 & n1336 ) | ( n1292 & n1336 ) ;
  assign n1338 = ( ~n1262 & n1292 ) | ( ~n1262 & n1336 ) | ( n1292 & n1336 ) ;
  assign n1339 = ( n1262 & ~n1337 ) | ( n1262 & n1338 ) | ( ~n1337 & n1338 ) ;
  assign n1340 = n301 & n823 ;
  assign n1341 = x8 & n1340 ;
  assign n1342 = x79 & n309 ;
  assign n1343 = x78 & n306 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = x77 & n359 ;
  assign n1346 = n1344 | n1345 ;
  assign n1347 = ( ~x8 & n1340 ) | ( ~x8 & n1346 ) | ( n1340 & n1346 ) ;
  assign n1348 = x8 & ~n1346 ;
  assign n1349 = ( ~n1341 & n1347 ) | ( ~n1341 & n1348 ) | ( n1347 & n1348 ) ;
  assign n1350 = ( n1264 & n1339 ) | ( n1264 & n1349 ) | ( n1339 & n1349 ) ;
  assign n1351 = ( ~n1264 & n1339 ) | ( ~n1264 & n1349 ) | ( n1339 & n1349 ) ;
  assign n1352 = ( n1264 & ~n1350 ) | ( n1264 & n1351 ) | ( ~n1350 & n1351 ) ;
  assign n1353 = n206 & n1006 ;
  assign n1354 = x5 & n1353 ;
  assign n1355 = x82 & n205 ;
  assign n1356 = x81 & n201 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = x80 & n221 ;
  assign n1359 = n1357 | n1358 ;
  assign n1360 = ( ~x5 & n1353 ) | ( ~x5 & n1359 ) | ( n1353 & n1359 ) ;
  assign n1361 = x5 & ~n1359 ;
  assign n1362 = ( ~n1354 & n1360 ) | ( ~n1354 & n1361 ) | ( n1360 & n1361 ) ;
  assign n1363 = ( n1278 & n1352 ) | ( n1278 & n1362 ) | ( n1352 & n1362 ) ;
  assign n1364 = ( ~n1278 & n1352 ) | ( ~n1278 & n1362 ) | ( n1352 & n1362 ) ;
  assign n1365 = ( n1278 & ~n1363 ) | ( n1278 & n1364 ) | ( ~n1363 & n1364 ) ;
  assign n1366 = ( ~x84 & x85 ) | ( ~x84 & n1189 ) | ( x85 & n1189 ) ;
  assign n1367 = ( x84 & x85 ) | ( x84 & n1189 ) | ( x85 & n1189 ) ;
  assign n1368 = ( x84 & n1366 ) | ( x84 & ~n1367 ) | ( n1366 & ~n1367 ) ;
  assign n1369 = x0 & n1368 ;
  assign n1370 = ( x1 & x2 ) | ( x1 & n1369 ) | ( x2 & n1369 ) ;
  assign n1371 = x84 & n172 ;
  assign n1372 = x85 | n1371 ;
  assign n1373 = ( n147 & n1371 ) | ( n147 & n1372 ) | ( n1371 & n1372 ) ;
  assign n1374 = ( ~x83 & n135 ) | ( ~x83 & n174 ) | ( n135 & n174 ) ;
  assign n1375 = n1373 | n1374 ;
  assign n1376 = n1370 | n1375 ;
  assign n1377 = n1370 & n1375 ;
  assign n1378 = n1376 & ~n1377 ;
  assign n1379 = ( n1280 & ~n1365 ) | ( n1280 & n1378 ) | ( ~n1365 & n1378 ) ;
  assign n1380 = ( n1280 & n1365 ) | ( n1280 & n1378 ) | ( n1365 & n1378 ) ;
  assign n1381 = ( n1365 & n1379 ) | ( n1365 & ~n1380 ) | ( n1379 & ~n1380 ) ;
  assign n1382 = ( ~x85 & x86 ) | ( ~x85 & n1367 ) | ( x86 & n1367 ) ;
  assign n1383 = ( x85 & x86 ) | ( x85 & n1367 ) | ( x86 & n1367 ) ;
  assign n1384 = ( x85 & n1382 ) | ( x85 & ~n1383 ) | ( n1382 & ~n1383 ) ;
  assign n1385 = x0 & n1384 ;
  assign n1386 = ( x1 & x2 ) | ( x1 & n1385 ) | ( x2 & n1385 ) ;
  assign n1387 = x85 & n172 ;
  assign n1388 = ( ~x84 & n135 ) | ( ~x84 & n174 ) | ( n135 & n174 ) ;
  assign n1389 = n1387 | n1388 ;
  assign n1390 = x86 & n147 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n1386 | n1391 ;
  assign n1393 = n1386 & n1391 ;
  assign n1394 = n1392 & ~n1393 ;
  assign n1395 = n449 & n626 ;
  assign n1396 = x11 & n1395 ;
  assign n1397 = x77 & n456 ;
  assign n1398 = x76 & n453 ;
  assign n1399 = n1397 | n1398 ;
  assign n1400 = x75 & n536 ;
  assign n1401 = n1399 | n1400 ;
  assign n1402 = ( ~x11 & n1395 ) | ( ~x11 & n1401 ) | ( n1395 & n1401 ) ;
  assign n1403 = x11 & ~n1401 ;
  assign n1404 = ( ~n1396 & n1402 ) | ( ~n1396 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1405 = n436 & n649 ;
  assign n1406 = x14 & n1405 ;
  assign n1407 = x74 & n656 ;
  assign n1408 = x73 & n653 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = x72 & n744 ;
  assign n1411 = n1409 | n1410 ;
  assign n1412 = ( ~x14 & n1405 ) | ( ~x14 & n1411 ) | ( n1405 & n1411 ) ;
  assign n1413 = x14 & ~n1411 ;
  assign n1414 = ( ~n1406 & n1412 ) | ( ~n1406 & n1413 ) | ( n1412 & n1413 ) ;
  assign n1415 = x68 & n1153 ;
  assign n1416 = x66 & n1217 ;
  assign n1417 = n1415 | n1416 ;
  assign n1418 = n193 & n1146 ;
  assign n1419 = n1417 | n1418 ;
  assign n1420 = x67 & n1150 ;
  assign n1421 = ( ~x20 & n1419 ) | ( ~x20 & n1420 ) | ( n1419 & n1420 ) ;
  assign n1422 = ( x20 & ~n1419 ) | ( x20 & n1420 ) | ( ~n1419 & n1420 ) ;
  assign n1423 = ~n1420 & n1422 ;
  assign n1424 = n1421 | n1423 ;
  assign n1425 = ~x22 & x23 ;
  assign n1426 = x22 & ~x23 ;
  assign n1427 = ( n1314 & n1425 ) | ( n1314 & n1426 ) | ( n1425 & n1426 ) ;
  assign n1428 = n302 & n1427 ;
  assign n1429 = ~x20 & x22 ;
  assign n1430 = x21 & x22 ;
  assign n1431 = ( n1313 & n1429 ) | ( n1313 & ~n1430 ) | ( n1429 & ~n1430 ) ;
  assign n1432 = x64 & n1431 ;
  assign n1433 = n1428 | n1432 ;
  assign n1434 = n1314 & ~n1427 ;
  assign n1435 = x65 & n1434 ;
  assign n1436 = n1433 | n1435 ;
  assign n1437 = n1315 | n1436 ;
  assign n1438 = ( x23 & n1315 ) | ( x23 & ~n1436 ) | ( n1315 & ~n1436 ) ;
  assign n1439 = x23 & ~n1436 ;
  assign n1440 = ( n1437 & ~n1438 ) | ( n1437 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1441 = ( ~n1319 & n1424 ) | ( ~n1319 & n1440 ) | ( n1424 & n1440 ) ;
  assign n1442 = ( n1319 & n1424 ) | ( n1319 & n1440 ) | ( n1424 & n1440 ) ;
  assign n1443 = ( n1319 & n1441 ) | ( n1319 & ~n1442 ) | ( n1441 & ~n1442 ) ;
  assign n1444 = n322 & n874 ;
  assign n1445 = x17 & n1444 ;
  assign n1446 = x71 & n881 ;
  assign n1447 = x70 & n878 ;
  assign n1448 = n1446 | n1447 ;
  assign n1449 = x69 & n959 ;
  assign n1450 = n1448 | n1449 ;
  assign n1451 = ( ~x17 & n1444 ) | ( ~x17 & n1450 ) | ( n1444 & n1450 ) ;
  assign n1452 = x17 & ~n1450 ;
  assign n1453 = ( ~n1445 & n1451 ) | ( ~n1445 & n1452 ) | ( n1451 & n1452 ) ;
  assign n1454 = ( n1321 & ~n1443 ) | ( n1321 & n1453 ) | ( ~n1443 & n1453 ) ;
  assign n1455 = ( n1321 & n1443 ) | ( n1321 & n1453 ) | ( n1443 & n1453 ) ;
  assign n1456 = ( n1443 & n1454 ) | ( n1443 & ~n1455 ) | ( n1454 & ~n1455 ) ;
  assign n1457 = ( n1335 & n1414 ) | ( n1335 & n1456 ) | ( n1414 & n1456 ) ;
  assign n1458 = ( ~n1335 & n1414 ) | ( ~n1335 & n1456 ) | ( n1414 & n1456 ) ;
  assign n1459 = ( n1335 & ~n1457 ) | ( n1335 & n1458 ) | ( ~n1457 & n1458 ) ;
  assign n1460 = ( n1337 & n1404 ) | ( n1337 & n1459 ) | ( n1404 & n1459 ) ;
  assign n1461 = ( ~n1337 & n1404 ) | ( ~n1337 & n1459 ) | ( n1404 & n1459 ) ;
  assign n1462 = ( n1337 & ~n1460 ) | ( n1337 & n1461 ) | ( ~n1460 & n1461 ) ;
  assign n1463 = n301 & n840 ;
  assign n1464 = x8 & n1463 ;
  assign n1465 = x80 & n309 ;
  assign n1466 = x79 & n306 ;
  assign n1467 = n1465 | n1466 ;
  assign n1468 = x78 & n359 ;
  assign n1469 = n1467 | n1468 ;
  assign n1470 = ( ~x8 & n1463 ) | ( ~x8 & n1469 ) | ( n1463 & n1469 ) ;
  assign n1471 = x8 & ~n1469 ;
  assign n1472 = ( ~n1464 & n1470 ) | ( ~n1464 & n1471 ) | ( n1470 & n1471 ) ;
  assign n1473 = ( n1350 & ~n1462 ) | ( n1350 & n1472 ) | ( ~n1462 & n1472 ) ;
  assign n1474 = ( n1350 & n1462 ) | ( n1350 & n1472 ) | ( n1462 & n1472 ) ;
  assign n1475 = ( n1462 & n1473 ) | ( n1462 & ~n1474 ) | ( n1473 & ~n1474 ) ;
  assign n1476 = n206 & n1093 ;
  assign n1477 = x5 & n1476 ;
  assign n1478 = x83 & n205 ;
  assign n1479 = x82 & n201 ;
  assign n1480 = n1478 | n1479 ;
  assign n1481 = x81 & n221 ;
  assign n1482 = n1480 | n1481 ;
  assign n1483 = ( ~x5 & n1476 ) | ( ~x5 & n1482 ) | ( n1476 & n1482 ) ;
  assign n1484 = x5 & ~n1482 ;
  assign n1485 = ( ~n1477 & n1483 ) | ( ~n1477 & n1484 ) | ( n1483 & n1484 ) ;
  assign n1486 = ( n1363 & ~n1475 ) | ( n1363 & n1485 ) | ( ~n1475 & n1485 ) ;
  assign n1487 = ( n1363 & n1475 ) | ( n1363 & n1485 ) | ( n1475 & n1485 ) ;
  assign n1488 = ( n1475 & n1486 ) | ( n1475 & ~n1487 ) | ( n1486 & ~n1487 ) ;
  assign n1489 = ( n1380 & n1394 ) | ( n1380 & n1488 ) | ( n1394 & n1488 ) ;
  assign n1490 = ( ~n1380 & n1394 ) | ( ~n1380 & n1488 ) | ( n1394 & n1488 ) ;
  assign n1491 = ( n1380 & ~n1489 ) | ( n1380 & n1490 ) | ( ~n1489 & n1490 ) ;
  assign n1492 = ( ~x86 & x87 ) | ( ~x86 & n1383 ) | ( x87 & n1383 ) ;
  assign n1493 = ( x86 & x87 ) | ( x86 & n1383 ) | ( x87 & n1383 ) ;
  assign n1494 = ( x86 & n1492 ) | ( x86 & ~n1493 ) | ( n1492 & ~n1493 ) ;
  assign n1495 = x0 & n1494 ;
  assign n1496 = ( x1 & x2 ) | ( x1 & n1495 ) | ( x2 & n1495 ) ;
  assign n1497 = x86 & n172 ;
  assign n1498 = x87 | n1497 ;
  assign n1499 = ( n147 & n1497 ) | ( n147 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1500 = ( ~x85 & n135 ) | ( ~x85 & n174 ) | ( n135 & n174 ) ;
  assign n1501 = n1499 | n1500 ;
  assign n1502 = n1496 | n1501 ;
  assign n1503 = n1496 & n1501 ;
  assign n1504 = n1502 & ~n1503 ;
  assign n1505 = n449 & n697 ;
  assign n1506 = x11 & n1505 ;
  assign n1507 = x78 & n456 ;
  assign n1508 = x77 & n453 ;
  assign n1509 = n1507 | n1508 ;
  assign n1510 = x76 & n536 ;
  assign n1511 = n1509 | n1510 ;
  assign n1512 = ( ~x11 & n1505 ) | ( ~x11 & n1511 ) | ( n1505 & n1511 ) ;
  assign n1513 = x11 & ~n1511 ;
  assign n1514 = ( ~n1506 & n1512 ) | ( ~n1506 & n1513 ) | ( n1512 & n1513 ) ;
  assign n1515 = n508 & n649 ;
  assign n1516 = x14 & n1515 ;
  assign n1517 = x75 & n656 ;
  assign n1518 = x74 & n653 ;
  assign n1519 = n1517 | n1518 ;
  assign n1520 = x73 & n744 ;
  assign n1521 = n1519 | n1520 ;
  assign n1522 = ( ~x14 & n1515 ) | ( ~x14 & n1521 ) | ( n1515 & n1521 ) ;
  assign n1523 = x14 & ~n1521 ;
  assign n1524 = ( ~n1516 & n1522 ) | ( ~n1516 & n1523 ) | ( n1522 & n1523 ) ;
  assign n1525 = x66 & n1434 ;
  assign n1526 = x65 & n1431 ;
  assign n1527 = n1525 | n1526 ;
  assign n1528 = n226 & n1427 ;
  assign n1529 = n1313 & n1426 ;
  assign n1530 = ~n1312 & n1425 ;
  assign n1531 = n1529 | n1530 ;
  assign n1532 = x64 & ~n1531 ;
  assign n1533 = ( x64 & n1528 ) | ( x64 & ~n1532 ) | ( n1528 & ~n1532 ) ;
  assign n1534 = n1527 | n1533 ;
  assign n1535 = ~x23 & n1534 ;
  assign n1536 = ( x23 & n1437 ) | ( x23 & n1534 ) | ( n1437 & n1534 ) ;
  assign n1537 = n1437 & n1534 ;
  assign n1538 = ( n1535 & n1536 ) | ( n1535 & ~n1537 ) | ( n1536 & ~n1537 ) ;
  assign n1539 = n240 & n1146 ;
  assign n1540 = x20 & n1539 ;
  assign n1541 = x69 & n1153 ;
  assign n1542 = x68 & n1150 ;
  assign n1543 = n1541 | n1542 ;
  assign n1544 = x67 & n1217 ;
  assign n1545 = n1543 | n1544 ;
  assign n1546 = ( ~x20 & n1539 ) | ( ~x20 & n1545 ) | ( n1539 & n1545 ) ;
  assign n1547 = x20 & ~n1545 ;
  assign n1548 = ( ~n1540 & n1546 ) | ( ~n1540 & n1547 ) | ( n1546 & n1547 ) ;
  assign n1549 = ( n1442 & n1538 ) | ( n1442 & n1548 ) | ( n1538 & n1548 ) ;
  assign n1550 = ( ~n1442 & n1538 ) | ( ~n1442 & n1548 ) | ( n1538 & n1548 ) ;
  assign n1551 = ( n1442 & ~n1549 ) | ( n1442 & n1550 ) | ( ~n1549 & n1550 ) ;
  assign n1552 = n372 & n874 ;
  assign n1553 = x17 & n1552 ;
  assign n1554 = x72 & n881 ;
  assign n1555 = x71 & n878 ;
  assign n1556 = n1554 | n1555 ;
  assign n1557 = x70 & n959 ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = ( ~x17 & n1552 ) | ( ~x17 & n1558 ) | ( n1552 & n1558 ) ;
  assign n1560 = x17 & ~n1558 ;
  assign n1561 = ( ~n1553 & n1559 ) | ( ~n1553 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1562 = ( n1455 & ~n1551 ) | ( n1455 & n1561 ) | ( ~n1551 & n1561 ) ;
  assign n1563 = ( n1455 & n1551 ) | ( n1455 & n1561 ) | ( n1551 & n1561 ) ;
  assign n1564 = ( n1551 & n1562 ) | ( n1551 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n1565 = ( n1457 & n1524 ) | ( n1457 & n1564 ) | ( n1524 & n1564 ) ;
  assign n1566 = ( ~n1457 & n1524 ) | ( ~n1457 & n1564 ) | ( n1524 & n1564 ) ;
  assign n1567 = ( n1457 & ~n1565 ) | ( n1457 & n1566 ) | ( ~n1565 & n1566 ) ;
  assign n1568 = ( n1460 & n1514 ) | ( n1460 & n1567 ) | ( n1514 & n1567 ) ;
  assign n1569 = ( ~n1460 & n1514 ) | ( ~n1460 & n1567 ) | ( n1514 & n1567 ) ;
  assign n1570 = ( n1460 & ~n1568 ) | ( n1460 & n1569 ) | ( ~n1568 & n1569 ) ;
  assign n1571 = n301 & n990 ;
  assign n1572 = x8 & n1571 ;
  assign n1573 = x81 & n309 ;
  assign n1574 = x80 & n306 ;
  assign n1575 = n1573 | n1574 ;
  assign n1576 = x79 & n359 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = ( ~x8 & n1571 ) | ( ~x8 & n1577 ) | ( n1571 & n1577 ) ;
  assign n1579 = x8 & ~n1577 ;
  assign n1580 = ( ~n1572 & n1578 ) | ( ~n1572 & n1579 ) | ( n1578 & n1579 ) ;
  assign n1581 = ( n1474 & ~n1570 ) | ( n1474 & n1580 ) | ( ~n1570 & n1580 ) ;
  assign n1582 = ( n1474 & n1570 ) | ( n1474 & n1580 ) | ( n1570 & n1580 ) ;
  assign n1583 = ( n1570 & n1581 ) | ( n1570 & ~n1582 ) | ( n1581 & ~n1582 ) ;
  assign n1584 = n206 & n1190 ;
  assign n1585 = x5 & n1584 ;
  assign n1586 = x84 & n205 ;
  assign n1587 = x83 & n201 ;
  assign n1588 = n1586 | n1587 ;
  assign n1589 = x82 & n221 ;
  assign n1590 = n1588 | n1589 ;
  assign n1591 = ( ~x5 & n1584 ) | ( ~x5 & n1590 ) | ( n1584 & n1590 ) ;
  assign n1592 = x5 & ~n1590 ;
  assign n1593 = ( ~n1585 & n1591 ) | ( ~n1585 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = ( n1487 & ~n1583 ) | ( n1487 & n1593 ) | ( ~n1583 & n1593 ) ;
  assign n1595 = ( n1487 & n1583 ) | ( n1487 & n1593 ) | ( n1583 & n1593 ) ;
  assign n1596 = ( n1583 & n1594 ) | ( n1583 & ~n1595 ) | ( n1594 & ~n1595 ) ;
  assign n1597 = ( n1489 & n1504 ) | ( n1489 & n1596 ) | ( n1504 & n1596 ) ;
  assign n1598 = ( ~n1489 & n1504 ) | ( ~n1489 & n1596 ) | ( n1504 & n1596 ) ;
  assign n1599 = ( n1489 & ~n1597 ) | ( n1489 & n1598 ) | ( ~n1597 & n1598 ) ;
  assign n1600 = ( ~x87 & x88 ) | ( ~x87 & n1493 ) | ( x88 & n1493 ) ;
  assign n1601 = ( x87 & x88 ) | ( x87 & n1493 ) | ( x88 & n1493 ) ;
  assign n1602 = ( x87 & n1600 ) | ( x87 & ~n1601 ) | ( n1600 & ~n1601 ) ;
  assign n1603 = x0 & n1602 ;
  assign n1604 = ( x1 & x2 ) | ( x1 & n1603 ) | ( x2 & n1603 ) ;
  assign n1605 = x87 & n172 ;
  assign n1606 = x88 | n1605 ;
  assign n1607 = ( n147 & n1605 ) | ( n147 & n1606 ) | ( n1605 & n1606 ) ;
  assign n1608 = ( ~x86 & n135 ) | ( ~x86 & n174 ) | ( n135 & n174 ) ;
  assign n1609 = n1607 | n1608 ;
  assign n1610 = n1604 | n1609 ;
  assign n1611 = n1604 & n1609 ;
  assign n1612 = n1610 & ~n1611 ;
  assign n1613 = n301 & n1006 ;
  assign n1614 = x8 & n1613 ;
  assign n1615 = x82 & n309 ;
  assign n1616 = x81 & n306 ;
  assign n1617 = n1615 | n1616 ;
  assign n1618 = x80 & n359 ;
  assign n1619 = n1617 | n1618 ;
  assign n1620 = ( ~x8 & n1613 ) | ( ~x8 & n1619 ) | ( n1613 & n1619 ) ;
  assign n1621 = x8 & ~n1619 ;
  assign n1622 = ( ~n1614 & n1620 ) | ( ~n1614 & n1621 ) | ( n1620 & n1621 ) ;
  assign n1623 = n565 & n649 ;
  assign n1624 = x14 & n1623 ;
  assign n1625 = x76 & n656 ;
  assign n1626 = x75 & n653 ;
  assign n1627 = n1625 | n1626 ;
  assign n1628 = x74 & n744 ;
  assign n1629 = n1627 | n1628 ;
  assign n1630 = ( ~x14 & n1623 ) | ( ~x14 & n1629 ) | ( n1623 & n1629 ) ;
  assign n1631 = x14 & ~n1629 ;
  assign n1632 = ( ~n1624 & n1630 ) | ( ~n1624 & n1631 ) | ( n1630 & n1631 ) ;
  assign n1633 = n276 & n1146 ;
  assign n1634 = x20 & n1633 ;
  assign n1635 = x70 & n1153 ;
  assign n1636 = x69 & n1150 ;
  assign n1637 = n1635 | n1636 ;
  assign n1638 = x68 & n1217 ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = ( ~x20 & n1633 ) | ( ~x20 & n1639 ) | ( n1633 & n1639 ) ;
  assign n1641 = x20 & ~n1639 ;
  assign n1642 = ( ~n1634 & n1640 ) | ( ~n1634 & n1641 ) | ( n1640 & n1641 ) ;
  assign n1643 = n1437 | n1534 ;
  assign n1644 = x23 & n1643 ;
  assign n1645 = x66 & n1431 ;
  assign n1646 = x67 & n1434 ;
  assign n1647 = x65 & n1531 ;
  assign n1648 = n1646 | n1647 ;
  assign n1649 = n169 & n1427 ;
  assign n1650 = n1648 | n1649 ;
  assign n1651 = n1645 | n1650 ;
  assign n1652 = x23 & x24 ;
  assign n1653 = x23 | x24 ;
  assign n1654 = ~n1652 & n1653 ;
  assign n1655 = x64 & n1654 ;
  assign n1656 = ( n1644 & ~n1651 ) | ( n1644 & n1655 ) | ( ~n1651 & n1655 ) ;
  assign n1657 = x23 & ~n1651 ;
  assign n1658 = ( ~n1644 & n1651 ) | ( ~n1644 & n1657 ) | ( n1651 & n1657 ) ;
  assign n1659 = ( n1655 & n1657 ) | ( n1655 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = ( n1656 & n1658 ) | ( n1656 & ~n1659 ) | ( n1658 & ~n1659 ) ;
  assign n1661 = ( n1549 & n1642 ) | ( n1549 & n1660 ) | ( n1642 & n1660 ) ;
  assign n1662 = ( ~n1549 & n1642 ) | ( ~n1549 & n1660 ) | ( n1642 & n1660 ) ;
  assign n1663 = ( n1549 & ~n1661 ) | ( n1549 & n1662 ) | ( ~n1661 & n1662 ) ;
  assign n1664 = n388 & n874 ;
  assign n1665 = x17 & n1664 ;
  assign n1666 = x73 & n881 ;
  assign n1667 = x72 & n878 ;
  assign n1668 = n1666 | n1667 ;
  assign n1669 = x71 & n959 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = ( ~x17 & n1664 ) | ( ~x17 & n1670 ) | ( n1664 & n1670 ) ;
  assign n1672 = x17 & ~n1670 ;
  assign n1673 = ( ~n1665 & n1671 ) | ( ~n1665 & n1672 ) | ( n1671 & n1672 ) ;
  assign n1674 = ( n1563 & ~n1663 ) | ( n1563 & n1673 ) | ( ~n1663 & n1673 ) ;
  assign n1675 = ( n1563 & n1663 ) | ( n1563 & n1673 ) | ( n1663 & n1673 ) ;
  assign n1676 = ( n1663 & n1674 ) | ( n1663 & ~n1675 ) | ( n1674 & ~n1675 ) ;
  assign n1677 = ( n1565 & n1632 ) | ( n1565 & n1676 ) | ( n1632 & n1676 ) ;
  assign n1678 = ( ~n1565 & n1632 ) | ( ~n1565 & n1676 ) | ( n1632 & n1676 ) ;
  assign n1679 = ( n1565 & ~n1677 ) | ( n1565 & n1678 ) | ( ~n1677 & n1678 ) ;
  assign n1680 = n449 & n823 ;
  assign n1681 = x11 & n1680 ;
  assign n1682 = x79 & n456 ;
  assign n1683 = x78 & n453 ;
  assign n1684 = n1682 | n1683 ;
  assign n1685 = x77 & n536 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = ( ~x11 & n1680 ) | ( ~x11 & n1686 ) | ( n1680 & n1686 ) ;
  assign n1688 = x11 & ~n1686 ;
  assign n1689 = ( ~n1681 & n1687 ) | ( ~n1681 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1690 = ( n1568 & ~n1679 ) | ( n1568 & n1689 ) | ( ~n1679 & n1689 ) ;
  assign n1691 = ( n1568 & n1679 ) | ( n1568 & n1689 ) | ( n1679 & n1689 ) ;
  assign n1692 = ( n1679 & n1690 ) | ( n1679 & ~n1691 ) | ( n1690 & ~n1691 ) ;
  assign n1693 = ( n1582 & n1622 ) | ( n1582 & n1692 ) | ( n1622 & n1692 ) ;
  assign n1694 = ( ~n1582 & n1622 ) | ( ~n1582 & n1692 ) | ( n1622 & n1692 ) ;
  assign n1695 = ( n1582 & ~n1693 ) | ( n1582 & n1694 ) | ( ~n1693 & n1694 ) ;
  assign n1696 = n206 & n1368 ;
  assign n1697 = x5 & n1696 ;
  assign n1698 = x84 & n201 ;
  assign n1699 = x83 & n221 ;
  assign n1700 = n1698 | n1699 ;
  assign n1701 = x85 & n205 ;
  assign n1702 = n1700 | n1701 ;
  assign n1703 = ( ~x5 & n1696 ) | ( ~x5 & n1702 ) | ( n1696 & n1702 ) ;
  assign n1704 = x5 & ~n1702 ;
  assign n1705 = ( ~n1697 & n1703 ) | ( ~n1697 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ( n1595 & ~n1695 ) | ( n1595 & n1705 ) | ( ~n1695 & n1705 ) ;
  assign n1707 = ( n1595 & n1695 ) | ( n1595 & n1705 ) | ( n1695 & n1705 ) ;
  assign n1708 = ( n1695 & n1706 ) | ( n1695 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1709 = ( n1597 & n1612 ) | ( n1597 & n1708 ) | ( n1612 & n1708 ) ;
  assign n1710 = ( ~n1597 & n1612 ) | ( ~n1597 & n1708 ) | ( n1612 & n1708 ) ;
  assign n1711 = ( n1597 & ~n1709 ) | ( n1597 & n1710 ) | ( ~n1709 & n1710 ) ;
  assign n1712 = n206 & n1384 ;
  assign n1713 = x5 & n1712 ;
  assign n1714 = x86 & n205 ;
  assign n1715 = x85 & n201 ;
  assign n1716 = n1714 | n1715 ;
  assign n1717 = x84 & n221 ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = ( ~x5 & n1712 ) | ( ~x5 & n1718 ) | ( n1712 & n1718 ) ;
  assign n1720 = x5 & ~n1718 ;
  assign n1721 = ( ~n1713 & n1719 ) | ( ~n1713 & n1720 ) | ( n1719 & n1720 ) ;
  assign n1722 = n449 & n840 ;
  assign n1723 = x11 & n1722 ;
  assign n1724 = x80 & n456 ;
  assign n1725 = x79 & n453 ;
  assign n1726 = n1724 | n1725 ;
  assign n1727 = x78 & n536 ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = ( ~x11 & n1722 ) | ( ~x11 & n1728 ) | ( n1722 & n1728 ) ;
  assign n1730 = x11 & ~n1728 ;
  assign n1731 = ( ~n1723 & n1729 ) | ( ~n1723 & n1730 ) | ( n1729 & n1730 ) ;
  assign n1732 = n436 & n874 ;
  assign n1733 = x17 & n1732 ;
  assign n1734 = x74 & n881 ;
  assign n1735 = x73 & n878 ;
  assign n1736 = n1734 | n1735 ;
  assign n1737 = x72 & n959 ;
  assign n1738 = n1736 | n1737 ;
  assign n1739 = ( ~x17 & n1732 ) | ( ~x17 & n1738 ) | ( n1732 & n1738 ) ;
  assign n1740 = x17 & ~n1738 ;
  assign n1741 = ( ~n1733 & n1739 ) | ( ~n1733 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1742 = x68 & n1434 ;
  assign n1743 = x66 & n1531 ;
  assign n1744 = n1742 | n1743 ;
  assign n1745 = n193 & n1427 ;
  assign n1746 = n1744 | n1745 ;
  assign n1747 = x67 & n1431 ;
  assign n1748 = ( ~x23 & n1746 ) | ( ~x23 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1749 = ( x23 & ~n1746 ) | ( x23 & n1747 ) | ( ~n1746 & n1747 ) ;
  assign n1750 = ~n1747 & n1749 ;
  assign n1751 = n1748 | n1750 ;
  assign n1752 = x25 & x26 ;
  assign n1753 = x25 | x26 ;
  assign n1754 = ~n1752 & n1753 ;
  assign n1755 = n1654 & n1754 ;
  assign n1756 = n302 & n1755 ;
  assign n1757 = ~x23 & x25 ;
  assign n1758 = x24 & x25 ;
  assign n1759 = ( n1652 & n1757 ) | ( n1652 & ~n1758 ) | ( n1757 & ~n1758 ) ;
  assign n1760 = x64 & n1759 ;
  assign n1761 = n1756 | n1760 ;
  assign n1762 = ( n1654 & n1752 ) | ( n1654 & ~n1753 ) | ( n1752 & ~n1753 ) ;
  assign n1763 = x65 & n1762 ;
  assign n1764 = n1761 | n1763 ;
  assign n1765 = n1655 | n1764 ;
  assign n1766 = ( x26 & n1655 ) | ( x26 & ~n1764 ) | ( n1655 & ~n1764 ) ;
  assign n1767 = x26 & ~n1764 ;
  assign n1768 = ( n1765 & ~n1766 ) | ( n1765 & n1767 ) | ( ~n1766 & n1767 ) ;
  assign n1769 = ( ~n1659 & n1751 ) | ( ~n1659 & n1768 ) | ( n1751 & n1768 ) ;
  assign n1770 = ( n1659 & n1751 ) | ( n1659 & n1768 ) | ( n1751 & n1768 ) ;
  assign n1771 = ( n1659 & n1769 ) | ( n1659 & ~n1770 ) | ( n1769 & ~n1770 ) ;
  assign n1772 = n322 & n1146 ;
  assign n1773 = x20 & n1772 ;
  assign n1774 = x71 & n1153 ;
  assign n1775 = x70 & n1150 ;
  assign n1776 = n1774 | n1775 ;
  assign n1777 = x69 & n1217 ;
  assign n1778 = n1776 | n1777 ;
  assign n1779 = ( ~x20 & n1772 ) | ( ~x20 & n1778 ) | ( n1772 & n1778 ) ;
  assign n1780 = x20 & ~n1778 ;
  assign n1781 = ( ~n1773 & n1779 ) | ( ~n1773 & n1780 ) | ( n1779 & n1780 ) ;
  assign n1782 = ( n1661 & ~n1771 ) | ( n1661 & n1781 ) | ( ~n1771 & n1781 ) ;
  assign n1783 = ( n1661 & n1771 ) | ( n1661 & n1781 ) | ( n1771 & n1781 ) ;
  assign n1784 = ( n1771 & n1782 ) | ( n1771 & ~n1783 ) | ( n1782 & ~n1783 ) ;
  assign n1785 = ( n1675 & n1741 ) | ( n1675 & n1784 ) | ( n1741 & n1784 ) ;
  assign n1786 = ( ~n1675 & n1741 ) | ( ~n1675 & n1784 ) | ( n1741 & n1784 ) ;
  assign n1787 = ( n1675 & ~n1785 ) | ( n1675 & n1786 ) | ( ~n1785 & n1786 ) ;
  assign n1788 = n626 & n649 ;
  assign n1789 = x14 & n1788 ;
  assign n1790 = x77 & n656 ;
  assign n1791 = x76 & n653 ;
  assign n1792 = n1790 | n1791 ;
  assign n1793 = x75 & n744 ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = ( ~x14 & n1788 ) | ( ~x14 & n1794 ) | ( n1788 & n1794 ) ;
  assign n1796 = x14 & ~n1794 ;
  assign n1797 = ( ~n1789 & n1795 ) | ( ~n1789 & n1796 ) | ( n1795 & n1796 ) ;
  assign n1798 = ( n1677 & ~n1787 ) | ( n1677 & n1797 ) | ( ~n1787 & n1797 ) ;
  assign n1799 = ( n1677 & n1787 ) | ( n1677 & n1797 ) | ( n1787 & n1797 ) ;
  assign n1800 = ( n1787 & n1798 ) | ( n1787 & ~n1799 ) | ( n1798 & ~n1799 ) ;
  assign n1801 = ( n1691 & n1731 ) | ( n1691 & n1800 ) | ( n1731 & n1800 ) ;
  assign n1802 = ( ~n1691 & n1731 ) | ( ~n1691 & n1800 ) | ( n1731 & n1800 ) ;
  assign n1803 = ( n1691 & ~n1801 ) | ( n1691 & n1802 ) | ( ~n1801 & n1802 ) ;
  assign n1804 = n301 & n1093 ;
  assign n1805 = x8 & n1804 ;
  assign n1806 = x83 & n309 ;
  assign n1807 = x82 & n306 ;
  assign n1808 = n1806 | n1807 ;
  assign n1809 = x81 & n359 ;
  assign n1810 = n1808 | n1809 ;
  assign n1811 = ( ~x8 & n1804 ) | ( ~x8 & n1810 ) | ( n1804 & n1810 ) ;
  assign n1812 = x8 & ~n1810 ;
  assign n1813 = ( ~n1805 & n1811 ) | ( ~n1805 & n1812 ) | ( n1811 & n1812 ) ;
  assign n1814 = ( n1693 & ~n1803 ) | ( n1693 & n1813 ) | ( ~n1803 & n1813 ) ;
  assign n1815 = ( n1693 & n1803 ) | ( n1693 & n1813 ) | ( n1803 & n1813 ) ;
  assign n1816 = ( n1803 & n1814 ) | ( n1803 & ~n1815 ) | ( n1814 & ~n1815 ) ;
  assign n1817 = ( ~n1707 & n1721 ) | ( ~n1707 & n1816 ) | ( n1721 & n1816 ) ;
  assign n1818 = ( n1707 & n1721 ) | ( n1707 & n1816 ) | ( n1721 & n1816 ) ;
  assign n1819 = ( n1707 & n1817 ) | ( n1707 & ~n1818 ) | ( n1817 & ~n1818 ) ;
  assign n1820 = ( ~x88 & x89 ) | ( ~x88 & n1601 ) | ( x89 & n1601 ) ;
  assign n1821 = ( x88 & x89 ) | ( x88 & n1601 ) | ( x89 & n1601 ) ;
  assign n1822 = ( x88 & n1820 ) | ( x88 & ~n1821 ) | ( n1820 & ~n1821 ) ;
  assign n1823 = x0 & n1822 ;
  assign n1824 = ( x1 & x2 ) | ( x1 & n1823 ) | ( x2 & n1823 ) ;
  assign n1825 = x88 & n172 ;
  assign n1826 = x89 | n1825 ;
  assign n1827 = ( n147 & n1825 ) | ( n147 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1828 = ( ~x87 & n135 ) | ( ~x87 & n174 ) | ( n135 & n174 ) ;
  assign n1829 = n1827 | n1828 ;
  assign n1830 = n1824 | n1829 ;
  assign n1831 = n1824 & n1829 ;
  assign n1832 = n1830 & ~n1831 ;
  assign n1833 = ( n1709 & ~n1819 ) | ( n1709 & n1832 ) | ( ~n1819 & n1832 ) ;
  assign n1834 = ( n1709 & n1819 ) | ( n1709 & n1832 ) | ( n1819 & n1832 ) ;
  assign n1835 = ( n1819 & n1833 ) | ( n1819 & ~n1834 ) | ( n1833 & ~n1834 ) ;
  assign n1836 = ( ~x89 & x90 ) | ( ~x89 & n1821 ) | ( x90 & n1821 ) ;
  assign n1837 = ( x89 & x90 ) | ( x89 & n1821 ) | ( x90 & n1821 ) ;
  assign n1838 = ( x89 & n1836 ) | ( x89 & ~n1837 ) | ( n1836 & ~n1837 ) ;
  assign n1839 = x0 & n1838 ;
  assign n1840 = ( x1 & x2 ) | ( x1 & n1839 ) | ( x2 & n1839 ) ;
  assign n1841 = x89 & n172 ;
  assign n1842 = ( ~x88 & n135 ) | ( ~x88 & n174 ) | ( n135 & n174 ) ;
  assign n1843 = n1841 | n1842 ;
  assign n1844 = x90 & n147 ;
  assign n1845 = n1843 | n1844 ;
  assign n1846 = n1840 | n1845 ;
  assign n1847 = n1840 & n1845 ;
  assign n1848 = n1846 & ~n1847 ;
  assign n1849 = n206 & n1494 ;
  assign n1850 = x5 & n1849 ;
  assign n1851 = x87 & n205 ;
  assign n1852 = x86 & n201 ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = x85 & n221 ;
  assign n1855 = n1853 | n1854 ;
  assign n1856 = ( ~x5 & n1849 ) | ( ~x5 & n1855 ) | ( n1849 & n1855 ) ;
  assign n1857 = x5 & ~n1855 ;
  assign n1858 = ( ~n1850 & n1856 ) | ( ~n1850 & n1857 ) | ( n1856 & n1857 ) ;
  assign n1859 = n649 & n697 ;
  assign n1860 = x14 & n1859 ;
  assign n1861 = x78 & n656 ;
  assign n1862 = x77 & n653 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = x76 & n744 ;
  assign n1865 = n1863 | n1864 ;
  assign n1866 = ( ~x14 & n1859 ) | ( ~x14 & n1865 ) | ( n1859 & n1865 ) ;
  assign n1867 = x14 & ~n1865 ;
  assign n1868 = ( ~n1860 & n1866 ) | ( ~n1860 & n1867 ) | ( n1866 & n1867 ) ;
  assign n1869 = n372 & n1146 ;
  assign n1870 = x20 & n1869 ;
  assign n1871 = x72 & n1153 ;
  assign n1872 = x71 & n1150 ;
  assign n1873 = n1871 | n1872 ;
  assign n1874 = x70 & n1217 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = ( ~x20 & n1869 ) | ( ~x20 & n1875 ) | ( n1869 & n1875 ) ;
  assign n1877 = x20 & ~n1875 ;
  assign n1878 = ( ~n1870 & n1876 ) | ( ~n1870 & n1877 ) | ( n1876 & n1877 ) ;
  assign n1879 = n240 & n1427 ;
  assign n1880 = x23 & n1879 ;
  assign n1881 = x69 & n1434 ;
  assign n1882 = x68 & n1431 ;
  assign n1883 = n1881 | n1882 ;
  assign n1884 = x67 & n1531 ;
  assign n1885 = n1883 | n1884 ;
  assign n1886 = ( ~x23 & n1879 ) | ( ~x23 & n1885 ) | ( n1879 & n1885 ) ;
  assign n1887 = x23 & ~n1885 ;
  assign n1888 = ( ~n1880 & n1886 ) | ( ~n1880 & n1887 ) | ( n1886 & n1887 ) ;
  assign n1889 = x65 & n1759 ;
  assign n1890 = n226 & n1755 ;
  assign n1891 = n1889 | n1890 ;
  assign n1892 = x66 & n1762 ;
  assign n1893 = n1891 | n1892 ;
  assign n1894 = ~n1654 & n1754 ;
  assign n1895 = ~n1759 & n1894 ;
  assign n1896 = x64 & n1895 ;
  assign n1897 = n1893 | n1896 ;
  assign n1898 = x26 & ~n1765 ;
  assign n1899 = ( x26 & ~n1897 ) | ( x26 & n1898 ) | ( ~n1897 & n1898 ) ;
  assign n1900 = ~n1897 & n1898 ;
  assign n1901 = ( x26 & n1897 ) | ( x26 & ~n1900 ) | ( n1897 & ~n1900 ) ;
  assign n1902 = ( ~x26 & n1899 ) | ( ~x26 & n1901 ) | ( n1899 & n1901 ) ;
  assign n1903 = ( n1770 & ~n1888 ) | ( n1770 & n1902 ) | ( ~n1888 & n1902 ) ;
  assign n1904 = ( n1770 & n1888 ) | ( n1770 & n1902 ) | ( n1888 & n1902 ) ;
  assign n1905 = ( n1888 & n1903 ) | ( n1888 & ~n1904 ) | ( n1903 & ~n1904 ) ;
  assign n1906 = ( n1783 & n1878 ) | ( n1783 & n1905 ) | ( n1878 & n1905 ) ;
  assign n1907 = ( ~n1783 & n1878 ) | ( ~n1783 & n1905 ) | ( n1878 & n1905 ) ;
  assign n1908 = ( n1783 & ~n1906 ) | ( n1783 & n1907 ) | ( ~n1906 & n1907 ) ;
  assign n1909 = n508 & n874 ;
  assign n1910 = x17 & n1909 ;
  assign n1911 = x75 & n881 ;
  assign n1912 = x74 & n878 ;
  assign n1913 = n1911 | n1912 ;
  assign n1914 = x73 & n959 ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = ( ~x17 & n1909 ) | ( ~x17 & n1915 ) | ( n1909 & n1915 ) ;
  assign n1917 = x17 & ~n1915 ;
  assign n1918 = ( ~n1910 & n1916 ) | ( ~n1910 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = ( n1785 & ~n1908 ) | ( n1785 & n1918 ) | ( ~n1908 & n1918 ) ;
  assign n1920 = ( n1785 & n1908 ) | ( n1785 & n1918 ) | ( n1908 & n1918 ) ;
  assign n1921 = ( n1908 & n1919 ) | ( n1908 & ~n1920 ) | ( n1919 & ~n1920 ) ;
  assign n1922 = ( n1799 & n1868 ) | ( n1799 & n1921 ) | ( n1868 & n1921 ) ;
  assign n1923 = ( ~n1799 & n1868 ) | ( ~n1799 & n1921 ) | ( n1868 & n1921 ) ;
  assign n1924 = ( n1799 & ~n1922 ) | ( n1799 & n1923 ) | ( ~n1922 & n1923 ) ;
  assign n1925 = n449 & n990 ;
  assign n1926 = x11 & n1925 ;
  assign n1927 = x80 & n453 ;
  assign n1928 = x79 & n536 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = x81 & n456 ;
  assign n1931 = n1929 | n1930 ;
  assign n1932 = ( ~x11 & n1925 ) | ( ~x11 & n1931 ) | ( n1925 & n1931 ) ;
  assign n1933 = x11 & ~n1931 ;
  assign n1934 = ( ~n1926 & n1932 ) | ( ~n1926 & n1933 ) | ( n1932 & n1933 ) ;
  assign n1935 = ( n1801 & n1924 ) | ( n1801 & n1934 ) | ( n1924 & n1934 ) ;
  assign n1936 = ( ~n1801 & n1924 ) | ( ~n1801 & n1934 ) | ( n1924 & n1934 ) ;
  assign n1937 = ( n1801 & ~n1935 ) | ( n1801 & n1936 ) | ( ~n1935 & n1936 ) ;
  assign n1938 = n301 & n1190 ;
  assign n1939 = x8 & n1938 ;
  assign n1940 = x84 & n309 ;
  assign n1941 = x83 & n306 ;
  assign n1942 = n1940 | n1941 ;
  assign n1943 = x82 & n359 ;
  assign n1944 = n1942 | n1943 ;
  assign n1945 = ( ~x8 & n1938 ) | ( ~x8 & n1944 ) | ( n1938 & n1944 ) ;
  assign n1946 = x8 & ~n1944 ;
  assign n1947 = ( ~n1939 & n1945 ) | ( ~n1939 & n1946 ) | ( n1945 & n1946 ) ;
  assign n1948 = ( ~n1815 & n1937 ) | ( ~n1815 & n1947 ) | ( n1937 & n1947 ) ;
  assign n1949 = ( n1815 & n1937 ) | ( n1815 & n1947 ) | ( n1937 & n1947 ) ;
  assign n1950 = ( n1815 & n1948 ) | ( n1815 & ~n1949 ) | ( n1948 & ~n1949 ) ;
  assign n1951 = ( n1818 & ~n1858 ) | ( n1818 & n1950 ) | ( ~n1858 & n1950 ) ;
  assign n1952 = ( n1818 & n1858 ) | ( n1818 & n1950 ) | ( n1858 & n1950 ) ;
  assign n1953 = ( n1858 & n1951 ) | ( n1858 & ~n1952 ) | ( n1951 & ~n1952 ) ;
  assign n1954 = ( n1834 & n1848 ) | ( n1834 & n1953 ) | ( n1848 & n1953 ) ;
  assign n1955 = ( ~n1834 & n1848 ) | ( ~n1834 & n1953 ) | ( n1848 & n1953 ) ;
  assign n1956 = ( n1834 & ~n1954 ) | ( n1834 & n1955 ) | ( ~n1954 & n1955 ) ;
  assign n1957 = ( ~x90 & x91 ) | ( ~x90 & n1837 ) | ( x91 & n1837 ) ;
  assign n1958 = ( x90 & x91 ) | ( x90 & n1837 ) | ( x91 & n1837 ) ;
  assign n1959 = ( x90 & n1957 ) | ( x90 & ~n1958 ) | ( n1957 & ~n1958 ) ;
  assign n1960 = x0 & n1959 ;
  assign n1961 = ( x1 & x2 ) | ( x1 & n1960 ) | ( x2 & n1960 ) ;
  assign n1962 = x90 & n172 ;
  assign n1963 = x91 | n1962 ;
  assign n1964 = ( n147 & n1962 ) | ( n147 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1965 = ( ~x89 & n135 ) | ( ~x89 & n174 ) | ( n135 & n174 ) ;
  assign n1966 = n1964 | n1965 ;
  assign n1967 = n1961 | n1966 ;
  assign n1968 = n1961 & n1966 ;
  assign n1969 = n1967 & ~n1968 ;
  assign n1970 = n301 & n1368 ;
  assign n1971 = x8 & n1970 ;
  assign n1972 = x85 & n309 ;
  assign n1973 = x84 & n306 ;
  assign n1974 = n1972 | n1973 ;
  assign n1975 = x83 & n359 ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = ( ~x8 & n1970 ) | ( ~x8 & n1976 ) | ( n1970 & n1976 ) ;
  assign n1978 = x8 & ~n1976 ;
  assign n1979 = ( ~n1971 & n1977 ) | ( ~n1971 & n1978 ) | ( n1977 & n1978 ) ;
  assign n1980 = n565 & n874 ;
  assign n1981 = x17 & n1980 ;
  assign n1982 = x76 & n881 ;
  assign n1983 = x75 & n878 ;
  assign n1984 = n1982 | n1983 ;
  assign n1985 = x74 & n959 ;
  assign n1986 = n1984 | n1985 ;
  assign n1987 = ( ~x17 & n1980 ) | ( ~x17 & n1986 ) | ( n1980 & n1986 ) ;
  assign n1988 = x17 & ~n1986 ;
  assign n1989 = ( ~n1981 & n1987 ) | ( ~n1981 & n1988 ) | ( n1987 & n1988 ) ;
  assign n1990 = n169 & n1755 ;
  assign n1991 = x26 & n1990 ;
  assign n1992 = x67 & n1762 ;
  assign n1993 = x66 & n1759 ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = x65 & n1895 ;
  assign n1996 = n1994 | n1995 ;
  assign n1997 = ( ~x26 & n1990 ) | ( ~x26 & n1996 ) | ( n1990 & n1996 ) ;
  assign n1998 = x26 & ~n1996 ;
  assign n1999 = ( ~n1991 & n1997 ) | ( ~n1991 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2000 = x26 | x27 ;
  assign n2001 = x26 & x27 ;
  assign n2002 = n2000 & ~n2001 ;
  assign n2003 = x64 & n2002 ;
  assign n2004 = ( ~n1900 & n1999 ) | ( ~n1900 & n2003 ) | ( n1999 & n2003 ) ;
  assign n2005 = ( n1900 & n1999 ) | ( n1900 & n2003 ) | ( n1999 & n2003 ) ;
  assign n2006 = ( n1900 & n2004 ) | ( n1900 & ~n2005 ) | ( n2004 & ~n2005 ) ;
  assign n2007 = n276 & n1427 ;
  assign n2008 = x23 & n2007 ;
  assign n2009 = x70 & n1434 ;
  assign n2010 = x69 & n1431 ;
  assign n2011 = n2009 | n2010 ;
  assign n2012 = x68 & n1531 ;
  assign n2013 = n2011 | n2012 ;
  assign n2014 = ( ~x23 & n2007 ) | ( ~x23 & n2013 ) | ( n2007 & n2013 ) ;
  assign n2015 = x23 & ~n2013 ;
  assign n2016 = ( ~n2008 & n2014 ) | ( ~n2008 & n2015 ) | ( n2014 & n2015 ) ;
  assign n2017 = ( n1904 & n2006 ) | ( n1904 & n2016 ) | ( n2006 & n2016 ) ;
  assign n2018 = ( ~n1904 & n2006 ) | ( ~n1904 & n2016 ) | ( n2006 & n2016 ) ;
  assign n2019 = ( n1904 & ~n2017 ) | ( n1904 & n2018 ) | ( ~n2017 & n2018 ) ;
  assign n2020 = n388 & n1146 ;
  assign n2021 = x20 & n2020 ;
  assign n2022 = x73 & n1153 ;
  assign n2023 = x72 & n1150 ;
  assign n2024 = n2022 | n2023 ;
  assign n2025 = x71 & n1217 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = ( ~x20 & n2020 ) | ( ~x20 & n2026 ) | ( n2020 & n2026 ) ;
  assign n2028 = x20 & ~n2026 ;
  assign n2029 = ( ~n2021 & n2027 ) | ( ~n2021 & n2028 ) | ( n2027 & n2028 ) ;
  assign n2030 = ( n1906 & ~n2019 ) | ( n1906 & n2029 ) | ( ~n2019 & n2029 ) ;
  assign n2031 = ( n1906 & n2019 ) | ( n1906 & n2029 ) | ( n2019 & n2029 ) ;
  assign n2032 = ( n2019 & n2030 ) | ( n2019 & ~n2031 ) | ( n2030 & ~n2031 ) ;
  assign n2033 = ( n1920 & n1989 ) | ( n1920 & n2032 ) | ( n1989 & n2032 ) ;
  assign n2034 = ( ~n1920 & n1989 ) | ( ~n1920 & n2032 ) | ( n1989 & n2032 ) ;
  assign n2035 = ( n1920 & ~n2033 ) | ( n1920 & n2034 ) | ( ~n2033 & n2034 ) ;
  assign n2036 = n649 & n823 ;
  assign n2037 = x14 & n2036 ;
  assign n2038 = x79 & n656 ;
  assign n2039 = x78 & n653 ;
  assign n2040 = n2038 | n2039 ;
  assign n2041 = x77 & n744 ;
  assign n2042 = n2040 | n2041 ;
  assign n2043 = ( ~x14 & n2036 ) | ( ~x14 & n2042 ) | ( n2036 & n2042 ) ;
  assign n2044 = x14 & ~n2042 ;
  assign n2045 = ( ~n2037 & n2043 ) | ( ~n2037 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2046 = ( n1922 & ~n2035 ) | ( n1922 & n2045 ) | ( ~n2035 & n2045 ) ;
  assign n2047 = ( n1922 & n2035 ) | ( n1922 & n2045 ) | ( n2035 & n2045 ) ;
  assign n2048 = ( n2035 & n2046 ) | ( n2035 & ~n2047 ) | ( n2046 & ~n2047 ) ;
  assign n2049 = n449 & n1006 ;
  assign n2050 = x11 & n2049 ;
  assign n2051 = x82 & n456 ;
  assign n2052 = x81 & n453 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = x80 & n536 ;
  assign n2055 = n2053 | n2054 ;
  assign n2056 = ( ~x11 & n2049 ) | ( ~x11 & n2055 ) | ( n2049 & n2055 ) ;
  assign n2057 = x11 & ~n2055 ;
  assign n2058 = ( ~n2050 & n2056 ) | ( ~n2050 & n2057 ) | ( n2056 & n2057 ) ;
  assign n2059 = ( n1935 & ~n2048 ) | ( n1935 & n2058 ) | ( ~n2048 & n2058 ) ;
  assign n2060 = ( n1935 & n2048 ) | ( n1935 & n2058 ) | ( n2048 & n2058 ) ;
  assign n2061 = ( n2048 & n2059 ) | ( n2048 & ~n2060 ) | ( n2059 & ~n2060 ) ;
  assign n2062 = ( n1949 & n1979 ) | ( n1949 & n2061 ) | ( n1979 & n2061 ) ;
  assign n2063 = ( ~n1949 & n1979 ) | ( ~n1949 & n2061 ) | ( n1979 & n2061 ) ;
  assign n2064 = ( n1949 & ~n2062 ) | ( n1949 & n2063 ) | ( ~n2062 & n2063 ) ;
  assign n2065 = n206 & n1602 ;
  assign n2066 = x5 & n2065 ;
  assign n2067 = x88 & n205 ;
  assign n2068 = x87 & n201 ;
  assign n2069 = n2067 | n2068 ;
  assign n2070 = x86 & n221 ;
  assign n2071 = n2069 | n2070 ;
  assign n2072 = ( ~x5 & n2065 ) | ( ~x5 & n2071 ) | ( n2065 & n2071 ) ;
  assign n2073 = x5 & ~n2071 ;
  assign n2074 = ( ~n2066 & n2072 ) | ( ~n2066 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2075 = ( n1952 & ~n2064 ) | ( n1952 & n2074 ) | ( ~n2064 & n2074 ) ;
  assign n2076 = ( n1952 & n2064 ) | ( n1952 & n2074 ) | ( n2064 & n2074 ) ;
  assign n2077 = ( n2064 & n2075 ) | ( n2064 & ~n2076 ) | ( n2075 & ~n2076 ) ;
  assign n2078 = ( n1954 & n1969 ) | ( n1954 & n2077 ) | ( n1969 & n2077 ) ;
  assign n2079 = ( ~n1954 & n1969 ) | ( ~n1954 & n2077 ) | ( n1969 & n2077 ) ;
  assign n2080 = ( n1954 & ~n2078 ) | ( n1954 & n2079 ) | ( ~n2078 & n2079 ) ;
  assign n2081 = ( ~x91 & x92 ) | ( ~x91 & n1958 ) | ( x92 & n1958 ) ;
  assign n2082 = ( x91 & x92 ) | ( x91 & n1958 ) | ( x92 & n1958 ) ;
  assign n2083 = ( x91 & n2081 ) | ( x91 & ~n2082 ) | ( n2081 & ~n2082 ) ;
  assign n2084 = x0 & n2083 ;
  assign n2085 = ( x1 & x2 ) | ( x1 & n2084 ) | ( x2 & n2084 ) ;
  assign n2086 = x91 & n172 ;
  assign n2087 = ( ~x90 & n135 ) | ( ~x90 & n174 ) | ( n135 & n174 ) ;
  assign n2088 = n2086 | n2087 ;
  assign n2089 = x92 & n147 ;
  assign n2090 = n2088 | n2089 ;
  assign n2091 = n2085 | n2090 ;
  assign n2092 = n2085 & n2090 ;
  assign n2093 = n2091 & ~n2092 ;
  assign n2094 = n206 & n1822 ;
  assign n2095 = x5 & n2094 ;
  assign n2096 = x89 & n205 ;
  assign n2097 = x88 & n201 ;
  assign n2098 = n2096 | n2097 ;
  assign n2099 = x87 & n221 ;
  assign n2100 = n2098 | n2099 ;
  assign n2101 = ( ~x5 & n2094 ) | ( ~x5 & n2100 ) | ( n2094 & n2100 ) ;
  assign n2102 = x5 & ~n2100 ;
  assign n2103 = ( ~n2095 & n2101 ) | ( ~n2095 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2104 = n649 & n840 ;
  assign n2105 = x14 & n2104 ;
  assign n2106 = x80 & n656 ;
  assign n2107 = x79 & n653 ;
  assign n2108 = n2106 | n2107 ;
  assign n2109 = x78 & n744 ;
  assign n2110 = n2108 | n2109 ;
  assign n2111 = ( ~x14 & n2104 ) | ( ~x14 & n2110 ) | ( n2104 & n2110 ) ;
  assign n2112 = x14 & ~n2110 ;
  assign n2113 = ( ~n2105 & n2111 ) | ( ~n2105 & n2112 ) | ( n2111 & n2112 ) ;
  assign n2114 = n626 & n874 ;
  assign n2115 = x17 & n2114 ;
  assign n2116 = x77 & n881 ;
  assign n2117 = x76 & n878 ;
  assign n2118 = n2116 | n2117 ;
  assign n2119 = x75 & n959 ;
  assign n2120 = n2118 | n2119 ;
  assign n2121 = ( ~x17 & n2114 ) | ( ~x17 & n2120 ) | ( n2114 & n2120 ) ;
  assign n2122 = x17 & ~n2120 ;
  assign n2123 = ( ~n2115 & n2121 ) | ( ~n2115 & n2122 ) | ( n2121 & n2122 ) ;
  assign n2124 = n1999 & n2005 ;
  assign n2125 = n193 & n1755 ;
  assign n2126 = x26 & n2125 ;
  assign n2127 = x68 & n1762 ;
  assign n2128 = x67 & n1759 ;
  assign n2129 = n2127 | n2128 ;
  assign n2130 = x66 & n1895 ;
  assign n2131 = n2129 | n2130 ;
  assign n2132 = ( ~x26 & n2125 ) | ( ~x26 & n2131 ) | ( n2125 & n2131 ) ;
  assign n2133 = x26 & ~n2131 ;
  assign n2134 = ( ~n2126 & n2132 ) | ( ~n2126 & n2133 ) | ( n2132 & n2133 ) ;
  assign n2135 = ~x28 & x29 ;
  assign n2136 = x28 & ~x29 ;
  assign n2137 = ( n2002 & n2135 ) | ( n2002 & n2136 ) | ( n2135 & n2136 ) ;
  assign n2138 = n302 & n2137 ;
  assign n2139 = ~x26 & x28 ;
  assign n2140 = x27 & x28 ;
  assign n2141 = ( n2001 & n2139 ) | ( n2001 & ~n2140 ) | ( n2139 & ~n2140 ) ;
  assign n2142 = x64 & n2141 ;
  assign n2143 = n2138 | n2142 ;
  assign n2144 = n2002 & ~n2137 ;
  assign n2145 = x65 & n2144 ;
  assign n2146 = n2143 | n2145 ;
  assign n2147 = n2003 | n2146 ;
  assign n2148 = ( x29 & n2003 ) | ( x29 & ~n2146 ) | ( n2003 & ~n2146 ) ;
  assign n2149 = x29 & ~n2146 ;
  assign n2150 = ( n2147 & ~n2148 ) | ( n2147 & n2149 ) | ( ~n2148 & n2149 ) ;
  assign n2151 = ( n2124 & n2134 ) | ( n2124 & n2150 ) | ( n2134 & n2150 ) ;
  assign n2152 = ( ~n2124 & n2134 ) | ( ~n2124 & n2150 ) | ( n2134 & n2150 ) ;
  assign n2153 = ( n2124 & ~n2151 ) | ( n2124 & n2152 ) | ( ~n2151 & n2152 ) ;
  assign n2154 = n322 & n1427 ;
  assign n2155 = x23 & n2154 ;
  assign n2156 = x71 & n1434 ;
  assign n2157 = x70 & n1431 ;
  assign n2158 = n2156 | n2157 ;
  assign n2159 = x69 & n1531 ;
  assign n2160 = n2158 | n2159 ;
  assign n2161 = ( ~x23 & n2154 ) | ( ~x23 & n2160 ) | ( n2154 & n2160 ) ;
  assign n2162 = x23 & ~n2160 ;
  assign n2163 = ( ~n2155 & n2161 ) | ( ~n2155 & n2162 ) | ( n2161 & n2162 ) ;
  assign n2164 = ( n2017 & n2153 ) | ( n2017 & n2163 ) | ( n2153 & n2163 ) ;
  assign n2165 = ( ~n2017 & n2153 ) | ( ~n2017 & n2163 ) | ( n2153 & n2163 ) ;
  assign n2166 = ( n2017 & ~n2164 ) | ( n2017 & n2165 ) | ( ~n2164 & n2165 ) ;
  assign n2167 = n436 & n1146 ;
  assign n2168 = x20 & n2167 ;
  assign n2169 = x74 & n1153 ;
  assign n2170 = x73 & n1150 ;
  assign n2171 = n2169 | n2170 ;
  assign n2172 = x72 & n1217 ;
  assign n2173 = n2171 | n2172 ;
  assign n2174 = ( ~x20 & n2167 ) | ( ~x20 & n2173 ) | ( n2167 & n2173 ) ;
  assign n2175 = x20 & ~n2173 ;
  assign n2176 = ( ~n2168 & n2174 ) | ( ~n2168 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2177 = ( n2031 & ~n2166 ) | ( n2031 & n2176 ) | ( ~n2166 & n2176 ) ;
  assign n2178 = ( n2031 & n2166 ) | ( n2031 & n2176 ) | ( n2166 & n2176 ) ;
  assign n2179 = ( n2166 & n2177 ) | ( n2166 & ~n2178 ) | ( n2177 & ~n2178 ) ;
  assign n2180 = ( n2033 & n2123 ) | ( n2033 & n2179 ) | ( n2123 & n2179 ) ;
  assign n2181 = ( ~n2033 & n2123 ) | ( ~n2033 & n2179 ) | ( n2123 & n2179 ) ;
  assign n2182 = ( n2033 & ~n2180 ) | ( n2033 & n2181 ) | ( ~n2180 & n2181 ) ;
  assign n2183 = ( n2047 & n2113 ) | ( n2047 & n2182 ) | ( n2113 & n2182 ) ;
  assign n2184 = ( ~n2047 & n2113 ) | ( ~n2047 & n2182 ) | ( n2113 & n2182 ) ;
  assign n2185 = ( n2047 & ~n2183 ) | ( n2047 & n2184 ) | ( ~n2183 & n2184 ) ;
  assign n2186 = n449 & n1093 ;
  assign n2187 = x11 & n2186 ;
  assign n2188 = x83 & n456 ;
  assign n2189 = x82 & n453 ;
  assign n2190 = n2188 | n2189 ;
  assign n2191 = x81 & n536 ;
  assign n2192 = n2190 | n2191 ;
  assign n2193 = ( ~x11 & n2186 ) | ( ~x11 & n2192 ) | ( n2186 & n2192 ) ;
  assign n2194 = x11 & ~n2192 ;
  assign n2195 = ( ~n2187 & n2193 ) | ( ~n2187 & n2194 ) | ( n2193 & n2194 ) ;
  assign n2196 = ( n2060 & n2185 ) | ( n2060 & n2195 ) | ( n2185 & n2195 ) ;
  assign n2197 = ( ~n2060 & n2185 ) | ( ~n2060 & n2195 ) | ( n2185 & n2195 ) ;
  assign n2198 = ( n2060 & ~n2196 ) | ( n2060 & n2197 ) | ( ~n2196 & n2197 ) ;
  assign n2199 = n301 & n1384 ;
  assign n2200 = x8 & n2199 ;
  assign n2201 = x86 & n309 ;
  assign n2202 = x85 & n306 ;
  assign n2203 = n2201 | n2202 ;
  assign n2204 = x84 & n359 ;
  assign n2205 = n2203 | n2204 ;
  assign n2206 = ( ~x8 & n2199 ) | ( ~x8 & n2205 ) | ( n2199 & n2205 ) ;
  assign n2207 = x8 & ~n2205 ;
  assign n2208 = ( ~n2200 & n2206 ) | ( ~n2200 & n2207 ) | ( n2206 & n2207 ) ;
  assign n2209 = ( ~n2062 & n2198 ) | ( ~n2062 & n2208 ) | ( n2198 & n2208 ) ;
  assign n2210 = ( n2062 & n2198 ) | ( n2062 & n2208 ) | ( n2198 & n2208 ) ;
  assign n2211 = ( n2062 & n2209 ) | ( n2062 & ~n2210 ) | ( n2209 & ~n2210 ) ;
  assign n2212 = ( n2076 & ~n2103 ) | ( n2076 & n2211 ) | ( ~n2103 & n2211 ) ;
  assign n2213 = ( n2076 & n2103 ) | ( n2076 & n2211 ) | ( n2103 & n2211 ) ;
  assign n2214 = ( n2103 & n2212 ) | ( n2103 & ~n2213 ) | ( n2212 & ~n2213 ) ;
  assign n2215 = ( n2078 & n2093 ) | ( n2078 & n2214 ) | ( n2093 & n2214 ) ;
  assign n2216 = ( ~n2078 & n2093 ) | ( ~n2078 & n2214 ) | ( n2093 & n2214 ) ;
  assign n2217 = ( n2078 & ~n2215 ) | ( n2078 & n2216 ) | ( ~n2215 & n2216 ) ;
  assign n2218 = ( ~x92 & x93 ) | ( ~x92 & n2082 ) | ( x93 & n2082 ) ;
  assign n2219 = ( x92 & x93 ) | ( x92 & n2082 ) | ( x93 & n2082 ) ;
  assign n2220 = ( x92 & n2218 ) | ( x92 & ~n2219 ) | ( n2218 & ~n2219 ) ;
  assign n2221 = x0 & n2220 ;
  assign n2222 = ( x1 & x2 ) | ( x1 & n2221 ) | ( x2 & n2221 ) ;
  assign n2223 = x92 & n172 ;
  assign n2224 = ( ~x91 & n135 ) | ( ~x91 & n174 ) | ( n135 & n174 ) ;
  assign n2225 = n2223 | n2224 ;
  assign n2226 = x93 & n147 ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = n2222 | n2227 ;
  assign n2229 = n2222 & n2227 ;
  assign n2230 = n2228 & ~n2229 ;
  assign n2231 = n206 & n1838 ;
  assign n2232 = x5 & n2231 ;
  assign n2233 = x90 & n205 ;
  assign n2234 = x89 & n201 ;
  assign n2235 = n2233 | n2234 ;
  assign n2236 = x88 & n221 ;
  assign n2237 = n2235 | n2236 ;
  assign n2238 = ( ~x5 & n2231 ) | ( ~x5 & n2237 ) | ( n2231 & n2237 ) ;
  assign n2239 = x5 & ~n2237 ;
  assign n2240 = ( ~n2232 & n2238 ) | ( ~n2232 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2241 = n301 & n1494 ;
  assign n2242 = x8 & n2241 ;
  assign n2243 = x87 & n309 ;
  assign n2244 = x86 & n306 ;
  assign n2245 = n2243 | n2244 ;
  assign n2246 = x85 & n359 ;
  assign n2247 = n2245 | n2246 ;
  assign n2248 = ( ~x8 & n2241 ) | ( ~x8 & n2247 ) | ( n2241 & n2247 ) ;
  assign n2249 = x8 & ~n2247 ;
  assign n2250 = ( ~n2242 & n2248 ) | ( ~n2242 & n2249 ) | ( n2248 & n2249 ) ;
  assign n2251 = n508 & n1146 ;
  assign n2252 = x20 & n2251 ;
  assign n2253 = x75 & n1153 ;
  assign n2254 = x74 & n1150 ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = x73 & n1217 ;
  assign n2257 = n2255 | n2256 ;
  assign n2258 = ( ~x20 & n2251 ) | ( ~x20 & n2257 ) | ( n2251 & n2257 ) ;
  assign n2259 = x20 & ~n2257 ;
  assign n2260 = ( ~n2252 & n2258 ) | ( ~n2252 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2261 = x66 & n2144 ;
  assign n2262 = x65 & n2141 ;
  assign n2263 = n2261 | n2262 ;
  assign n2264 = n226 & n2137 ;
  assign n2265 = n2001 & n2136 ;
  assign n2266 = ~n2000 & n2135 ;
  assign n2267 = n2265 | n2266 ;
  assign n2268 = x64 & ~n2267 ;
  assign n2269 = ( x64 & n2264 ) | ( x64 & ~n2268 ) | ( n2264 & ~n2268 ) ;
  assign n2270 = n2263 | n2269 ;
  assign n2271 = ~x29 & n2270 ;
  assign n2272 = ( x29 & n2147 ) | ( x29 & n2270 ) | ( n2147 & n2270 ) ;
  assign n2273 = n2147 & n2270 ;
  assign n2274 = ( n2271 & n2272 ) | ( n2271 & ~n2273 ) | ( n2272 & ~n2273 ) ;
  assign n2275 = n240 & n1755 ;
  assign n2276 = x26 & n2275 ;
  assign n2277 = x69 & n1762 ;
  assign n2278 = x68 & n1759 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = x67 & n1895 ;
  assign n2281 = n2279 | n2280 ;
  assign n2282 = ( ~x26 & n2275 ) | ( ~x26 & n2281 ) | ( n2275 & n2281 ) ;
  assign n2283 = x26 & ~n2281 ;
  assign n2284 = ( ~n2276 & n2282 ) | ( ~n2276 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2285 = ( n2151 & n2274 ) | ( n2151 & n2284 ) | ( n2274 & n2284 ) ;
  assign n2286 = ( ~n2151 & n2274 ) | ( ~n2151 & n2284 ) | ( n2274 & n2284 ) ;
  assign n2287 = ( n2151 & ~n2285 ) | ( n2151 & n2286 ) | ( ~n2285 & n2286 ) ;
  assign n2288 = n372 & n1427 ;
  assign n2289 = x23 & n2288 ;
  assign n2290 = x72 & n1434 ;
  assign n2291 = x71 & n1431 ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = x70 & n1531 ;
  assign n2294 = n2292 | n2293 ;
  assign n2295 = ( ~x23 & n2288 ) | ( ~x23 & n2294 ) | ( n2288 & n2294 ) ;
  assign n2296 = x23 & ~n2294 ;
  assign n2297 = ( ~n2289 & n2295 ) | ( ~n2289 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = ( n2164 & ~n2287 ) | ( n2164 & n2297 ) | ( ~n2287 & n2297 ) ;
  assign n2299 = ( n2164 & n2287 ) | ( n2164 & n2297 ) | ( n2287 & n2297 ) ;
  assign n2300 = ( n2287 & n2298 ) | ( n2287 & ~n2299 ) | ( n2298 & ~n2299 ) ;
  assign n2301 = ( n2178 & n2260 ) | ( n2178 & n2300 ) | ( n2260 & n2300 ) ;
  assign n2302 = ( ~n2178 & n2260 ) | ( ~n2178 & n2300 ) | ( n2260 & n2300 ) ;
  assign n2303 = ( n2178 & ~n2301 ) | ( n2178 & n2302 ) | ( ~n2301 & n2302 ) ;
  assign n2304 = n697 & n874 ;
  assign n2305 = x17 & n2304 ;
  assign n2306 = x78 & n881 ;
  assign n2307 = x77 & n878 ;
  assign n2308 = n2306 | n2307 ;
  assign n2309 = x76 & n959 ;
  assign n2310 = n2308 | n2309 ;
  assign n2311 = ( ~x17 & n2304 ) | ( ~x17 & n2310 ) | ( n2304 & n2310 ) ;
  assign n2312 = x17 & ~n2310 ;
  assign n2313 = ( ~n2305 & n2311 ) | ( ~n2305 & n2312 ) | ( n2311 & n2312 ) ;
  assign n2314 = ( n2180 & n2303 ) | ( n2180 & n2313 ) | ( n2303 & n2313 ) ;
  assign n2315 = ( ~n2180 & n2303 ) | ( ~n2180 & n2313 ) | ( n2303 & n2313 ) ;
  assign n2316 = ( n2180 & ~n2314 ) | ( n2180 & n2315 ) | ( ~n2314 & n2315 ) ;
  assign n2317 = n649 & n990 ;
  assign n2318 = x14 & n2317 ;
  assign n2319 = x81 & n656 ;
  assign n2320 = x80 & n653 ;
  assign n2321 = n2319 | n2320 ;
  assign n2322 = x79 & n744 ;
  assign n2323 = n2321 | n2322 ;
  assign n2324 = ( ~x14 & n2317 ) | ( ~x14 & n2323 ) | ( n2317 & n2323 ) ;
  assign n2325 = x14 & ~n2323 ;
  assign n2326 = ( ~n2318 & n2324 ) | ( ~n2318 & n2325 ) | ( n2324 & n2325 ) ;
  assign n2327 = ( n2183 & ~n2316 ) | ( n2183 & n2326 ) | ( ~n2316 & n2326 ) ;
  assign n2328 = ( n2183 & n2316 ) | ( n2183 & n2326 ) | ( n2316 & n2326 ) ;
  assign n2329 = ( n2316 & n2327 ) | ( n2316 & ~n2328 ) | ( n2327 & ~n2328 ) ;
  assign n2330 = n449 & n1190 ;
  assign n2331 = x11 & n2330 ;
  assign n2332 = x84 & n456 ;
  assign n2333 = x83 & n453 ;
  assign n2334 = n2332 | n2333 ;
  assign n2335 = x82 & n536 ;
  assign n2336 = n2334 | n2335 ;
  assign n2337 = ( ~x11 & n2330 ) | ( ~x11 & n2336 ) | ( n2330 & n2336 ) ;
  assign n2338 = x11 & ~n2336 ;
  assign n2339 = ( ~n2331 & n2337 ) | ( ~n2331 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2340 = ( n2196 & ~n2329 ) | ( n2196 & n2339 ) | ( ~n2329 & n2339 ) ;
  assign n2341 = ( n2196 & n2329 ) | ( n2196 & n2339 ) | ( n2329 & n2339 ) ;
  assign n2342 = ( n2329 & n2340 ) | ( n2329 & ~n2341 ) | ( n2340 & ~n2341 ) ;
  assign n2343 = ( n2210 & n2250 ) | ( n2210 & n2342 ) | ( n2250 & n2342 ) ;
  assign n2344 = ( ~n2210 & n2250 ) | ( ~n2210 & n2342 ) | ( n2250 & n2342 ) ;
  assign n2345 = ( n2210 & ~n2343 ) | ( n2210 & n2344 ) | ( ~n2343 & n2344 ) ;
  assign n2346 = ( n2213 & ~n2240 ) | ( n2213 & n2345 ) | ( ~n2240 & n2345 ) ;
  assign n2347 = ( n2213 & n2240 ) | ( n2213 & n2345 ) | ( n2240 & n2345 ) ;
  assign n2348 = ( n2240 & n2346 ) | ( n2240 & ~n2347 ) | ( n2346 & ~n2347 ) ;
  assign n2349 = ( n2215 & n2230 ) | ( n2215 & n2348 ) | ( n2230 & n2348 ) ;
  assign n2350 = ( n2215 & ~n2230 ) | ( n2215 & n2348 ) | ( ~n2230 & n2348 ) ;
  assign n2351 = ( n2230 & ~n2349 ) | ( n2230 & n2350 ) | ( ~n2349 & n2350 ) ;
  assign n2352 = n206 & n1959 ;
  assign n2353 = x5 & n2352 ;
  assign n2354 = x91 & n205 ;
  assign n2355 = x90 & n201 ;
  assign n2356 = n2354 | n2355 ;
  assign n2357 = x89 & n221 ;
  assign n2358 = n2356 | n2357 ;
  assign n2359 = ( ~x5 & n2352 ) | ( ~x5 & n2358 ) | ( n2352 & n2358 ) ;
  assign n2360 = x5 & ~n2358 ;
  assign n2361 = ( ~n2353 & n2359 ) | ( ~n2353 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2362 = n301 & n1602 ;
  assign n2363 = x8 & n2362 ;
  assign n2364 = x88 & n309 ;
  assign n2365 = x87 & n306 ;
  assign n2366 = n2364 | n2365 ;
  assign n2367 = x86 & n359 ;
  assign n2368 = n2366 | n2367 ;
  assign n2369 = ( ~x8 & n2362 ) | ( ~x8 & n2368 ) | ( n2362 & n2368 ) ;
  assign n2370 = x8 & ~n2368 ;
  assign n2371 = ( ~n2363 & n2369 ) | ( ~n2363 & n2370 ) | ( n2369 & n2370 ) ;
  assign n2372 = n276 & n1755 ;
  assign n2373 = x26 & n2372 ;
  assign n2374 = x70 & n1762 ;
  assign n2375 = x69 & n1759 ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = x68 & n1895 ;
  assign n2378 = n2376 | n2377 ;
  assign n2379 = ( ~x26 & n2372 ) | ( ~x26 & n2378 ) | ( n2372 & n2378 ) ;
  assign n2380 = x26 & ~n2378 ;
  assign n2381 = ( ~n2373 & n2379 ) | ( ~n2373 & n2380 ) | ( n2379 & n2380 ) ;
  assign n2382 = n2147 | n2270 ;
  assign n2383 = x29 & n2382 ;
  assign n2384 = x66 & n2141 ;
  assign n2385 = n169 & n2137 ;
  assign n2386 = x67 & n2144 ;
  assign n2387 = x65 & ~n2267 ;
  assign n2388 = ( x65 & n2386 ) | ( x65 & ~n2387 ) | ( n2386 & ~n2387 ) ;
  assign n2389 = n2385 | n2388 ;
  assign n2390 = n2384 | n2389 ;
  assign n2391 = x29 | x30 ;
  assign n2392 = x29 & x30 ;
  assign n2393 = n2391 & ~n2392 ;
  assign n2394 = x64 & n2393 ;
  assign n2395 = ( n2383 & ~n2390 ) | ( n2383 & n2394 ) | ( ~n2390 & n2394 ) ;
  assign n2396 = x29 & ~n2390 ;
  assign n2397 = ( ~n2383 & n2390 ) | ( ~n2383 & n2396 ) | ( n2390 & n2396 ) ;
  assign n2398 = ( n2394 & n2396 ) | ( n2394 & n2397 ) | ( n2396 & n2397 ) ;
  assign n2399 = ( n2395 & n2397 ) | ( n2395 & ~n2398 ) | ( n2397 & ~n2398 ) ;
  assign n2400 = ( n2285 & n2381 ) | ( n2285 & n2399 ) | ( n2381 & n2399 ) ;
  assign n2401 = ( ~n2285 & n2381 ) | ( ~n2285 & n2399 ) | ( n2381 & n2399 ) ;
  assign n2402 = ( n2285 & ~n2400 ) | ( n2285 & n2401 ) | ( ~n2400 & n2401 ) ;
  assign n2403 = n388 & n1427 ;
  assign n2404 = x23 & n2403 ;
  assign n2405 = x73 & n1434 ;
  assign n2406 = x72 & n1431 ;
  assign n2407 = n2405 | n2406 ;
  assign n2408 = x71 & n1531 ;
  assign n2409 = n2407 | n2408 ;
  assign n2410 = ( ~x23 & n2403 ) | ( ~x23 & n2409 ) | ( n2403 & n2409 ) ;
  assign n2411 = x23 & ~n2409 ;
  assign n2412 = ( ~n2404 & n2410 ) | ( ~n2404 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = ( ~n2299 & n2402 ) | ( ~n2299 & n2412 ) | ( n2402 & n2412 ) ;
  assign n2414 = ( n2299 & n2402 ) | ( n2299 & n2412 ) | ( n2402 & n2412 ) ;
  assign n2415 = ( n2299 & n2413 ) | ( n2299 & ~n2414 ) | ( n2413 & ~n2414 ) ;
  assign n2416 = n565 & n1146 ;
  assign n2417 = x20 & n2416 ;
  assign n2418 = x76 & n1153 ;
  assign n2419 = x75 & n1150 ;
  assign n2420 = n2418 | n2419 ;
  assign n2421 = x74 & n1217 ;
  assign n2422 = n2420 | n2421 ;
  assign n2423 = ( ~x20 & n2416 ) | ( ~x20 & n2422 ) | ( n2416 & n2422 ) ;
  assign n2424 = x20 & ~n2422 ;
  assign n2425 = ( ~n2417 & n2423 ) | ( ~n2417 & n2424 ) | ( n2423 & n2424 ) ;
  assign n2426 = ( ~n2301 & n2415 ) | ( ~n2301 & n2425 ) | ( n2415 & n2425 ) ;
  assign n2427 = ( n2301 & n2415 ) | ( n2301 & n2425 ) | ( n2415 & n2425 ) ;
  assign n2428 = ( n2301 & n2426 ) | ( n2301 & ~n2427 ) | ( n2426 & ~n2427 ) ;
  assign n2429 = n823 & n874 ;
  assign n2430 = x17 & n2429 ;
  assign n2431 = x79 & n881 ;
  assign n2432 = x78 & n878 ;
  assign n2433 = n2431 | n2432 ;
  assign n2434 = x77 & n959 ;
  assign n2435 = n2433 | n2434 ;
  assign n2436 = ( ~x17 & n2429 ) | ( ~x17 & n2435 ) | ( n2429 & n2435 ) ;
  assign n2437 = x17 & ~n2435 ;
  assign n2438 = ( ~n2430 & n2436 ) | ( ~n2430 & n2437 ) | ( n2436 & n2437 ) ;
  assign n2439 = ( n2314 & n2428 ) | ( n2314 & n2438 ) | ( n2428 & n2438 ) ;
  assign n2440 = ( ~n2314 & n2428 ) | ( ~n2314 & n2438 ) | ( n2428 & n2438 ) ;
  assign n2441 = ( n2314 & ~n2439 ) | ( n2314 & n2440 ) | ( ~n2439 & n2440 ) ;
  assign n2442 = n649 & n1006 ;
  assign n2443 = x14 & n2442 ;
  assign n2444 = x82 & n656 ;
  assign n2445 = x81 & n653 ;
  assign n2446 = n2444 | n2445 ;
  assign n2447 = x80 & n744 ;
  assign n2448 = n2446 | n2447 ;
  assign n2449 = ( ~x14 & n2442 ) | ( ~x14 & n2448 ) | ( n2442 & n2448 ) ;
  assign n2450 = x14 & ~n2448 ;
  assign n2451 = ( ~n2443 & n2449 ) | ( ~n2443 & n2450 ) | ( n2449 & n2450 ) ;
  assign n2452 = ( n2328 & ~n2441 ) | ( n2328 & n2451 ) | ( ~n2441 & n2451 ) ;
  assign n2453 = ( n2328 & n2441 ) | ( n2328 & n2451 ) | ( n2441 & n2451 ) ;
  assign n2454 = ( n2441 & n2452 ) | ( n2441 & ~n2453 ) | ( n2452 & ~n2453 ) ;
  assign n2455 = n449 & n1368 ;
  assign n2456 = x11 & n2455 ;
  assign n2457 = x85 & n456 ;
  assign n2458 = x84 & n453 ;
  assign n2459 = n2457 | n2458 ;
  assign n2460 = x83 & n536 ;
  assign n2461 = n2459 | n2460 ;
  assign n2462 = ( ~x11 & n2455 ) | ( ~x11 & n2461 ) | ( n2455 & n2461 ) ;
  assign n2463 = x11 & ~n2461 ;
  assign n2464 = ( ~n2456 & n2462 ) | ( ~n2456 & n2463 ) | ( n2462 & n2463 ) ;
  assign n2465 = ( n2341 & ~n2454 ) | ( n2341 & n2464 ) | ( ~n2454 & n2464 ) ;
  assign n2466 = ( n2341 & n2454 ) | ( n2341 & n2464 ) | ( n2454 & n2464 ) ;
  assign n2467 = ( n2454 & n2465 ) | ( n2454 & ~n2466 ) | ( n2465 & ~n2466 ) ;
  assign n2468 = ( n2343 & n2371 ) | ( n2343 & n2467 ) | ( n2371 & n2467 ) ;
  assign n2469 = ( ~n2343 & n2371 ) | ( ~n2343 & n2467 ) | ( n2371 & n2467 ) ;
  assign n2470 = ( n2343 & ~n2468 ) | ( n2343 & n2469 ) | ( ~n2468 & n2469 ) ;
  assign n2471 = ( n2347 & n2361 ) | ( n2347 & n2470 ) | ( n2361 & n2470 ) ;
  assign n2472 = ( ~n2347 & n2361 ) | ( ~n2347 & n2470 ) | ( n2361 & n2470 ) ;
  assign n2473 = ( n2347 & ~n2471 ) | ( n2347 & n2472 ) | ( ~n2471 & n2472 ) ;
  assign n2474 = ( ~x93 & x94 ) | ( ~x93 & n2219 ) | ( x94 & n2219 ) ;
  assign n2475 = ( x93 & x94 ) | ( x93 & n2219 ) | ( x94 & n2219 ) ;
  assign n2476 = ( x93 & n2474 ) | ( x93 & ~n2475 ) | ( n2474 & ~n2475 ) ;
  assign n2477 = x0 & n2476 ;
  assign n2478 = ( x1 & x2 ) | ( x1 & n2477 ) | ( x2 & n2477 ) ;
  assign n2479 = x93 & n172 ;
  assign n2480 = ( ~x92 & n135 ) | ( ~x92 & n174 ) | ( n135 & n174 ) ;
  assign n2481 = n2479 | n2480 ;
  assign n2482 = x94 & n147 ;
  assign n2483 = n2481 | n2482 ;
  assign n2484 = n2478 | n2483 ;
  assign n2485 = n2478 & n2483 ;
  assign n2486 = n2484 & ~n2485 ;
  assign n2487 = ( n2349 & ~n2473 ) | ( n2349 & n2486 ) | ( ~n2473 & n2486 ) ;
  assign n2488 = ( n2349 & n2473 ) | ( n2349 & n2486 ) | ( n2473 & n2486 ) ;
  assign n2489 = ( n2473 & n2487 ) | ( n2473 & ~n2488 ) | ( n2487 & ~n2488 ) ;
  assign n2490 = ( ~x94 & x95 ) | ( ~x94 & n2475 ) | ( x95 & n2475 ) ;
  assign n2491 = ( x94 & x95 ) | ( x94 & n2475 ) | ( x95 & n2475 ) ;
  assign n2492 = ( x94 & n2490 ) | ( x94 & ~n2491 ) | ( n2490 & ~n2491 ) ;
  assign n2493 = x0 & n2492 ;
  assign n2494 = ( x1 & x2 ) | ( x1 & n2493 ) | ( x2 & n2493 ) ;
  assign n2495 = x94 & n172 ;
  assign n2496 = x95 | n2495 ;
  assign n2497 = ( n147 & n2495 ) | ( n147 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2498 = ( ~x93 & n135 ) | ( ~x93 & n174 ) | ( n135 & n174 ) ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = n2494 | n2499 ;
  assign n2501 = n2494 & n2499 ;
  assign n2502 = n2500 & ~n2501 ;
  assign n2503 = n301 & n1822 ;
  assign n2504 = x8 & n2503 ;
  assign n2505 = x89 & n309 ;
  assign n2506 = x88 & n306 ;
  assign n2507 = n2505 | n2506 ;
  assign n2508 = x87 & n359 ;
  assign n2509 = n2507 | n2508 ;
  assign n2510 = ( ~x8 & n2503 ) | ( ~x8 & n2509 ) | ( n2503 & n2509 ) ;
  assign n2511 = x8 & ~n2509 ;
  assign n2512 = ( ~n2504 & n2510 ) | ( ~n2504 & n2511 ) | ( n2510 & n2511 ) ;
  assign n2513 = n649 & n1093 ;
  assign n2514 = x14 & n2513 ;
  assign n2515 = x83 & n656 ;
  assign n2516 = x82 & n653 ;
  assign n2517 = n2515 | n2516 ;
  assign n2518 = x81 & n744 ;
  assign n2519 = n2517 | n2518 ;
  assign n2520 = ( ~x14 & n2513 ) | ( ~x14 & n2519 ) | ( n2513 & n2519 ) ;
  assign n2521 = x14 & ~n2519 ;
  assign n2522 = ( ~n2514 & n2520 ) | ( ~n2514 & n2521 ) | ( n2520 & n2521 ) ;
  assign n2523 = n626 & n1146 ;
  assign n2524 = x20 & n2523 ;
  assign n2525 = x77 & n1153 ;
  assign n2526 = x76 & n1150 ;
  assign n2527 = n2525 | n2526 ;
  assign n2528 = x75 & n1217 ;
  assign n2529 = n2527 | n2528 ;
  assign n2530 = ( ~x20 & n2523 ) | ( ~x20 & n2529 ) | ( n2523 & n2529 ) ;
  assign n2531 = x20 & ~n2529 ;
  assign n2532 = ( ~n2524 & n2530 ) | ( ~n2524 & n2531 ) | ( n2530 & n2531 ) ;
  assign n2533 = n322 & n1755 ;
  assign n2534 = x26 & n2533 ;
  assign n2535 = x71 & n1762 ;
  assign n2536 = x70 & n1759 ;
  assign n2537 = n2535 | n2536 ;
  assign n2538 = x69 & n1895 ;
  assign n2539 = n2537 | n2538 ;
  assign n2540 = ( ~x26 & n2533 ) | ( ~x26 & n2539 ) | ( n2533 & n2539 ) ;
  assign n2541 = x26 & ~n2539 ;
  assign n2542 = ( ~n2534 & n2540 ) | ( ~n2534 & n2541 ) | ( n2540 & n2541 ) ;
  assign n2543 = ~x31 & x32 ;
  assign n2544 = x31 & ~x32 ;
  assign n2545 = ( n2393 & n2543 ) | ( n2393 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2546 = n302 & n2545 ;
  assign n2547 = ~x29 & x31 ;
  assign n2548 = x30 & x31 ;
  assign n2549 = ( n2392 & n2547 ) | ( n2392 & ~n2548 ) | ( n2547 & ~n2548 ) ;
  assign n2550 = x64 & n2549 ;
  assign n2551 = n2546 | n2550 ;
  assign n2552 = n2393 & ~n2545 ;
  assign n2553 = x65 & n2552 ;
  assign n2554 = n2551 | n2553 ;
  assign n2555 = n2394 | n2554 ;
  assign n2556 = ( x32 & n2394 ) | ( x32 & ~n2554 ) | ( n2394 & ~n2554 ) ;
  assign n2557 = x32 & ~n2554 ;
  assign n2558 = ( n2555 & ~n2556 ) | ( n2555 & n2557 ) | ( ~n2556 & n2557 ) ;
  assign n2559 = x68 & n2144 ;
  assign n2560 = x29 & n2559 ;
  assign n2561 = x67 & n2141 ;
  assign n2562 = x66 & n2267 ;
  assign n2563 = n2561 | n2562 ;
  assign n2564 = n193 & n2137 ;
  assign n2565 = n2563 | n2564 ;
  assign n2566 = ( ~x29 & n2559 ) | ( ~x29 & n2565 ) | ( n2559 & n2565 ) ;
  assign n2567 = x29 & ~n2565 ;
  assign n2568 = ( ~n2560 & n2566 ) | ( ~n2560 & n2567 ) | ( n2566 & n2567 ) ;
  assign n2569 = ( n2398 & ~n2558 ) | ( n2398 & n2568 ) | ( ~n2558 & n2568 ) ;
  assign n2570 = ( n2398 & n2558 ) | ( n2398 & n2568 ) | ( n2558 & n2568 ) ;
  assign n2571 = ( n2558 & n2569 ) | ( n2558 & ~n2570 ) | ( n2569 & ~n2570 ) ;
  assign n2572 = ( ~n2400 & n2542 ) | ( ~n2400 & n2571 ) | ( n2542 & n2571 ) ;
  assign n2573 = ( n2400 & n2542 ) | ( n2400 & n2571 ) | ( n2542 & n2571 ) ;
  assign n2574 = ( n2400 & n2572 ) | ( n2400 & ~n2573 ) | ( n2572 & ~n2573 ) ;
  assign n2575 = n436 & n1427 ;
  assign n2576 = x23 & n2575 ;
  assign n2577 = x74 & n1434 ;
  assign n2578 = x73 & n1431 ;
  assign n2579 = n2577 | n2578 ;
  assign n2580 = x72 & n1531 ;
  assign n2581 = n2579 | n2580 ;
  assign n2582 = ( ~x23 & n2575 ) | ( ~x23 & n2581 ) | ( n2575 & n2581 ) ;
  assign n2583 = x23 & ~n2581 ;
  assign n2584 = ( ~n2576 & n2582 ) | ( ~n2576 & n2583 ) | ( n2582 & n2583 ) ;
  assign n2585 = ( n2414 & ~n2574 ) | ( n2414 & n2584 ) | ( ~n2574 & n2584 ) ;
  assign n2586 = ( n2414 & n2574 ) | ( n2414 & n2584 ) | ( n2574 & n2584 ) ;
  assign n2587 = ( n2574 & n2585 ) | ( n2574 & ~n2586 ) | ( n2585 & ~n2586 ) ;
  assign n2588 = ( n2427 & n2532 ) | ( n2427 & n2587 ) | ( n2532 & n2587 ) ;
  assign n2589 = ( ~n2427 & n2532 ) | ( ~n2427 & n2587 ) | ( n2532 & n2587 ) ;
  assign n2590 = ( n2427 & ~n2588 ) | ( n2427 & n2589 ) | ( ~n2588 & n2589 ) ;
  assign n2591 = n840 & n874 ;
  assign n2592 = x17 & n2591 ;
  assign n2593 = x80 & n881 ;
  assign n2594 = x79 & n878 ;
  assign n2595 = n2593 | n2594 ;
  assign n2596 = x78 & n959 ;
  assign n2597 = n2595 | n2596 ;
  assign n2598 = ( ~x17 & n2591 ) | ( ~x17 & n2597 ) | ( n2591 & n2597 ) ;
  assign n2599 = x17 & ~n2597 ;
  assign n2600 = ( ~n2592 & n2598 ) | ( ~n2592 & n2599 ) | ( n2598 & n2599 ) ;
  assign n2601 = ( n2439 & ~n2590 ) | ( n2439 & n2600 ) | ( ~n2590 & n2600 ) ;
  assign n2602 = ( n2439 & n2590 ) | ( n2439 & n2600 ) | ( n2590 & n2600 ) ;
  assign n2603 = ( n2590 & n2601 ) | ( n2590 & ~n2602 ) | ( n2601 & ~n2602 ) ;
  assign n2604 = ( n2453 & n2522 ) | ( n2453 & n2603 ) | ( n2522 & n2603 ) ;
  assign n2605 = ( ~n2453 & n2522 ) | ( ~n2453 & n2603 ) | ( n2522 & n2603 ) ;
  assign n2606 = ( n2453 & ~n2604 ) | ( n2453 & n2605 ) | ( ~n2604 & n2605 ) ;
  assign n2607 = n449 & n1384 ;
  assign n2608 = x11 & n2607 ;
  assign n2609 = x86 & n456 ;
  assign n2610 = x85 & n453 ;
  assign n2611 = n2609 | n2610 ;
  assign n2612 = x84 & n536 ;
  assign n2613 = n2611 | n2612 ;
  assign n2614 = ( ~x11 & n2607 ) | ( ~x11 & n2613 ) | ( n2607 & n2613 ) ;
  assign n2615 = x11 & ~n2613 ;
  assign n2616 = ( ~n2608 & n2614 ) | ( ~n2608 & n2615 ) | ( n2614 & n2615 ) ;
  assign n2617 = ( n2466 & ~n2606 ) | ( n2466 & n2616 ) | ( ~n2606 & n2616 ) ;
  assign n2618 = ( n2466 & n2606 ) | ( n2466 & n2616 ) | ( n2606 & n2616 ) ;
  assign n2619 = ( n2606 & n2617 ) | ( n2606 & ~n2618 ) | ( n2617 & ~n2618 ) ;
  assign n2620 = ( n2468 & n2512 ) | ( n2468 & n2619 ) | ( n2512 & n2619 ) ;
  assign n2621 = ( ~n2468 & n2512 ) | ( ~n2468 & n2619 ) | ( n2512 & n2619 ) ;
  assign n2622 = ( n2468 & ~n2620 ) | ( n2468 & n2621 ) | ( ~n2620 & n2621 ) ;
  assign n2623 = n206 & n2083 ;
  assign n2624 = x5 & n2623 ;
  assign n2625 = x92 & n205 ;
  assign n2626 = x91 & n201 ;
  assign n2627 = n2625 | n2626 ;
  assign n2628 = x90 & n221 ;
  assign n2629 = n2627 | n2628 ;
  assign n2630 = ( ~x5 & n2623 ) | ( ~x5 & n2629 ) | ( n2623 & n2629 ) ;
  assign n2631 = x5 & ~n2629 ;
  assign n2632 = ( ~n2624 & n2630 ) | ( ~n2624 & n2631 ) | ( n2630 & n2631 ) ;
  assign n2633 = ( n2471 & ~n2622 ) | ( n2471 & n2632 ) | ( ~n2622 & n2632 ) ;
  assign n2634 = ( n2471 & n2622 ) | ( n2471 & n2632 ) | ( n2622 & n2632 ) ;
  assign n2635 = ( n2622 & n2633 ) | ( n2622 & ~n2634 ) | ( n2633 & ~n2634 ) ;
  assign n2636 = ( n2488 & n2502 ) | ( n2488 & n2635 ) | ( n2502 & n2635 ) ;
  assign n2637 = ( n2488 & ~n2502 ) | ( n2488 & n2635 ) | ( ~n2502 & n2635 ) ;
  assign n2638 = ( n2502 & ~n2636 ) | ( n2502 & n2637 ) | ( ~n2636 & n2637 ) ;
  assign n2639 = n301 & n1838 ;
  assign n2640 = x8 & n2639 ;
  assign n2641 = x90 & n309 ;
  assign n2642 = x89 & n306 ;
  assign n2643 = n2641 | n2642 ;
  assign n2644 = x88 & n359 ;
  assign n2645 = n2643 | n2644 ;
  assign n2646 = ( ~x8 & n2639 ) | ( ~x8 & n2645 ) | ( n2639 & n2645 ) ;
  assign n2647 = x8 & ~n2645 ;
  assign n2648 = ( ~n2640 & n2646 ) | ( ~n2640 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2649 = n449 & n1494 ;
  assign n2650 = x11 & n2649 ;
  assign n2651 = x87 & n456 ;
  assign n2652 = x86 & n453 ;
  assign n2653 = n2651 | n2652 ;
  assign n2654 = x85 & n536 ;
  assign n2655 = n2653 | n2654 ;
  assign n2656 = ( ~x11 & n2649 ) | ( ~x11 & n2655 ) | ( n2649 & n2655 ) ;
  assign n2657 = x11 & ~n2655 ;
  assign n2658 = ( ~n2650 & n2656 ) | ( ~n2650 & n2657 ) | ( n2656 & n2657 ) ;
  assign n2659 = n649 & n1190 ;
  assign n2660 = x14 & n2659 ;
  assign n2661 = x84 & n656 ;
  assign n2662 = x83 & n653 ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = x82 & n744 ;
  assign n2665 = n2663 | n2664 ;
  assign n2666 = ( ~x14 & n2659 ) | ( ~x14 & n2665 ) | ( n2659 & n2665 ) ;
  assign n2667 = x14 & ~n2665 ;
  assign n2668 = ( ~n2660 & n2666 ) | ( ~n2660 & n2667 ) | ( n2666 & n2667 ) ;
  assign n2669 = n874 & n990 ;
  assign n2670 = x17 & n2669 ;
  assign n2671 = x81 & n881 ;
  assign n2672 = x80 & n878 ;
  assign n2673 = n2671 | n2672 ;
  assign n2674 = x79 & n959 ;
  assign n2675 = n2673 | n2674 ;
  assign n2676 = ( ~x17 & n2669 ) | ( ~x17 & n2675 ) | ( n2669 & n2675 ) ;
  assign n2677 = x17 & ~n2675 ;
  assign n2678 = ( ~n2670 & n2676 ) | ( ~n2670 & n2677 ) | ( n2676 & n2677 ) ;
  assign n2679 = n508 & n1427 ;
  assign n2680 = x23 & n2679 ;
  assign n2681 = x75 & n1434 ;
  assign n2682 = x74 & n1431 ;
  assign n2683 = n2681 | n2682 ;
  assign n2684 = x73 & n1531 ;
  assign n2685 = n2683 | n2684 ;
  assign n2686 = ( ~x23 & n2679 ) | ( ~x23 & n2685 ) | ( n2679 & n2685 ) ;
  assign n2687 = x23 & ~n2685 ;
  assign n2688 = ( ~n2680 & n2686 ) | ( ~n2680 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = x66 & n2552 ;
  assign n2690 = x65 & n2549 ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = n226 & n2545 ;
  assign n2693 = n2691 | n2692 ;
  assign n2694 = n2392 & n2544 ;
  assign n2695 = ~n2391 & n2543 ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = x64 & n2696 ;
  assign n2698 = n2693 | n2697 ;
  assign n2699 = ~x32 & n2698 ;
  assign n2700 = ( x32 & n2555 ) | ( x32 & n2698 ) | ( n2555 & n2698 ) ;
  assign n2701 = n2555 & n2698 ;
  assign n2702 = ( n2699 & n2700 ) | ( n2699 & ~n2701 ) | ( n2700 & ~n2701 ) ;
  assign n2703 = n240 & n2137 ;
  assign n2704 = x29 & n2703 ;
  assign n2705 = x69 & n2144 ;
  assign n2706 = x68 & n2141 ;
  assign n2707 = n2705 | n2706 ;
  assign n2708 = x67 & n2267 ;
  assign n2709 = n2707 | n2708 ;
  assign n2710 = ( ~x29 & n2703 ) | ( ~x29 & n2709 ) | ( n2703 & n2709 ) ;
  assign n2711 = x29 & ~n2709 ;
  assign n2712 = ( ~n2704 & n2710 ) | ( ~n2704 & n2711 ) | ( n2710 & n2711 ) ;
  assign n2713 = ( n2570 & n2702 ) | ( n2570 & n2712 ) | ( n2702 & n2712 ) ;
  assign n2714 = ( ~n2570 & n2702 ) | ( ~n2570 & n2712 ) | ( n2702 & n2712 ) ;
  assign n2715 = ( n2570 & ~n2713 ) | ( n2570 & n2714 ) | ( ~n2713 & n2714 ) ;
  assign n2716 = n372 & n1755 ;
  assign n2717 = x26 & n2716 ;
  assign n2718 = x72 & n1762 ;
  assign n2719 = x71 & n1759 ;
  assign n2720 = n2718 | n2719 ;
  assign n2721 = x70 & n1895 ;
  assign n2722 = n2720 | n2721 ;
  assign n2723 = ( ~x26 & n2716 ) | ( ~x26 & n2722 ) | ( n2716 & n2722 ) ;
  assign n2724 = x26 & ~n2722 ;
  assign n2725 = ( ~n2717 & n2723 ) | ( ~n2717 & n2724 ) | ( n2723 & n2724 ) ;
  assign n2726 = ( n2573 & ~n2715 ) | ( n2573 & n2725 ) | ( ~n2715 & n2725 ) ;
  assign n2727 = ( n2573 & n2715 ) | ( n2573 & n2725 ) | ( n2715 & n2725 ) ;
  assign n2728 = ( n2715 & n2726 ) | ( n2715 & ~n2727 ) | ( n2726 & ~n2727 ) ;
  assign n2729 = ( n2586 & n2688 ) | ( n2586 & n2728 ) | ( n2688 & n2728 ) ;
  assign n2730 = ( ~n2586 & n2688 ) | ( ~n2586 & n2728 ) | ( n2688 & n2728 ) ;
  assign n2731 = ( n2586 & ~n2729 ) | ( n2586 & n2730 ) | ( ~n2729 & n2730 ) ;
  assign n2732 = n697 & n1146 ;
  assign n2733 = x20 & n2732 ;
  assign n2734 = x78 & n1153 ;
  assign n2735 = x77 & n1150 ;
  assign n2736 = n2734 | n2735 ;
  assign n2737 = x76 & n1217 ;
  assign n2738 = n2736 | n2737 ;
  assign n2739 = ( ~x20 & n2732 ) | ( ~x20 & n2738 ) | ( n2732 & n2738 ) ;
  assign n2740 = x20 & ~n2738 ;
  assign n2741 = ( ~n2733 & n2739 ) | ( ~n2733 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2742 = ( n2588 & ~n2731 ) | ( n2588 & n2741 ) | ( ~n2731 & n2741 ) ;
  assign n2743 = ( n2588 & n2731 ) | ( n2588 & n2741 ) | ( n2731 & n2741 ) ;
  assign n2744 = ( n2731 & n2742 ) | ( n2731 & ~n2743 ) | ( n2742 & ~n2743 ) ;
  assign n2745 = ( n2602 & n2678 ) | ( n2602 & n2744 ) | ( n2678 & n2744 ) ;
  assign n2746 = ( ~n2602 & n2678 ) | ( ~n2602 & n2744 ) | ( n2678 & n2744 ) ;
  assign n2747 = ( n2602 & ~n2745 ) | ( n2602 & n2746 ) | ( ~n2745 & n2746 ) ;
  assign n2748 = ( n2604 & n2668 ) | ( n2604 & n2747 ) | ( n2668 & n2747 ) ;
  assign n2749 = ( ~n2604 & n2668 ) | ( ~n2604 & n2747 ) | ( n2668 & n2747 ) ;
  assign n2750 = ( n2604 & ~n2748 ) | ( n2604 & n2749 ) | ( ~n2748 & n2749 ) ;
  assign n2751 = ( n2618 & ~n2658 ) | ( n2618 & n2750 ) | ( ~n2658 & n2750 ) ;
  assign n2752 = ( n2618 & n2658 ) | ( n2618 & n2750 ) | ( n2658 & n2750 ) ;
  assign n2753 = ( n2658 & n2751 ) | ( n2658 & ~n2752 ) | ( n2751 & ~n2752 ) ;
  assign n2754 = ( n2620 & n2648 ) | ( n2620 & n2753 ) | ( n2648 & n2753 ) ;
  assign n2755 = ( ~n2620 & n2648 ) | ( ~n2620 & n2753 ) | ( n2648 & n2753 ) ;
  assign n2756 = ( n2620 & ~n2754 ) | ( n2620 & n2755 ) | ( ~n2754 & n2755 ) ;
  assign n2757 = n206 & n2220 ;
  assign n2758 = x5 & n2757 ;
  assign n2759 = x93 & n205 ;
  assign n2760 = x92 & n201 ;
  assign n2761 = n2759 | n2760 ;
  assign n2762 = x91 & n221 ;
  assign n2763 = n2761 | n2762 ;
  assign n2764 = ( ~x5 & n2757 ) | ( ~x5 & n2763 ) | ( n2757 & n2763 ) ;
  assign n2765 = x5 & ~n2763 ;
  assign n2766 = ( ~n2758 & n2764 ) | ( ~n2758 & n2765 ) | ( n2764 & n2765 ) ;
  assign n2767 = ( n2634 & n2756 ) | ( n2634 & n2766 ) | ( n2756 & n2766 ) ;
  assign n2768 = ( ~n2634 & n2756 ) | ( ~n2634 & n2766 ) | ( n2756 & n2766 ) ;
  assign n2769 = ( n2634 & ~n2767 ) | ( n2634 & n2768 ) | ( ~n2767 & n2768 ) ;
  assign n2770 = ( ~x95 & x96 ) | ( ~x95 & n2491 ) | ( x96 & n2491 ) ;
  assign n2771 = ( x95 & x96 ) | ( x95 & n2491 ) | ( x96 & n2491 ) ;
  assign n2772 = ( x95 & n2770 ) | ( x95 & ~n2771 ) | ( n2770 & ~n2771 ) ;
  assign n2773 = x0 & n2772 ;
  assign n2774 = ( x1 & x2 ) | ( x1 & n2773 ) | ( x2 & n2773 ) ;
  assign n2775 = x95 & n172 ;
  assign n2776 = ( ~x94 & n135 ) | ( ~x94 & n174 ) | ( n135 & n174 ) ;
  assign n2777 = n2775 | n2776 ;
  assign n2778 = x96 & n147 ;
  assign n2779 = n2777 | n2778 ;
  assign n2780 = n2774 | n2779 ;
  assign n2781 = n2774 & n2779 ;
  assign n2782 = n2780 & ~n2781 ;
  assign n2783 = ( n2636 & ~n2769 ) | ( n2636 & n2782 ) | ( ~n2769 & n2782 ) ;
  assign n2784 = ( n2636 & n2769 ) | ( n2636 & n2782 ) | ( n2769 & n2782 ) ;
  assign n2785 = ( n2769 & n2783 ) | ( n2769 & ~n2784 ) | ( n2783 & ~n2784 ) ;
  assign n2786 = ( ~x96 & x97 ) | ( ~x96 & n2771 ) | ( x97 & n2771 ) ;
  assign n2787 = ( x96 & x97 ) | ( x96 & n2771 ) | ( x97 & n2771 ) ;
  assign n2788 = ( x96 & n2786 ) | ( x96 & ~n2787 ) | ( n2786 & ~n2787 ) ;
  assign n2789 = x0 & n2788 ;
  assign n2790 = ( x1 & x2 ) | ( x1 & n2789 ) | ( x2 & n2789 ) ;
  assign n2791 = x96 & n172 ;
  assign n2792 = ( ~x95 & n135 ) | ( ~x95 & n174 ) | ( n135 & n174 ) ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = x97 & n147 ;
  assign n2795 = n2793 | n2794 ;
  assign n2796 = n2790 | n2795 ;
  assign n2797 = n2790 & n2795 ;
  assign n2798 = n2796 & ~n2797 ;
  assign n2799 = n206 & n2476 ;
  assign n2800 = x5 & n2799 ;
  assign n2801 = x94 & n205 ;
  assign n2802 = x93 & n201 ;
  assign n2803 = n2801 | n2802 ;
  assign n2804 = x92 & n221 ;
  assign n2805 = n2803 | n2804 ;
  assign n2806 = ( ~x5 & n2799 ) | ( ~x5 & n2805 ) | ( n2799 & n2805 ) ;
  assign n2807 = x5 & ~n2805 ;
  assign n2808 = ( ~n2800 & n2806 ) | ( ~n2800 & n2807 ) | ( n2806 & n2807 ) ;
  assign n2809 = n301 & n1959 ;
  assign n2810 = x8 & n2809 ;
  assign n2811 = x91 & n309 ;
  assign n2812 = x90 & n306 ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = x89 & n359 ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = ( ~x8 & n2809 ) | ( ~x8 & n2815 ) | ( n2809 & n2815 ) ;
  assign n2817 = x8 & ~n2815 ;
  assign n2818 = ( ~n2810 & n2816 ) | ( ~n2810 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2819 = n823 & n1146 ;
  assign n2820 = x20 & n2819 ;
  assign n2821 = x79 & n1153 ;
  assign n2822 = x78 & n1150 ;
  assign n2823 = n2821 | n2822 ;
  assign n2824 = x77 & n1217 ;
  assign n2825 = n2823 | n2824 ;
  assign n2826 = ( ~x20 & n2819 ) | ( ~x20 & n2825 ) | ( n2819 & n2825 ) ;
  assign n2827 = x20 & ~n2825 ;
  assign n2828 = ( ~n2820 & n2826 ) | ( ~n2820 & n2827 ) | ( n2826 & n2827 ) ;
  assign n2829 = n565 & n1427 ;
  assign n2830 = x23 & n2829 ;
  assign n2831 = x76 & n1434 ;
  assign n2832 = x75 & n1431 ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = x74 & n1531 ;
  assign n2835 = n2833 | n2834 ;
  assign n2836 = ( ~x23 & n2829 ) | ( ~x23 & n2835 ) | ( n2829 & n2835 ) ;
  assign n2837 = x23 & ~n2835 ;
  assign n2838 = ( ~n2830 & n2836 ) | ( ~n2830 & n2837 ) | ( n2836 & n2837 ) ;
  assign n2839 = n276 & n2137 ;
  assign n2840 = x29 & n2839 ;
  assign n2841 = x70 & n2144 ;
  assign n2842 = x69 & n2141 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = x68 & n2267 ;
  assign n2845 = n2843 | n2844 ;
  assign n2846 = ( ~x29 & n2839 ) | ( ~x29 & n2845 ) | ( n2839 & n2845 ) ;
  assign n2847 = x29 & ~n2845 ;
  assign n2848 = ( ~n2840 & n2846 ) | ( ~n2840 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = n2555 | n2698 ;
  assign n2850 = x32 & n2849 ;
  assign n2851 = x66 & n2549 ;
  assign n2852 = n169 & n2545 ;
  assign n2853 = x67 & n2552 ;
  assign n2854 = x65 & ~n2696 ;
  assign n2855 = ( x65 & n2853 ) | ( x65 & ~n2854 ) | ( n2853 & ~n2854 ) ;
  assign n2856 = n2852 | n2855 ;
  assign n2857 = n2851 | n2856 ;
  assign n2858 = x32 | x33 ;
  assign n2859 = x32 & x33 ;
  assign n2860 = n2858 & ~n2859 ;
  assign n2861 = x64 & n2860 ;
  assign n2862 = ( n2850 & ~n2857 ) | ( n2850 & n2861 ) | ( ~n2857 & n2861 ) ;
  assign n2863 = x32 & ~n2857 ;
  assign n2864 = ( ~n2850 & n2857 ) | ( ~n2850 & n2863 ) | ( n2857 & n2863 ) ;
  assign n2865 = ( n2861 & n2863 ) | ( n2861 & n2864 ) | ( n2863 & n2864 ) ;
  assign n2866 = ( n2862 & n2864 ) | ( n2862 & ~n2865 ) | ( n2864 & ~n2865 ) ;
  assign n2867 = ( n2713 & n2848 ) | ( n2713 & n2866 ) | ( n2848 & n2866 ) ;
  assign n2868 = ( ~n2713 & n2848 ) | ( ~n2713 & n2866 ) | ( n2848 & n2866 ) ;
  assign n2869 = ( n2713 & ~n2867 ) | ( n2713 & n2868 ) | ( ~n2867 & n2868 ) ;
  assign n2870 = n388 & n1755 ;
  assign n2871 = x26 & n2870 ;
  assign n2872 = x73 & n1762 ;
  assign n2873 = x72 & n1759 ;
  assign n2874 = n2872 | n2873 ;
  assign n2875 = x71 & n1895 ;
  assign n2876 = n2874 | n2875 ;
  assign n2877 = ( ~x26 & n2870 ) | ( ~x26 & n2876 ) | ( n2870 & n2876 ) ;
  assign n2878 = x26 & ~n2876 ;
  assign n2879 = ( ~n2871 & n2877 ) | ( ~n2871 & n2878 ) | ( n2877 & n2878 ) ;
  assign n2880 = ( n2727 & ~n2869 ) | ( n2727 & n2879 ) | ( ~n2869 & n2879 ) ;
  assign n2881 = ( n2727 & n2869 ) | ( n2727 & n2879 ) | ( n2869 & n2879 ) ;
  assign n2882 = ( n2869 & n2880 ) | ( n2869 & ~n2881 ) | ( n2880 & ~n2881 ) ;
  assign n2883 = ( n2729 & n2838 ) | ( n2729 & n2882 ) | ( n2838 & n2882 ) ;
  assign n2884 = ( ~n2729 & n2838 ) | ( ~n2729 & n2882 ) | ( n2838 & n2882 ) ;
  assign n2885 = ( n2729 & ~n2883 ) | ( n2729 & n2884 ) | ( ~n2883 & n2884 ) ;
  assign n2886 = ( n2743 & n2828 ) | ( n2743 & n2885 ) | ( n2828 & n2885 ) ;
  assign n2887 = ( ~n2743 & n2828 ) | ( ~n2743 & n2885 ) | ( n2828 & n2885 ) ;
  assign n2888 = ( n2743 & ~n2886 ) | ( n2743 & n2887 ) | ( ~n2886 & n2887 ) ;
  assign n2889 = n874 & n1006 ;
  assign n2890 = x17 & n2889 ;
  assign n2891 = x82 & n881 ;
  assign n2892 = x81 & n878 ;
  assign n2893 = n2891 | n2892 ;
  assign n2894 = x80 & n959 ;
  assign n2895 = n2893 | n2894 ;
  assign n2896 = ( ~x17 & n2889 ) | ( ~x17 & n2895 ) | ( n2889 & n2895 ) ;
  assign n2897 = x17 & ~n2895 ;
  assign n2898 = ( ~n2890 & n2896 ) | ( ~n2890 & n2897 ) | ( n2896 & n2897 ) ;
  assign n2899 = ( n2745 & n2888 ) | ( n2745 & n2898 ) | ( n2888 & n2898 ) ;
  assign n2900 = ( ~n2745 & n2888 ) | ( ~n2745 & n2898 ) | ( n2888 & n2898 ) ;
  assign n2901 = ( n2745 & ~n2899 ) | ( n2745 & n2900 ) | ( ~n2899 & n2900 ) ;
  assign n2902 = n649 & n1368 ;
  assign n2903 = x14 & n2902 ;
  assign n2904 = x85 & n656 ;
  assign n2905 = x84 & n653 ;
  assign n2906 = n2904 | n2905 ;
  assign n2907 = x83 & n744 ;
  assign n2908 = n2906 | n2907 ;
  assign n2909 = ( ~x14 & n2902 ) | ( ~x14 & n2908 ) | ( n2902 & n2908 ) ;
  assign n2910 = x14 & ~n2908 ;
  assign n2911 = ( ~n2903 & n2909 ) | ( ~n2903 & n2910 ) | ( n2909 & n2910 ) ;
  assign n2912 = ( n2748 & ~n2901 ) | ( n2748 & n2911 ) | ( ~n2901 & n2911 ) ;
  assign n2913 = ( n2748 & n2901 ) | ( n2748 & n2911 ) | ( n2901 & n2911 ) ;
  assign n2914 = ( n2901 & n2912 ) | ( n2901 & ~n2913 ) | ( n2912 & ~n2913 ) ;
  assign n2915 = n449 & n1602 ;
  assign n2916 = x11 & n2915 ;
  assign n2917 = x88 & n456 ;
  assign n2918 = x87 & n453 ;
  assign n2919 = n2917 | n2918 ;
  assign n2920 = x86 & n536 ;
  assign n2921 = n2919 | n2920 ;
  assign n2922 = ( ~x11 & n2915 ) | ( ~x11 & n2921 ) | ( n2915 & n2921 ) ;
  assign n2923 = x11 & ~n2921 ;
  assign n2924 = ( ~n2916 & n2922 ) | ( ~n2916 & n2923 ) | ( n2922 & n2923 ) ;
  assign n2925 = ( n2752 & ~n2914 ) | ( n2752 & n2924 ) | ( ~n2914 & n2924 ) ;
  assign n2926 = ( n2752 & n2914 ) | ( n2752 & n2924 ) | ( n2914 & n2924 ) ;
  assign n2927 = ( n2914 & n2925 ) | ( n2914 & ~n2926 ) | ( n2925 & ~n2926 ) ;
  assign n2928 = ( n2754 & n2818 ) | ( n2754 & n2927 ) | ( n2818 & n2927 ) ;
  assign n2929 = ( ~n2754 & n2818 ) | ( ~n2754 & n2927 ) | ( n2818 & n2927 ) ;
  assign n2930 = ( n2754 & ~n2928 ) | ( n2754 & n2929 ) | ( ~n2928 & n2929 ) ;
  assign n2931 = ( n2767 & ~n2808 ) | ( n2767 & n2930 ) | ( ~n2808 & n2930 ) ;
  assign n2932 = ( n2767 & n2808 ) | ( n2767 & n2930 ) | ( n2808 & n2930 ) ;
  assign n2933 = ( n2808 & n2931 ) | ( n2808 & ~n2932 ) | ( n2931 & ~n2932 ) ;
  assign n2934 = ( n2784 & n2798 ) | ( n2784 & n2933 ) | ( n2798 & n2933 ) ;
  assign n2935 = ( ~n2784 & n2798 ) | ( ~n2784 & n2933 ) | ( n2798 & n2933 ) ;
  assign n2936 = ( n2784 & ~n2934 ) | ( n2784 & n2935 ) | ( ~n2934 & n2935 ) ;
  assign n2937 = ( ~x97 & x98 ) | ( ~x97 & n2787 ) | ( x98 & n2787 ) ;
  assign n2938 = ( x97 & x98 ) | ( x97 & n2787 ) | ( x98 & n2787 ) ;
  assign n2939 = ( x97 & n2937 ) | ( x97 & ~n2938 ) | ( n2937 & ~n2938 ) ;
  assign n2940 = x0 & n2939 ;
  assign n2941 = ( x1 & x2 ) | ( x1 & n2940 ) | ( x2 & n2940 ) ;
  assign n2942 = x97 & n172 ;
  assign n2943 = ( ~x96 & n135 ) | ( ~x96 & n174 ) | ( n135 & n174 ) ;
  assign n2944 = n2942 | n2943 ;
  assign n2945 = x98 & n147 ;
  assign n2946 = n2944 | n2945 ;
  assign n2947 = n2941 | n2946 ;
  assign n2948 = n2941 & n2946 ;
  assign n2949 = n2947 & ~n2948 ;
  assign n2950 = n874 & n1093 ;
  assign n2951 = x17 & n2950 ;
  assign n2952 = x83 & n881 ;
  assign n2953 = x82 & n878 ;
  assign n2954 = n2952 | n2953 ;
  assign n2955 = x81 & n959 ;
  assign n2956 = n2954 | n2955 ;
  assign n2957 = ( ~x17 & n2950 ) | ( ~x17 & n2956 ) | ( n2950 & n2956 ) ;
  assign n2958 = x17 & ~n2956 ;
  assign n2959 = ( ~n2951 & n2957 ) | ( ~n2951 & n2958 ) | ( n2957 & n2958 ) ;
  assign n2960 = n840 & n1146 ;
  assign n2961 = x20 & n2960 ;
  assign n2962 = x80 & n1153 ;
  assign n2963 = x79 & n1150 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = x78 & n1217 ;
  assign n2966 = n2964 | n2965 ;
  assign n2967 = ( ~x20 & n2960 ) | ( ~x20 & n2966 ) | ( n2960 & n2966 ) ;
  assign n2968 = x20 & ~n2966 ;
  assign n2969 = ( ~n2961 & n2967 ) | ( ~n2961 & n2968 ) | ( n2967 & n2968 ) ;
  assign n2970 = n322 & n2137 ;
  assign n2971 = x29 & n2970 ;
  assign n2972 = x71 & n2144 ;
  assign n2973 = x70 & n2141 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = x69 & n2267 ;
  assign n2976 = n2974 | n2975 ;
  assign n2977 = ( ~x29 & n2970 ) | ( ~x29 & n2976 ) | ( n2970 & n2976 ) ;
  assign n2978 = x29 & ~n2976 ;
  assign n2979 = ( ~n2971 & n2977 ) | ( ~n2971 & n2978 ) | ( n2977 & n2978 ) ;
  assign n2980 = ~x34 & x35 ;
  assign n2981 = x34 & ~x35 ;
  assign n2982 = ( n2860 & n2980 ) | ( n2860 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2983 = n302 & n2982 ;
  assign n2984 = ~x32 & x34 ;
  assign n2985 = x33 & x34 ;
  assign n2986 = ( n2859 & n2984 ) | ( n2859 & ~n2985 ) | ( n2984 & ~n2985 ) ;
  assign n2987 = x64 & n2986 ;
  assign n2988 = n2983 | n2987 ;
  assign n2989 = n2860 & ~n2982 ;
  assign n2990 = x65 & n2989 ;
  assign n2991 = n2988 | n2990 ;
  assign n2992 = n2861 | n2991 ;
  assign n2993 = ( x35 & n2861 ) | ( x35 & ~n2991 ) | ( n2861 & ~n2991 ) ;
  assign n2994 = x35 & ~n2991 ;
  assign n2995 = ( n2992 & ~n2993 ) | ( n2992 & n2994 ) | ( ~n2993 & n2994 ) ;
  assign n2996 = x68 & n2552 ;
  assign n2997 = x32 & n2996 ;
  assign n2998 = x67 & n2549 ;
  assign n2999 = x66 & n2696 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = n193 & n2545 ;
  assign n3002 = n3000 | n3001 ;
  assign n3003 = ( ~x32 & n2996 ) | ( ~x32 & n3002 ) | ( n2996 & n3002 ) ;
  assign n3004 = x32 & ~n3002 ;
  assign n3005 = ( ~n2997 & n3003 ) | ( ~n2997 & n3004 ) | ( n3003 & n3004 ) ;
  assign n3006 = ( n2865 & ~n2995 ) | ( n2865 & n3005 ) | ( ~n2995 & n3005 ) ;
  assign n3007 = ( n2865 & n2995 ) | ( n2865 & n3005 ) | ( n2995 & n3005 ) ;
  assign n3008 = ( n2995 & n3006 ) | ( n2995 & ~n3007 ) | ( n3006 & ~n3007 ) ;
  assign n3009 = ( n2867 & n2979 ) | ( n2867 & n3008 ) | ( n2979 & n3008 ) ;
  assign n3010 = ( ~n2867 & n2979 ) | ( ~n2867 & n3008 ) | ( n2979 & n3008 ) ;
  assign n3011 = ( n2867 & ~n3009 ) | ( n2867 & n3010 ) | ( ~n3009 & n3010 ) ;
  assign n3012 = n436 & n1755 ;
  assign n3013 = x26 & n3012 ;
  assign n3014 = x74 & n1762 ;
  assign n3015 = x73 & n1759 ;
  assign n3016 = n3014 | n3015 ;
  assign n3017 = x72 & n1895 ;
  assign n3018 = n3016 | n3017 ;
  assign n3019 = ( ~x26 & n3012 ) | ( ~x26 & n3018 ) | ( n3012 & n3018 ) ;
  assign n3020 = x26 & ~n3018 ;
  assign n3021 = ( ~n3013 & n3019 ) | ( ~n3013 & n3020 ) | ( n3019 & n3020 ) ;
  assign n3022 = ( n2881 & n3011 ) | ( n2881 & n3021 ) | ( n3011 & n3021 ) ;
  assign n3023 = ( ~n2881 & n3011 ) | ( ~n2881 & n3021 ) | ( n3011 & n3021 ) ;
  assign n3024 = ( n2881 & ~n3022 ) | ( n2881 & n3023 ) | ( ~n3022 & n3023 ) ;
  assign n3025 = n626 & n1427 ;
  assign n3026 = x23 & n3025 ;
  assign n3027 = x77 & n1434 ;
  assign n3028 = x76 & n1431 ;
  assign n3029 = n3027 | n3028 ;
  assign n3030 = x75 & n1531 ;
  assign n3031 = n3029 | n3030 ;
  assign n3032 = ( ~x23 & n3025 ) | ( ~x23 & n3031 ) | ( n3025 & n3031 ) ;
  assign n3033 = x23 & ~n3031 ;
  assign n3034 = ( ~n3026 & n3032 ) | ( ~n3026 & n3033 ) | ( n3032 & n3033 ) ;
  assign n3035 = ( n2883 & ~n3024 ) | ( n2883 & n3034 ) | ( ~n3024 & n3034 ) ;
  assign n3036 = ( n2883 & n3024 ) | ( n2883 & n3034 ) | ( n3024 & n3034 ) ;
  assign n3037 = ( n3024 & n3035 ) | ( n3024 & ~n3036 ) | ( n3035 & ~n3036 ) ;
  assign n3038 = ( n2886 & n2969 ) | ( n2886 & n3037 ) | ( n2969 & n3037 ) ;
  assign n3039 = ( ~n2886 & n2969 ) | ( ~n2886 & n3037 ) | ( n2969 & n3037 ) ;
  assign n3040 = ( n2886 & ~n3038 ) | ( n2886 & n3039 ) | ( ~n3038 & n3039 ) ;
  assign n3041 = ( n2899 & n2959 ) | ( n2899 & n3040 ) | ( n2959 & n3040 ) ;
  assign n3042 = ( ~n2899 & n2959 ) | ( ~n2899 & n3040 ) | ( n2959 & n3040 ) ;
  assign n3043 = ( n2899 & ~n3041 ) | ( n2899 & n3042 ) | ( ~n3041 & n3042 ) ;
  assign n3044 = n649 & n1384 ;
  assign n3045 = x14 & n3044 ;
  assign n3046 = x86 & n656 ;
  assign n3047 = x85 & n653 ;
  assign n3048 = n3046 | n3047 ;
  assign n3049 = x84 & n744 ;
  assign n3050 = n3048 | n3049 ;
  assign n3051 = ( ~x14 & n3044 ) | ( ~x14 & n3050 ) | ( n3044 & n3050 ) ;
  assign n3052 = x14 & ~n3050 ;
  assign n3053 = ( ~n3045 & n3051 ) | ( ~n3045 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3054 = ( n2913 & n3043 ) | ( n2913 & n3053 ) | ( n3043 & n3053 ) ;
  assign n3055 = ( ~n2913 & n3043 ) | ( ~n2913 & n3053 ) | ( n3043 & n3053 ) ;
  assign n3056 = ( n2913 & ~n3054 ) | ( n2913 & n3055 ) | ( ~n3054 & n3055 ) ;
  assign n3057 = n449 & n1822 ;
  assign n3058 = x11 & n3057 ;
  assign n3059 = x89 & n456 ;
  assign n3060 = x88 & n453 ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = x87 & n536 ;
  assign n3063 = n3061 | n3062 ;
  assign n3064 = ( ~x11 & n3057 ) | ( ~x11 & n3063 ) | ( n3057 & n3063 ) ;
  assign n3065 = x11 & ~n3063 ;
  assign n3066 = ( ~n3058 & n3064 ) | ( ~n3058 & n3065 ) | ( n3064 & n3065 ) ;
  assign n3067 = ( n2926 & n3056 ) | ( n2926 & n3066 ) | ( n3056 & n3066 ) ;
  assign n3068 = ( ~n2926 & n3056 ) | ( ~n2926 & n3066 ) | ( n3056 & n3066 ) ;
  assign n3069 = ( n2926 & ~n3067 ) | ( n2926 & n3068 ) | ( ~n3067 & n3068 ) ;
  assign n3070 = n301 & n2083 ;
  assign n3071 = x8 & n3070 ;
  assign n3072 = x92 & n309 ;
  assign n3073 = x91 & n306 ;
  assign n3074 = n3072 | n3073 ;
  assign n3075 = x90 & n359 ;
  assign n3076 = n3074 | n3075 ;
  assign n3077 = ( ~x8 & n3070 ) | ( ~x8 & n3076 ) | ( n3070 & n3076 ) ;
  assign n3078 = x8 & ~n3076 ;
  assign n3079 = ( ~n3071 & n3077 ) | ( ~n3071 & n3078 ) | ( n3077 & n3078 ) ;
  assign n3080 = ( n2928 & ~n3069 ) | ( n2928 & n3079 ) | ( ~n3069 & n3079 ) ;
  assign n3081 = ( n2928 & n3069 ) | ( n2928 & n3079 ) | ( n3069 & n3079 ) ;
  assign n3082 = ( n3069 & n3080 ) | ( n3069 & ~n3081 ) | ( n3080 & ~n3081 ) ;
  assign n3083 = n206 & n2492 ;
  assign n3084 = x5 & n3083 ;
  assign n3085 = x95 & n205 ;
  assign n3086 = x94 & n201 ;
  assign n3087 = n3085 | n3086 ;
  assign n3088 = x93 & n221 ;
  assign n3089 = n3087 | n3088 ;
  assign n3090 = ( ~x5 & n3083 ) | ( ~x5 & n3089 ) | ( n3083 & n3089 ) ;
  assign n3091 = x5 & ~n3089 ;
  assign n3092 = ( ~n3084 & n3090 ) | ( ~n3084 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3093 = ( n2932 & ~n3082 ) | ( n2932 & n3092 ) | ( ~n3082 & n3092 ) ;
  assign n3094 = ( n2932 & n3082 ) | ( n2932 & n3092 ) | ( n3082 & n3092 ) ;
  assign n3095 = ( n3082 & n3093 ) | ( n3082 & ~n3094 ) | ( n3093 & ~n3094 ) ;
  assign n3096 = ( n2934 & n2949 ) | ( n2934 & n3095 ) | ( n2949 & n3095 ) ;
  assign n3097 = ( ~n2934 & n2949 ) | ( ~n2934 & n3095 ) | ( n2949 & n3095 ) ;
  assign n3098 = ( n2934 & ~n3096 ) | ( n2934 & n3097 ) | ( ~n3096 & n3097 ) ;
  assign n3099 = n301 & n2220 ;
  assign n3100 = x8 & n3099 ;
  assign n3101 = x93 & n309 ;
  assign n3102 = x92 & n306 ;
  assign n3103 = n3101 | n3102 ;
  assign n3104 = x91 & n359 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = ( ~x8 & n3099 ) | ( ~x8 & n3105 ) | ( n3099 & n3105 ) ;
  assign n3107 = x8 & ~n3105 ;
  assign n3108 = ( ~n3100 & n3106 ) | ( ~n3100 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3109 = n449 & n1838 ;
  assign n3110 = x11 & n3109 ;
  assign n3111 = x90 & n456 ;
  assign n3112 = x89 & n453 ;
  assign n3113 = n3111 | n3112 ;
  assign n3114 = x88 & n536 ;
  assign n3115 = n3113 | n3114 ;
  assign n3116 = ( ~x11 & n3109 ) | ( ~x11 & n3115 ) | ( n3109 & n3115 ) ;
  assign n3117 = x11 & ~n3115 ;
  assign n3118 = ( ~n3110 & n3116 ) | ( ~n3110 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3119 = n990 & n1146 ;
  assign n3120 = x20 & n3119 ;
  assign n3121 = x81 & n1153 ;
  assign n3122 = x80 & n1150 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = x79 & n1217 ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = ( ~x20 & n3119 ) | ( ~x20 & n3125 ) | ( n3119 & n3125 ) ;
  assign n3127 = x20 & ~n3125 ;
  assign n3128 = ( ~n3120 & n3126 ) | ( ~n3120 & n3127 ) | ( n3126 & n3127 ) ;
  assign n3129 = n372 & n2137 ;
  assign n3130 = x29 & n3129 ;
  assign n3131 = x72 & n2144 ;
  assign n3132 = x71 & n2141 ;
  assign n3133 = n3131 | n3132 ;
  assign n3134 = x70 & n2267 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = ( ~x29 & n3129 ) | ( ~x29 & n3135 ) | ( n3129 & n3135 ) ;
  assign n3137 = x29 & ~n3135 ;
  assign n3138 = ( ~n3130 & n3136 ) | ( ~n3130 & n3137 ) | ( n3136 & n3137 ) ;
  assign n3139 = n240 & n2545 ;
  assign n3140 = x32 & n3139 ;
  assign n3141 = x69 & n2552 ;
  assign n3142 = x68 & n2549 ;
  assign n3143 = n3141 | n3142 ;
  assign n3144 = x67 & n2696 ;
  assign n3145 = n3143 | n3144 ;
  assign n3146 = ( ~x32 & n3139 ) | ( ~x32 & n3145 ) | ( n3139 & n3145 ) ;
  assign n3147 = x32 & ~n3145 ;
  assign n3148 = ( ~n3140 & n3146 ) | ( ~n3140 & n3147 ) | ( n3146 & n3147 ) ;
  assign n3149 = ~n3138 & n3148 ;
  assign n3150 = n3138 & ~n3148 ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = x65 & n2986 ;
  assign n3153 = n226 & n2982 ;
  assign n3154 = n3152 | n3153 ;
  assign n3155 = x66 & n2989 ;
  assign n3156 = n3154 | n3155 ;
  assign n3157 = n2859 & n2981 ;
  assign n3158 = ~n2858 & n2980 ;
  assign n3159 = n3157 | n3158 ;
  assign n3160 = x64 & n3159 ;
  assign n3161 = n3156 | n3160 ;
  assign n3162 = ~x35 & n3161 ;
  assign n3163 = ( x35 & n2992 ) | ( x35 & n3161 ) | ( n2992 & n3161 ) ;
  assign n3164 = n2992 & n3161 ;
  assign n3165 = ( n3162 & n3163 ) | ( n3162 & ~n3164 ) | ( n3163 & ~n3164 ) ;
  assign n3166 = n3007 & ~n3165 ;
  assign n3167 = ~n3007 & n3165 ;
  assign n3168 = n3166 | n3167 ;
  assign n3169 = ( ~n3009 & n3151 ) | ( ~n3009 & n3168 ) | ( n3151 & n3168 ) ;
  assign n3170 = ( n3009 & n3151 ) | ( n3009 & ~n3168 ) | ( n3151 & ~n3168 ) ;
  assign n3171 = ( ~n3151 & n3169 ) | ( ~n3151 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3172 = n508 & n1755 ;
  assign n3173 = x26 & n3172 ;
  assign n3174 = x75 & n1762 ;
  assign n3175 = x74 & n1759 ;
  assign n3176 = n3174 | n3175 ;
  assign n3177 = x73 & n1895 ;
  assign n3178 = n3176 | n3177 ;
  assign n3179 = ( ~x26 & n3172 ) | ( ~x26 & n3178 ) | ( n3172 & n3178 ) ;
  assign n3180 = x26 & ~n3178 ;
  assign n3181 = ( ~n3173 & n3179 ) | ( ~n3173 & n3180 ) | ( n3179 & n3180 ) ;
  assign n3182 = ( n3022 & n3171 ) | ( n3022 & n3181 ) | ( n3171 & n3181 ) ;
  assign n3183 = ( ~n3022 & n3171 ) | ( ~n3022 & n3181 ) | ( n3171 & n3181 ) ;
  assign n3184 = ( n3022 & ~n3182 ) | ( n3022 & n3183 ) | ( ~n3182 & n3183 ) ;
  assign n3185 = n697 & n1427 ;
  assign n3186 = x23 & n3185 ;
  assign n3187 = x78 & n1434 ;
  assign n3188 = x77 & n1431 ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = x76 & n1531 ;
  assign n3191 = n3189 | n3190 ;
  assign n3192 = ( ~x23 & n3185 ) | ( ~x23 & n3191 ) | ( n3185 & n3191 ) ;
  assign n3193 = x23 & ~n3191 ;
  assign n3194 = ( ~n3186 & n3192 ) | ( ~n3186 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3195 = ( n3036 & ~n3184 ) | ( n3036 & n3194 ) | ( ~n3184 & n3194 ) ;
  assign n3196 = ( n3036 & n3184 ) | ( n3036 & n3194 ) | ( n3184 & n3194 ) ;
  assign n3197 = ( n3184 & n3195 ) | ( n3184 & ~n3196 ) | ( n3195 & ~n3196 ) ;
  assign n3198 = ( ~n3038 & n3128 ) | ( ~n3038 & n3197 ) | ( n3128 & n3197 ) ;
  assign n3199 = ( n3038 & n3128 ) | ( n3038 & n3197 ) | ( n3128 & n3197 ) ;
  assign n3200 = ( n3038 & n3198 ) | ( n3038 & ~n3199 ) | ( n3198 & ~n3199 ) ;
  assign n3201 = n874 & n1190 ;
  assign n3202 = x17 & n3201 ;
  assign n3203 = x84 & n881 ;
  assign n3204 = x83 & n878 ;
  assign n3205 = n3203 | n3204 ;
  assign n3206 = x82 & n959 ;
  assign n3207 = n3205 | n3206 ;
  assign n3208 = ( ~x17 & n3201 ) | ( ~x17 & n3207 ) | ( n3201 & n3207 ) ;
  assign n3209 = x17 & ~n3207 ;
  assign n3210 = ( ~n3202 & n3208 ) | ( ~n3202 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = ( ~n3041 & n3200 ) | ( ~n3041 & n3210 ) | ( n3200 & n3210 ) ;
  assign n3212 = ( n3041 & n3200 ) | ( n3041 & n3210 ) | ( n3200 & n3210 ) ;
  assign n3213 = ( n3041 & n3211 ) | ( n3041 & ~n3212 ) | ( n3211 & ~n3212 ) ;
  assign n3214 = n649 & n1494 ;
  assign n3215 = x14 & n3214 ;
  assign n3216 = x87 & n656 ;
  assign n3217 = x86 & n653 ;
  assign n3218 = n3216 | n3217 ;
  assign n3219 = x85 & n744 ;
  assign n3220 = n3218 | n3219 ;
  assign n3221 = ( ~x14 & n3214 ) | ( ~x14 & n3220 ) | ( n3214 & n3220 ) ;
  assign n3222 = x14 & ~n3220 ;
  assign n3223 = ( ~n3215 & n3221 ) | ( ~n3215 & n3222 ) | ( n3221 & n3222 ) ;
  assign n3224 = ( ~n3054 & n3213 ) | ( ~n3054 & n3223 ) | ( n3213 & n3223 ) ;
  assign n3225 = ( n3054 & n3213 ) | ( n3054 & n3223 ) | ( n3213 & n3223 ) ;
  assign n3226 = ( n3054 & n3224 ) | ( n3054 & ~n3225 ) | ( n3224 & ~n3225 ) ;
  assign n3227 = ( n3067 & ~n3118 ) | ( n3067 & n3226 ) | ( ~n3118 & n3226 ) ;
  assign n3228 = ( n3067 & n3118 ) | ( n3067 & n3226 ) | ( n3118 & n3226 ) ;
  assign n3229 = ( n3118 & n3227 ) | ( n3118 & ~n3228 ) | ( n3227 & ~n3228 ) ;
  assign n3230 = ( n3081 & n3108 ) | ( n3081 & n3229 ) | ( n3108 & n3229 ) ;
  assign n3231 = ( ~n3081 & n3108 ) | ( ~n3081 & n3229 ) | ( n3108 & n3229 ) ;
  assign n3232 = ( n3081 & ~n3230 ) | ( n3081 & n3231 ) | ( ~n3230 & n3231 ) ;
  assign n3233 = n206 & n2772 ;
  assign n3234 = x5 & n3233 ;
  assign n3235 = x96 & n205 ;
  assign n3236 = x95 & n201 ;
  assign n3237 = n3235 | n3236 ;
  assign n3238 = x94 & n221 ;
  assign n3239 = n3237 | n3238 ;
  assign n3240 = ( ~x5 & n3233 ) | ( ~x5 & n3239 ) | ( n3233 & n3239 ) ;
  assign n3241 = x5 & ~n3239 ;
  assign n3242 = ( ~n3234 & n3240 ) | ( ~n3234 & n3241 ) | ( n3240 & n3241 ) ;
  assign n3243 = ( n3094 & n3232 ) | ( n3094 & n3242 ) | ( n3232 & n3242 ) ;
  assign n3244 = ( ~n3094 & n3232 ) | ( ~n3094 & n3242 ) | ( n3232 & n3242 ) ;
  assign n3245 = ( n3094 & ~n3243 ) | ( n3094 & n3244 ) | ( ~n3243 & n3244 ) ;
  assign n3246 = ( ~x98 & x99 ) | ( ~x98 & n2938 ) | ( x99 & n2938 ) ;
  assign n3247 = ( x98 & x99 ) | ( x98 & n2938 ) | ( x99 & n2938 ) ;
  assign n3248 = ( x98 & n3246 ) | ( x98 & ~n3247 ) | ( n3246 & ~n3247 ) ;
  assign n3249 = x0 & n3248 ;
  assign n3250 = ( x1 & x2 ) | ( x1 & n3249 ) | ( x2 & n3249 ) ;
  assign n3251 = x98 & n172 ;
  assign n3252 = ( ~x97 & n135 ) | ( ~x97 & n174 ) | ( n135 & n174 ) ;
  assign n3253 = n3251 | n3252 ;
  assign n3254 = x99 & n147 ;
  assign n3255 = n3253 | n3254 ;
  assign n3256 = n3250 | n3255 ;
  assign n3257 = n3250 & n3255 ;
  assign n3258 = n3256 & ~n3257 ;
  assign n3259 = ( n3096 & ~n3245 ) | ( n3096 & n3258 ) | ( ~n3245 & n3258 ) ;
  assign n3260 = ( n3096 & n3245 ) | ( n3096 & n3258 ) | ( n3245 & n3258 ) ;
  assign n3261 = ( n3245 & n3259 ) | ( n3245 & ~n3260 ) | ( n3259 & ~n3260 ) ;
  assign n3262 = ( ~x99 & x100 ) | ( ~x99 & n3247 ) | ( x100 & n3247 ) ;
  assign n3263 = ( x99 & x100 ) | ( x99 & n3247 ) | ( x100 & n3247 ) ;
  assign n3264 = ( x99 & n3262 ) | ( x99 & ~n3263 ) | ( n3262 & ~n3263 ) ;
  assign n3265 = x0 & n3264 ;
  assign n3266 = ( x1 & x2 ) | ( x1 & n3265 ) | ( x2 & n3265 ) ;
  assign n3267 = x99 & n172 ;
  assign n3268 = ( ~x98 & n135 ) | ( ~x98 & n174 ) | ( n135 & n174 ) ;
  assign n3269 = n3267 | n3268 ;
  assign n3270 = x100 & n147 ;
  assign n3271 = n3269 | n3270 ;
  assign n3272 = n3266 | n3271 ;
  assign n3273 = n3266 & n3271 ;
  assign n3274 = n3272 & ~n3273 ;
  assign n3275 = n206 & n2788 ;
  assign n3276 = x5 & n3275 ;
  assign n3277 = x97 & n205 ;
  assign n3278 = x96 & n201 ;
  assign n3279 = n3277 | n3278 ;
  assign n3280 = x95 & n221 ;
  assign n3281 = n3279 | n3280 ;
  assign n3282 = ( ~x5 & n3275 ) | ( ~x5 & n3281 ) | ( n3275 & n3281 ) ;
  assign n3283 = x5 & ~n3281 ;
  assign n3284 = ( ~n3276 & n3282 ) | ( ~n3276 & n3283 ) | ( n3282 & n3283 ) ;
  assign n3285 = n449 & n1959 ;
  assign n3286 = x11 & n3285 ;
  assign n3287 = x91 & n456 ;
  assign n3288 = x90 & n453 ;
  assign n3289 = n3287 | n3288 ;
  assign n3290 = x89 & n536 ;
  assign n3291 = n3289 | n3290 ;
  assign n3292 = ( ~x11 & n3285 ) | ( ~x11 & n3291 ) | ( n3285 & n3291 ) ;
  assign n3293 = x11 & ~n3291 ;
  assign n3294 = ( ~n3286 & n3292 ) | ( ~n3286 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3295 = n874 & n1368 ;
  assign n3296 = x17 & n3295 ;
  assign n3297 = x85 & n881 ;
  assign n3298 = x84 & n878 ;
  assign n3299 = n3297 | n3298 ;
  assign n3300 = x83 & n959 ;
  assign n3301 = n3299 | n3300 ;
  assign n3302 = ( ~x17 & n3295 ) | ( ~x17 & n3301 ) | ( n3295 & n3301 ) ;
  assign n3303 = x17 & ~n3301 ;
  assign n3304 = ( ~n3296 & n3302 ) | ( ~n3296 & n3303 ) | ( n3302 & n3303 ) ;
  assign n3305 = n1006 & n1146 ;
  assign n3306 = x20 & n3305 ;
  assign n3307 = x82 & n1153 ;
  assign n3308 = x81 & n1150 ;
  assign n3309 = n3307 | n3308 ;
  assign n3310 = x80 & n1217 ;
  assign n3311 = n3309 | n3310 ;
  assign n3312 = ( ~x20 & n3305 ) | ( ~x20 & n3311 ) | ( n3305 & n3311 ) ;
  assign n3313 = x20 & ~n3311 ;
  assign n3314 = ( ~n3306 & n3312 ) | ( ~n3306 & n3313 ) | ( n3312 & n3313 ) ;
  assign n3315 = ( n3007 & n3148 ) | ( n3007 & ~n3165 ) | ( n3148 & ~n3165 ) ;
  assign n3316 = ( n3007 & n3148 ) | ( n3007 & n3165 ) | ( n3148 & n3165 ) ;
  assign n3317 = ( n3165 & n3315 ) | ( n3165 & ~n3316 ) | ( n3315 & ~n3316 ) ;
  assign n3318 = ( n3009 & n3138 ) | ( n3009 & n3317 ) | ( n3138 & n3317 ) ;
  assign n3319 = n388 & n2137 ;
  assign n3320 = x29 & n3319 ;
  assign n3321 = x73 & n2144 ;
  assign n3322 = x72 & n2141 ;
  assign n3323 = n3321 | n3322 ;
  assign n3324 = x71 & n2267 ;
  assign n3325 = n3323 | n3324 ;
  assign n3326 = ( ~x29 & n3319 ) | ( ~x29 & n3325 ) | ( n3319 & n3325 ) ;
  assign n3327 = x29 & ~n3325 ;
  assign n3328 = ( ~n3320 & n3326 ) | ( ~n3320 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3329 = n276 & n2545 ;
  assign n3330 = x32 & n3329 ;
  assign n3331 = x70 & n2552 ;
  assign n3332 = x69 & n2549 ;
  assign n3333 = n3331 | n3332 ;
  assign n3334 = x68 & n2696 ;
  assign n3335 = n3333 | n3334 ;
  assign n3336 = ( ~x32 & n3329 ) | ( ~x32 & n3335 ) | ( n3329 & n3335 ) ;
  assign n3337 = x32 & ~n3335 ;
  assign n3338 = ( ~n3330 & n3336 ) | ( ~n3330 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3339 = n2992 | n3161 ;
  assign n3340 = x35 & n3339 ;
  assign n3341 = x67 & n2989 ;
  assign n3342 = x66 & n2986 ;
  assign n3343 = x65 & n3159 ;
  assign n3344 = n3342 | n3343 ;
  assign n3345 = n3341 | n3344 ;
  assign n3346 = n169 & n2982 ;
  assign n3347 = n3345 | n3346 ;
  assign n3348 = x35 | x36 ;
  assign n3349 = x35 & x36 ;
  assign n3350 = n3348 & ~n3349 ;
  assign n3351 = x64 & n3350 ;
  assign n3352 = ( n3340 & ~n3347 ) | ( n3340 & n3351 ) | ( ~n3347 & n3351 ) ;
  assign n3353 = x35 & ~n3347 ;
  assign n3354 = ( ~n3340 & n3347 ) | ( ~n3340 & n3353 ) | ( n3347 & n3353 ) ;
  assign n3355 = ( n3351 & n3353 ) | ( n3351 & n3354 ) | ( n3353 & n3354 ) ;
  assign n3356 = ( n3352 & n3354 ) | ( n3352 & ~n3355 ) | ( n3354 & ~n3355 ) ;
  assign n3357 = ( n3316 & n3338 ) | ( n3316 & n3356 ) | ( n3338 & n3356 ) ;
  assign n3358 = ( ~n3316 & n3338 ) | ( ~n3316 & n3356 ) | ( n3338 & n3356 ) ;
  assign n3359 = ( n3316 & ~n3357 ) | ( n3316 & n3358 ) | ( ~n3357 & n3358 ) ;
  assign n3360 = ( n3318 & n3328 ) | ( n3318 & n3359 ) | ( n3328 & n3359 ) ;
  assign n3361 = ( ~n3318 & n3328 ) | ( ~n3318 & n3359 ) | ( n3328 & n3359 ) ;
  assign n3362 = ( n3318 & ~n3360 ) | ( n3318 & n3361 ) | ( ~n3360 & n3361 ) ;
  assign n3363 = n565 & n1755 ;
  assign n3364 = x26 & n3363 ;
  assign n3365 = x76 & n1762 ;
  assign n3366 = x75 & n1759 ;
  assign n3367 = n3365 | n3366 ;
  assign n3368 = x74 & n1895 ;
  assign n3369 = n3367 | n3368 ;
  assign n3370 = ( ~x26 & n3363 ) | ( ~x26 & n3369 ) | ( n3363 & n3369 ) ;
  assign n3371 = x26 & ~n3369 ;
  assign n3372 = ( ~n3364 & n3370 ) | ( ~n3364 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3373 = ( n3182 & n3362 ) | ( n3182 & n3372 ) | ( n3362 & n3372 ) ;
  assign n3374 = ( ~n3182 & n3362 ) | ( ~n3182 & n3372 ) | ( n3362 & n3372 ) ;
  assign n3375 = ( n3182 & ~n3373 ) | ( n3182 & n3374 ) | ( ~n3373 & n3374 ) ;
  assign n3376 = n823 & n1427 ;
  assign n3377 = x23 & n3376 ;
  assign n3378 = x79 & n1434 ;
  assign n3379 = x78 & n1431 ;
  assign n3380 = n3378 | n3379 ;
  assign n3381 = x77 & n1531 ;
  assign n3382 = n3380 | n3381 ;
  assign n3383 = ( ~x23 & n3376 ) | ( ~x23 & n3382 ) | ( n3376 & n3382 ) ;
  assign n3384 = x23 & ~n3382 ;
  assign n3385 = ( ~n3377 & n3383 ) | ( ~n3377 & n3384 ) | ( n3383 & n3384 ) ;
  assign n3386 = ( n3196 & ~n3375 ) | ( n3196 & n3385 ) | ( ~n3375 & n3385 ) ;
  assign n3387 = ( n3196 & n3375 ) | ( n3196 & n3385 ) | ( n3375 & n3385 ) ;
  assign n3388 = ( n3375 & n3386 ) | ( n3375 & ~n3387 ) | ( n3386 & ~n3387 ) ;
  assign n3389 = ( n3199 & n3314 ) | ( n3199 & n3388 ) | ( n3314 & n3388 ) ;
  assign n3390 = ( ~n3199 & n3314 ) | ( ~n3199 & n3388 ) | ( n3314 & n3388 ) ;
  assign n3391 = ( n3199 & ~n3389 ) | ( n3199 & n3390 ) | ( ~n3389 & n3390 ) ;
  assign n3392 = ( ~n3212 & n3304 ) | ( ~n3212 & n3391 ) | ( n3304 & n3391 ) ;
  assign n3393 = ( n3212 & n3304 ) | ( n3212 & n3391 ) | ( n3304 & n3391 ) ;
  assign n3394 = ( n3212 & n3392 ) | ( n3212 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = n649 & n1602 ;
  assign n3396 = x14 & n3395 ;
  assign n3397 = x88 & n656 ;
  assign n3398 = x87 & n653 ;
  assign n3399 = n3397 | n3398 ;
  assign n3400 = x86 & n744 ;
  assign n3401 = n3399 | n3400 ;
  assign n3402 = ( ~x14 & n3395 ) | ( ~x14 & n3401 ) | ( n3395 & n3401 ) ;
  assign n3403 = x14 & ~n3401 ;
  assign n3404 = ( ~n3396 & n3402 ) | ( ~n3396 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3405 = ( n3225 & ~n3394 ) | ( n3225 & n3404 ) | ( ~n3394 & n3404 ) ;
  assign n3406 = ( n3225 & n3394 ) | ( n3225 & n3404 ) | ( n3394 & n3404 ) ;
  assign n3407 = ( n3394 & n3405 ) | ( n3394 & ~n3406 ) | ( n3405 & ~n3406 ) ;
  assign n3408 = ( n3228 & n3294 ) | ( n3228 & n3407 ) | ( n3294 & n3407 ) ;
  assign n3409 = ( ~n3228 & n3294 ) | ( ~n3228 & n3407 ) | ( n3294 & n3407 ) ;
  assign n3410 = ( n3228 & ~n3408 ) | ( n3228 & n3409 ) | ( ~n3408 & n3409 ) ;
  assign n3411 = n301 & n2476 ;
  assign n3412 = x8 & n3411 ;
  assign n3413 = x94 & n309 ;
  assign n3414 = x93 & n306 ;
  assign n3415 = n3413 | n3414 ;
  assign n3416 = x92 & n359 ;
  assign n3417 = n3415 | n3416 ;
  assign n3418 = ( ~x8 & n3411 ) | ( ~x8 & n3417 ) | ( n3411 & n3417 ) ;
  assign n3419 = x8 & ~n3417 ;
  assign n3420 = ( ~n3412 & n3418 ) | ( ~n3412 & n3419 ) | ( n3418 & n3419 ) ;
  assign n3421 = ( n3230 & n3410 ) | ( n3230 & n3420 ) | ( n3410 & n3420 ) ;
  assign n3422 = ( ~n3230 & n3410 ) | ( ~n3230 & n3420 ) | ( n3410 & n3420 ) ;
  assign n3423 = ( n3230 & ~n3421 ) | ( n3230 & n3422 ) | ( ~n3421 & n3422 ) ;
  assign n3424 = ( n3243 & ~n3284 ) | ( n3243 & n3423 ) | ( ~n3284 & n3423 ) ;
  assign n3425 = ( n3243 & n3284 ) | ( n3243 & n3423 ) | ( n3284 & n3423 ) ;
  assign n3426 = ( n3284 & n3424 ) | ( n3284 & ~n3425 ) | ( n3424 & ~n3425 ) ;
  assign n3427 = ( n3260 & n3274 ) | ( n3260 & n3426 ) | ( n3274 & n3426 ) ;
  assign n3428 = ( ~n3260 & n3274 ) | ( ~n3260 & n3426 ) | ( n3274 & n3426 ) ;
  assign n3429 = ( n3260 & ~n3427 ) | ( n3260 & n3428 ) | ( ~n3427 & n3428 ) ;
  assign n3430 = n206 & n2939 ;
  assign n3431 = x5 & n3430 ;
  assign n3432 = x98 & n205 ;
  assign n3433 = x97 & n201 ;
  assign n3434 = n3432 | n3433 ;
  assign n3435 = x96 & n221 ;
  assign n3436 = n3434 | n3435 ;
  assign n3437 = ( ~x5 & n3430 ) | ( ~x5 & n3436 ) | ( n3430 & n3436 ) ;
  assign n3438 = x5 & ~n3436 ;
  assign n3439 = ( ~n3431 & n3437 ) | ( ~n3431 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3440 = n301 & n2492 ;
  assign n3441 = x8 & n3440 ;
  assign n3442 = x95 & n309 ;
  assign n3443 = x94 & n306 ;
  assign n3444 = n3442 | n3443 ;
  assign n3445 = x93 & n359 ;
  assign n3446 = n3444 | n3445 ;
  assign n3447 = ( ~x8 & n3440 ) | ( ~x8 & n3446 ) | ( n3440 & n3446 ) ;
  assign n3448 = x8 & ~n3446 ;
  assign n3449 = ( ~n3441 & n3447 ) | ( ~n3441 & n3448 ) | ( n3447 & n3448 ) ;
  assign n3450 = n649 & n1822 ;
  assign n3451 = x14 & n3450 ;
  assign n3452 = x89 & n656 ;
  assign n3453 = x88 & n653 ;
  assign n3454 = n3452 | n3453 ;
  assign n3455 = x87 & n744 ;
  assign n3456 = n3454 | n3455 ;
  assign n3457 = ( ~x14 & n3450 ) | ( ~x14 & n3456 ) | ( n3450 & n3456 ) ;
  assign n3458 = x14 & ~n3456 ;
  assign n3459 = ( ~n3451 & n3457 ) | ( ~n3451 & n3458 ) | ( n3457 & n3458 ) ;
  assign n3460 = n1093 & n1146 ;
  assign n3461 = x20 & n3460 ;
  assign n3462 = x83 & n1153 ;
  assign n3463 = x82 & n1150 ;
  assign n3464 = n3462 | n3463 ;
  assign n3465 = x81 & n1217 ;
  assign n3466 = n3464 | n3465 ;
  assign n3467 = ( ~x20 & n3460 ) | ( ~x20 & n3466 ) | ( n3460 & n3466 ) ;
  assign n3468 = x20 & ~n3466 ;
  assign n3469 = ( ~n3461 & n3467 ) | ( ~n3461 & n3468 ) | ( n3467 & n3468 ) ;
  assign n3470 = n626 & n1755 ;
  assign n3471 = x26 & n3470 ;
  assign n3472 = x77 & n1762 ;
  assign n3473 = x76 & n1759 ;
  assign n3474 = n3472 | n3473 ;
  assign n3475 = x75 & n1895 ;
  assign n3476 = n3474 | n3475 ;
  assign n3477 = ( ~x26 & n3470 ) | ( ~x26 & n3476 ) | ( n3470 & n3476 ) ;
  assign n3478 = x26 & ~n3476 ;
  assign n3479 = ( ~n3471 & n3477 ) | ( ~n3471 & n3478 ) | ( n3477 & n3478 ) ;
  assign n3480 = n322 & n2545 ;
  assign n3481 = x32 & n3480 ;
  assign n3482 = x71 & n2552 ;
  assign n3483 = x70 & n2549 ;
  assign n3484 = n3482 | n3483 ;
  assign n3485 = x69 & n2696 ;
  assign n3486 = n3484 | n3485 ;
  assign n3487 = ( ~x32 & n3480 ) | ( ~x32 & n3486 ) | ( n3480 & n3486 ) ;
  assign n3488 = x32 & ~n3486 ;
  assign n3489 = ( ~n3481 & n3487 ) | ( ~n3481 & n3488 ) | ( n3487 & n3488 ) ;
  assign n3490 = ~x37 & x38 ;
  assign n3491 = x37 & ~x38 ;
  assign n3492 = ( n3350 & n3490 ) | ( n3350 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3493 = n302 & n3492 ;
  assign n3494 = ~x35 & x37 ;
  assign n3495 = x36 & x37 ;
  assign n3496 = ( n3349 & n3494 ) | ( n3349 & ~n3495 ) | ( n3494 & ~n3495 ) ;
  assign n3497 = x64 & n3496 ;
  assign n3498 = n3493 | n3497 ;
  assign n3499 = n3350 & ~n3492 ;
  assign n3500 = x65 & n3499 ;
  assign n3501 = n3498 | n3500 ;
  assign n3502 = n3351 | n3501 ;
  assign n3503 = ( x38 & n3351 ) | ( x38 & ~n3501 ) | ( n3351 & ~n3501 ) ;
  assign n3504 = x38 & ~n3501 ;
  assign n3505 = ( n3502 & ~n3503 ) | ( n3502 & n3504 ) | ( ~n3503 & n3504 ) ;
  assign n3506 = n193 & n2982 ;
  assign n3507 = x35 & n3506 ;
  assign n3508 = x68 & n2989 ;
  assign n3509 = x67 & n2986 ;
  assign n3510 = n3508 | n3509 ;
  assign n3511 = x66 & n3159 ;
  assign n3512 = n3510 | n3511 ;
  assign n3513 = ( ~x35 & n3506 ) | ( ~x35 & n3512 ) | ( n3506 & n3512 ) ;
  assign n3514 = x35 & ~n3512 ;
  assign n3515 = ( ~n3507 & n3513 ) | ( ~n3507 & n3514 ) | ( n3513 & n3514 ) ;
  assign n3516 = ( n3355 & ~n3505 ) | ( n3355 & n3515 ) | ( ~n3505 & n3515 ) ;
  assign n3517 = ( n3355 & n3505 ) | ( n3355 & n3515 ) | ( n3505 & n3515 ) ;
  assign n3518 = ( n3505 & n3516 ) | ( n3505 & ~n3517 ) | ( n3516 & ~n3517 ) ;
  assign n3519 = ( ~n3357 & n3489 ) | ( ~n3357 & n3518 ) | ( n3489 & n3518 ) ;
  assign n3520 = ( n3357 & n3489 ) | ( n3357 & n3518 ) | ( n3489 & n3518 ) ;
  assign n3521 = ( n3357 & n3519 ) | ( n3357 & ~n3520 ) | ( n3519 & ~n3520 ) ;
  assign n3522 = n436 & n2137 ;
  assign n3523 = x29 & n3522 ;
  assign n3524 = x74 & n2144 ;
  assign n3525 = x73 & n2141 ;
  assign n3526 = n3524 | n3525 ;
  assign n3527 = x72 & n2267 ;
  assign n3528 = n3526 | n3527 ;
  assign n3529 = ( ~x29 & n3522 ) | ( ~x29 & n3528 ) | ( n3522 & n3528 ) ;
  assign n3530 = x29 & ~n3528 ;
  assign n3531 = ( ~n3523 & n3529 ) | ( ~n3523 & n3530 ) | ( n3529 & n3530 ) ;
  assign n3532 = ( n3360 & ~n3521 ) | ( n3360 & n3531 ) | ( ~n3521 & n3531 ) ;
  assign n3533 = ( n3360 & n3521 ) | ( n3360 & n3531 ) | ( n3521 & n3531 ) ;
  assign n3534 = ( n3521 & n3532 ) | ( n3521 & ~n3533 ) | ( n3532 & ~n3533 ) ;
  assign n3535 = ( n3373 & n3479 ) | ( n3373 & n3534 ) | ( n3479 & n3534 ) ;
  assign n3536 = ( ~n3373 & n3479 ) | ( ~n3373 & n3534 ) | ( n3479 & n3534 ) ;
  assign n3537 = ( n3373 & ~n3535 ) | ( n3373 & n3536 ) | ( ~n3535 & n3536 ) ;
  assign n3538 = n840 & n1427 ;
  assign n3539 = x23 & n3538 ;
  assign n3540 = x80 & n1434 ;
  assign n3541 = x79 & n1431 ;
  assign n3542 = n3540 | n3541 ;
  assign n3543 = x78 & n1531 ;
  assign n3544 = n3542 | n3543 ;
  assign n3545 = ( ~x23 & n3538 ) | ( ~x23 & n3544 ) | ( n3538 & n3544 ) ;
  assign n3546 = x23 & ~n3544 ;
  assign n3547 = ( ~n3539 & n3545 ) | ( ~n3539 & n3546 ) | ( n3545 & n3546 ) ;
  assign n3548 = ( n3387 & ~n3537 ) | ( n3387 & n3547 ) | ( ~n3537 & n3547 ) ;
  assign n3549 = ( n3387 & n3537 ) | ( n3387 & n3547 ) | ( n3537 & n3547 ) ;
  assign n3550 = ( n3537 & n3548 ) | ( n3537 & ~n3549 ) | ( n3548 & ~n3549 ) ;
  assign n3551 = ( n3389 & n3469 ) | ( n3389 & n3550 ) | ( n3469 & n3550 ) ;
  assign n3552 = ( ~n3389 & n3469 ) | ( ~n3389 & n3550 ) | ( n3469 & n3550 ) ;
  assign n3553 = ( n3389 & ~n3551 ) | ( n3389 & n3552 ) | ( ~n3551 & n3552 ) ;
  assign n3554 = n874 & n1384 ;
  assign n3555 = x17 & n3554 ;
  assign n3556 = x86 & n881 ;
  assign n3557 = x85 & n878 ;
  assign n3558 = n3556 | n3557 ;
  assign n3559 = x84 & n959 ;
  assign n3560 = n3558 | n3559 ;
  assign n3561 = ( ~x17 & n3554 ) | ( ~x17 & n3560 ) | ( n3554 & n3560 ) ;
  assign n3562 = x17 & ~n3560 ;
  assign n3563 = ( ~n3555 & n3561 ) | ( ~n3555 & n3562 ) | ( n3561 & n3562 ) ;
  assign n3564 = ( n3393 & ~n3553 ) | ( n3393 & n3563 ) | ( ~n3553 & n3563 ) ;
  assign n3565 = ( n3393 & n3553 ) | ( n3393 & n3563 ) | ( n3553 & n3563 ) ;
  assign n3566 = ( n3553 & n3564 ) | ( n3553 & ~n3565 ) | ( n3564 & ~n3565 ) ;
  assign n3567 = ( n3406 & n3459 ) | ( n3406 & n3566 ) | ( n3459 & n3566 ) ;
  assign n3568 = ( ~n3406 & n3459 ) | ( ~n3406 & n3566 ) | ( n3459 & n3566 ) ;
  assign n3569 = ( n3406 & ~n3567 ) | ( n3406 & n3568 ) | ( ~n3567 & n3568 ) ;
  assign n3570 = n449 & n2083 ;
  assign n3571 = x11 & n3570 ;
  assign n3572 = x92 & n456 ;
  assign n3573 = x91 & n453 ;
  assign n3574 = n3572 | n3573 ;
  assign n3575 = x90 & n536 ;
  assign n3576 = n3574 | n3575 ;
  assign n3577 = ( ~x11 & n3570 ) | ( ~x11 & n3576 ) | ( n3570 & n3576 ) ;
  assign n3578 = x11 & ~n3576 ;
  assign n3579 = ( ~n3571 & n3577 ) | ( ~n3571 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = ( n3408 & ~n3569 ) | ( n3408 & n3579 ) | ( ~n3569 & n3579 ) ;
  assign n3581 = ( n3408 & n3569 ) | ( n3408 & n3579 ) | ( n3569 & n3579 ) ;
  assign n3582 = ( n3569 & n3580 ) | ( n3569 & ~n3581 ) | ( n3580 & ~n3581 ) ;
  assign n3583 = ( n3421 & n3449 ) | ( n3421 & n3582 ) | ( n3449 & n3582 ) ;
  assign n3584 = ( ~n3421 & n3449 ) | ( ~n3421 & n3582 ) | ( n3449 & n3582 ) ;
  assign n3585 = ( n3421 & ~n3583 ) | ( n3421 & n3584 ) | ( ~n3583 & n3584 ) ;
  assign n3586 = ( ~n3425 & n3439 ) | ( ~n3425 & n3585 ) | ( n3439 & n3585 ) ;
  assign n3587 = ( n3425 & n3439 ) | ( n3425 & n3585 ) | ( n3439 & n3585 ) ;
  assign n3588 = ( n3425 & n3586 ) | ( n3425 & ~n3587 ) | ( n3586 & ~n3587 ) ;
  assign n3589 = ( ~x100 & x101 ) | ( ~x100 & n3263 ) | ( x101 & n3263 ) ;
  assign n3590 = ( x100 & x101 ) | ( x100 & n3263 ) | ( x101 & n3263 ) ;
  assign n3591 = ( x100 & n3589 ) | ( x100 & ~n3590 ) | ( n3589 & ~n3590 ) ;
  assign n3592 = x0 & n3591 ;
  assign n3593 = ( x1 & x2 ) | ( x1 & n3592 ) | ( x2 & n3592 ) ;
  assign n3594 = x100 & n172 ;
  assign n3595 = x101 | n3594 ;
  assign n3596 = ( n147 & n3594 ) | ( n147 & n3595 ) | ( n3594 & n3595 ) ;
  assign n3597 = ( ~x99 & n135 ) | ( ~x99 & n174 ) | ( n135 & n174 ) ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3593 | n3598 ;
  assign n3600 = n3593 & n3598 ;
  assign n3601 = n3599 & ~n3600 ;
  assign n3602 = ( n3427 & ~n3588 ) | ( n3427 & n3601 ) | ( ~n3588 & n3601 ) ;
  assign n3603 = ( n3427 & n3588 ) | ( n3427 & n3601 ) | ( n3588 & n3601 ) ;
  assign n3604 = ( n3588 & n3602 ) | ( n3588 & ~n3603 ) | ( n3602 & ~n3603 ) ;
  assign n3605 = n206 & n3248 ;
  assign n3606 = x5 & n3605 ;
  assign n3607 = x99 & n205 ;
  assign n3608 = x98 & n201 ;
  assign n3609 = n3607 | n3608 ;
  assign n3610 = x97 & n221 ;
  assign n3611 = n3609 | n3610 ;
  assign n3612 = ( ~x5 & n3605 ) | ( ~x5 & n3611 ) | ( n3605 & n3611 ) ;
  assign n3613 = x5 & ~n3611 ;
  assign n3614 = ( ~n3606 & n3612 ) | ( ~n3606 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3615 = n301 & n2772 ;
  assign n3616 = x8 & n3615 ;
  assign n3617 = x96 & n309 ;
  assign n3618 = x95 & n306 ;
  assign n3619 = n3617 | n3618 ;
  assign n3620 = x94 & n359 ;
  assign n3621 = n3619 | n3620 ;
  assign n3622 = ( ~x8 & n3615 ) | ( ~x8 & n3621 ) | ( n3615 & n3621 ) ;
  assign n3623 = x8 & ~n3621 ;
  assign n3624 = ( ~n3616 & n3622 ) | ( ~n3616 & n3623 ) | ( n3622 & n3623 ) ;
  assign n3625 = n874 & n1494 ;
  assign n3626 = x17 & n3625 ;
  assign n3627 = x87 & n881 ;
  assign n3628 = x86 & n878 ;
  assign n3629 = n3627 | n3628 ;
  assign n3630 = x85 & n959 ;
  assign n3631 = n3629 | n3630 ;
  assign n3632 = ( ~x17 & n3625 ) | ( ~x17 & n3631 ) | ( n3625 & n3631 ) ;
  assign n3633 = x17 & ~n3631 ;
  assign n3634 = ( ~n3626 & n3632 ) | ( ~n3626 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3635 = n990 & n1427 ;
  assign n3636 = x23 & n3635 ;
  assign n3637 = x81 & n1434 ;
  assign n3638 = x80 & n1431 ;
  assign n3639 = n3637 | n3638 ;
  assign n3640 = x79 & n1531 ;
  assign n3641 = n3639 | n3640 ;
  assign n3642 = ( ~x23 & n3635 ) | ( ~x23 & n3641 ) | ( n3635 & n3641 ) ;
  assign n3643 = x23 & ~n3641 ;
  assign n3644 = ( ~n3636 & n3642 ) | ( ~n3636 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3645 = n508 & n2137 ;
  assign n3646 = x29 & n3645 ;
  assign n3647 = x75 & n2144 ;
  assign n3648 = x74 & n2141 ;
  assign n3649 = n3647 | n3648 ;
  assign n3650 = x73 & n2267 ;
  assign n3651 = n3649 | n3650 ;
  assign n3652 = ( ~x29 & n3645 ) | ( ~x29 & n3651 ) | ( n3645 & n3651 ) ;
  assign n3653 = x29 & ~n3651 ;
  assign n3654 = ( ~n3646 & n3652 ) | ( ~n3646 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = x66 & n3499 ;
  assign n3656 = x65 & n3496 ;
  assign n3657 = n3655 | n3656 ;
  assign n3658 = n226 & n3492 ;
  assign n3659 = n3657 | n3658 ;
  assign n3660 = n3349 & n3491 ;
  assign n3661 = ~n3348 & n3490 ;
  assign n3662 = n3660 | n3661 ;
  assign n3663 = x64 & n3662 ;
  assign n3664 = n3659 | n3663 ;
  assign n3665 = ~x38 & n3664 ;
  assign n3666 = ( x38 & n3502 ) | ( x38 & n3664 ) | ( n3502 & n3664 ) ;
  assign n3667 = n3502 & n3664 ;
  assign n3668 = ( n3665 & n3666 ) | ( n3665 & ~n3667 ) | ( n3666 & ~n3667 ) ;
  assign n3669 = n240 & n2982 ;
  assign n3670 = x35 & n3669 ;
  assign n3671 = x69 & n2989 ;
  assign n3672 = x68 & n2986 ;
  assign n3673 = n3671 | n3672 ;
  assign n3674 = x67 & n3159 ;
  assign n3675 = n3673 | n3674 ;
  assign n3676 = ( ~x35 & n3669 ) | ( ~x35 & n3675 ) | ( n3669 & n3675 ) ;
  assign n3677 = x35 & ~n3675 ;
  assign n3678 = ( ~n3670 & n3676 ) | ( ~n3670 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3679 = ( n3517 & n3668 ) | ( n3517 & n3678 ) | ( n3668 & n3678 ) ;
  assign n3680 = ( ~n3517 & n3668 ) | ( ~n3517 & n3678 ) | ( n3668 & n3678 ) ;
  assign n3681 = ( n3517 & ~n3679 ) | ( n3517 & n3680 ) | ( ~n3679 & n3680 ) ;
  assign n3682 = n372 & n2545 ;
  assign n3683 = x32 & n3682 ;
  assign n3684 = x72 & n2552 ;
  assign n3685 = x71 & n2549 ;
  assign n3686 = n3684 | n3685 ;
  assign n3687 = x70 & n2696 ;
  assign n3688 = n3686 | n3687 ;
  assign n3689 = ( ~x32 & n3682 ) | ( ~x32 & n3688 ) | ( n3682 & n3688 ) ;
  assign n3690 = x32 & ~n3688 ;
  assign n3691 = ( ~n3683 & n3689 ) | ( ~n3683 & n3690 ) | ( n3689 & n3690 ) ;
  assign n3692 = ( n3520 & ~n3681 ) | ( n3520 & n3691 ) | ( ~n3681 & n3691 ) ;
  assign n3693 = ( n3520 & n3681 ) | ( n3520 & n3691 ) | ( n3681 & n3691 ) ;
  assign n3694 = ( n3681 & n3692 ) | ( n3681 & ~n3693 ) | ( n3692 & ~n3693 ) ;
  assign n3695 = ( n3533 & n3654 ) | ( n3533 & n3694 ) | ( n3654 & n3694 ) ;
  assign n3696 = ( ~n3533 & n3654 ) | ( ~n3533 & n3694 ) | ( n3654 & n3694 ) ;
  assign n3697 = ( n3533 & ~n3695 ) | ( n3533 & n3696 ) | ( ~n3695 & n3696 ) ;
  assign n3698 = n697 & n1755 ;
  assign n3699 = x26 & n3698 ;
  assign n3700 = x78 & n1762 ;
  assign n3701 = x77 & n1759 ;
  assign n3702 = n3700 | n3701 ;
  assign n3703 = x76 & n1895 ;
  assign n3704 = n3702 | n3703 ;
  assign n3705 = ( ~x26 & n3698 ) | ( ~x26 & n3704 ) | ( n3698 & n3704 ) ;
  assign n3706 = x26 & ~n3704 ;
  assign n3707 = ( ~n3699 & n3705 ) | ( ~n3699 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3708 = ( n3535 & ~n3697 ) | ( n3535 & n3707 ) | ( ~n3697 & n3707 ) ;
  assign n3709 = ( n3535 & n3697 ) | ( n3535 & n3707 ) | ( n3697 & n3707 ) ;
  assign n3710 = ( n3697 & n3708 ) | ( n3697 & ~n3709 ) | ( n3708 & ~n3709 ) ;
  assign n3711 = ( ~n3549 & n3644 ) | ( ~n3549 & n3710 ) | ( n3644 & n3710 ) ;
  assign n3712 = ( n3549 & n3644 ) | ( n3549 & n3710 ) | ( n3644 & n3710 ) ;
  assign n3713 = ( n3549 & n3711 ) | ( n3549 & ~n3712 ) | ( n3711 & ~n3712 ) ;
  assign n3714 = n1146 & n1190 ;
  assign n3715 = x20 & n3714 ;
  assign n3716 = x83 & n1150 ;
  assign n3717 = x82 & n1217 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = x84 & n1153 ;
  assign n3720 = n3718 | n3719 ;
  assign n3721 = ( ~x20 & n3714 ) | ( ~x20 & n3720 ) | ( n3714 & n3720 ) ;
  assign n3722 = x20 & ~n3720 ;
  assign n3723 = ( ~n3715 & n3721 ) | ( ~n3715 & n3722 ) | ( n3721 & n3722 ) ;
  assign n3724 = ( n3551 & ~n3713 ) | ( n3551 & n3723 ) | ( ~n3713 & n3723 ) ;
  assign n3725 = ( n3551 & n3713 ) | ( n3551 & n3723 ) | ( n3713 & n3723 ) ;
  assign n3726 = ( n3713 & n3724 ) | ( n3713 & ~n3725 ) | ( n3724 & ~n3725 ) ;
  assign n3727 = ( ~n3565 & n3634 ) | ( ~n3565 & n3726 ) | ( n3634 & n3726 ) ;
  assign n3728 = ( n3565 & n3634 ) | ( n3565 & n3726 ) | ( n3634 & n3726 ) ;
  assign n3729 = ( n3565 & n3727 ) | ( n3565 & ~n3728 ) | ( n3727 & ~n3728 ) ;
  assign n3730 = n649 & n1838 ;
  assign n3731 = x14 & n3730 ;
  assign n3732 = x90 & n656 ;
  assign n3733 = x89 & n653 ;
  assign n3734 = n3732 | n3733 ;
  assign n3735 = x88 & n744 ;
  assign n3736 = n3734 | n3735 ;
  assign n3737 = ( ~x14 & n3730 ) | ( ~x14 & n3736 ) | ( n3730 & n3736 ) ;
  assign n3738 = x14 & ~n3736 ;
  assign n3739 = ( ~n3731 & n3737 ) | ( ~n3731 & n3738 ) | ( n3737 & n3738 ) ;
  assign n3740 = ( n3567 & ~n3729 ) | ( n3567 & n3739 ) | ( ~n3729 & n3739 ) ;
  assign n3741 = ( n3567 & n3729 ) | ( n3567 & n3739 ) | ( n3729 & n3739 ) ;
  assign n3742 = ( n3729 & n3740 ) | ( n3729 & ~n3741 ) | ( n3740 & ~n3741 ) ;
  assign n3743 = n449 & n2220 ;
  assign n3744 = x11 & n3743 ;
  assign n3745 = x93 & n456 ;
  assign n3746 = x92 & n453 ;
  assign n3747 = n3745 | n3746 ;
  assign n3748 = x91 & n536 ;
  assign n3749 = n3747 | n3748 ;
  assign n3750 = ( ~x11 & n3743 ) | ( ~x11 & n3749 ) | ( n3743 & n3749 ) ;
  assign n3751 = x11 & ~n3749 ;
  assign n3752 = ( ~n3744 & n3750 ) | ( ~n3744 & n3751 ) | ( n3750 & n3751 ) ;
  assign n3753 = ( n3581 & ~n3742 ) | ( n3581 & n3752 ) | ( ~n3742 & n3752 ) ;
  assign n3754 = ( n3581 & n3742 ) | ( n3581 & n3752 ) | ( n3742 & n3752 ) ;
  assign n3755 = ( n3742 & n3753 ) | ( n3742 & ~n3754 ) | ( n3753 & ~n3754 ) ;
  assign n3756 = ( n3583 & n3624 ) | ( n3583 & n3755 ) | ( n3624 & n3755 ) ;
  assign n3757 = ( ~n3583 & n3624 ) | ( ~n3583 & n3755 ) | ( n3624 & n3755 ) ;
  assign n3758 = ( n3583 & ~n3756 ) | ( n3583 & n3757 ) | ( ~n3756 & n3757 ) ;
  assign n3759 = ( n3587 & n3614 ) | ( n3587 & n3758 ) | ( n3614 & n3758 ) ;
  assign n3760 = ( ~n3587 & n3614 ) | ( ~n3587 & n3758 ) | ( n3614 & n3758 ) ;
  assign n3761 = ( n3587 & ~n3759 ) | ( n3587 & n3760 ) | ( ~n3759 & n3760 ) ;
  assign n3762 = ( ~x101 & x102 ) | ( ~x101 & n3590 ) | ( x102 & n3590 ) ;
  assign n3763 = ( x101 & x102 ) | ( x101 & n3590 ) | ( x102 & n3590 ) ;
  assign n3764 = ( x101 & n3762 ) | ( x101 & ~n3763 ) | ( n3762 & ~n3763 ) ;
  assign n3765 = x0 & n3764 ;
  assign n3766 = ( x1 & x2 ) | ( x1 & n3765 ) | ( x2 & n3765 ) ;
  assign n3767 = x101 & n172 ;
  assign n3768 = x102 | n3767 ;
  assign n3769 = ( n147 & n3767 ) | ( n147 & n3768 ) | ( n3767 & n3768 ) ;
  assign n3770 = ( ~x100 & n135 ) | ( ~x100 & n174 ) | ( n135 & n174 ) ;
  assign n3771 = n3769 | n3770 ;
  assign n3772 = n3766 | n3771 ;
  assign n3773 = n3766 & n3771 ;
  assign n3774 = n3772 & ~n3773 ;
  assign n3775 = ( n3603 & n3761 ) | ( n3603 & n3774 ) | ( n3761 & n3774 ) ;
  assign n3776 = ( ~n3603 & n3761 ) | ( ~n3603 & n3774 ) | ( n3761 & n3774 ) ;
  assign n3777 = ( n3603 & ~n3775 ) | ( n3603 & n3776 ) | ( ~n3775 & n3776 ) ;
  assign n3778 = n301 & n2788 ;
  assign n3779 = x8 & n3778 ;
  assign n3780 = x97 & n309 ;
  assign n3781 = x96 & n306 ;
  assign n3782 = n3780 | n3781 ;
  assign n3783 = x95 & n359 ;
  assign n3784 = n3782 | n3783 ;
  assign n3785 = ( ~x8 & n3778 ) | ( ~x8 & n3784 ) | ( n3778 & n3784 ) ;
  assign n3786 = x8 & ~n3784 ;
  assign n3787 = ( ~n3779 & n3785 ) | ( ~n3779 & n3786 ) | ( n3785 & n3786 ) ;
  assign n3788 = n649 & n1959 ;
  assign n3789 = x14 & n3788 ;
  assign n3790 = x91 & n656 ;
  assign n3791 = x90 & n653 ;
  assign n3792 = n3790 | n3791 ;
  assign n3793 = x89 & n744 ;
  assign n3794 = n3792 | n3793 ;
  assign n3795 = ( ~x14 & n3788 ) | ( ~x14 & n3794 ) | ( n3788 & n3794 ) ;
  assign n3796 = x14 & ~n3794 ;
  assign n3797 = ( ~n3789 & n3795 ) | ( ~n3789 & n3796 ) | ( n3795 & n3796 ) ;
  assign n3798 = n1146 & n1368 ;
  assign n3799 = x20 & n3798 ;
  assign n3800 = x85 & n1153 ;
  assign n3801 = x84 & n1150 ;
  assign n3802 = n3800 | n3801 ;
  assign n3803 = x83 & n1217 ;
  assign n3804 = n3802 | n3803 ;
  assign n3805 = ( ~x20 & n3798 ) | ( ~x20 & n3804 ) | ( n3798 & n3804 ) ;
  assign n3806 = x20 & ~n3804 ;
  assign n3807 = ( ~n3799 & n3805 ) | ( ~n3799 & n3806 ) | ( n3805 & n3806 ) ;
  assign n3808 = n823 & n1755 ;
  assign n3809 = x26 & n3808 ;
  assign n3810 = x79 & n1762 ;
  assign n3811 = x78 & n1759 ;
  assign n3812 = n3810 | n3811 ;
  assign n3813 = x77 & n1895 ;
  assign n3814 = n3812 | n3813 ;
  assign n3815 = ( ~x26 & n3808 ) | ( ~x26 & n3814 ) | ( n3808 & n3814 ) ;
  assign n3816 = x26 & ~n3814 ;
  assign n3817 = ( ~n3809 & n3815 ) | ( ~n3809 & n3816 ) | ( n3815 & n3816 ) ;
  assign n3818 = n565 & n2137 ;
  assign n3819 = x29 & n3818 ;
  assign n3820 = x76 & n2144 ;
  assign n3821 = x75 & n2141 ;
  assign n3822 = n3820 | n3821 ;
  assign n3823 = x74 & n2267 ;
  assign n3824 = n3822 | n3823 ;
  assign n3825 = ( ~x29 & n3818 ) | ( ~x29 & n3824 ) | ( n3818 & n3824 ) ;
  assign n3826 = x29 & ~n3824 ;
  assign n3827 = ( ~n3819 & n3825 ) | ( ~n3819 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3828 = n276 & n2982 ;
  assign n3829 = x35 & n3828 ;
  assign n3830 = x70 & n2989 ;
  assign n3831 = x69 & n2986 ;
  assign n3832 = n3830 | n3831 ;
  assign n3833 = x68 & n3159 ;
  assign n3834 = n3832 | n3833 ;
  assign n3835 = ( ~x35 & n3828 ) | ( ~x35 & n3834 ) | ( n3828 & n3834 ) ;
  assign n3836 = x35 & ~n3834 ;
  assign n3837 = ( ~n3829 & n3835 ) | ( ~n3829 & n3836 ) | ( n3835 & n3836 ) ;
  assign n3838 = n3502 | n3664 ;
  assign n3839 = x38 & n3838 ;
  assign n3840 = x66 & n3496 ;
  assign n3841 = x67 & n3499 ;
  assign n3842 = x65 & n3662 ;
  assign n3843 = n3841 | n3842 ;
  assign n3844 = n169 & n3492 ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = n3840 | n3845 ;
  assign n3847 = x38 | x39 ;
  assign n3848 = x38 & x39 ;
  assign n3849 = n3847 & ~n3848 ;
  assign n3850 = x64 & n3849 ;
  assign n3851 = ( n3839 & ~n3846 ) | ( n3839 & n3850 ) | ( ~n3846 & n3850 ) ;
  assign n3852 = x38 & ~n3846 ;
  assign n3853 = ( ~n3839 & n3846 ) | ( ~n3839 & n3852 ) | ( n3846 & n3852 ) ;
  assign n3854 = ( n3850 & n3852 ) | ( n3850 & n3853 ) | ( n3852 & n3853 ) ;
  assign n3855 = ( n3851 & n3853 ) | ( n3851 & ~n3854 ) | ( n3853 & ~n3854 ) ;
  assign n3856 = ( n3679 & n3837 ) | ( n3679 & n3855 ) | ( n3837 & n3855 ) ;
  assign n3857 = ( ~n3679 & n3837 ) | ( ~n3679 & n3855 ) | ( n3837 & n3855 ) ;
  assign n3858 = ( n3679 & ~n3856 ) | ( n3679 & n3857 ) | ( ~n3856 & n3857 ) ;
  assign n3859 = n388 & n2545 ;
  assign n3860 = x32 & n3859 ;
  assign n3861 = x73 & n2552 ;
  assign n3862 = x72 & n2549 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = x71 & n2696 ;
  assign n3865 = n3863 | n3864 ;
  assign n3866 = ( ~x32 & n3859 ) | ( ~x32 & n3865 ) | ( n3859 & n3865 ) ;
  assign n3867 = x32 & ~n3865 ;
  assign n3868 = ( ~n3860 & n3866 ) | ( ~n3860 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = ( n3693 & ~n3858 ) | ( n3693 & n3868 ) | ( ~n3858 & n3868 ) ;
  assign n3870 = ( n3693 & n3858 ) | ( n3693 & n3868 ) | ( n3858 & n3868 ) ;
  assign n3871 = ( n3858 & n3869 ) | ( n3858 & ~n3870 ) | ( n3869 & ~n3870 ) ;
  assign n3872 = ( n3695 & n3827 ) | ( n3695 & n3871 ) | ( n3827 & n3871 ) ;
  assign n3873 = ( ~n3695 & n3827 ) | ( ~n3695 & n3871 ) | ( n3827 & n3871 ) ;
  assign n3874 = ( n3695 & ~n3872 ) | ( n3695 & n3873 ) | ( ~n3872 & n3873 ) ;
  assign n3875 = ( n3709 & n3817 ) | ( n3709 & n3874 ) | ( n3817 & n3874 ) ;
  assign n3876 = ( ~n3709 & n3817 ) | ( ~n3709 & n3874 ) | ( n3817 & n3874 ) ;
  assign n3877 = ( n3709 & ~n3875 ) | ( n3709 & n3876 ) | ( ~n3875 & n3876 ) ;
  assign n3878 = n1006 & n1427 ;
  assign n3879 = x23 & n3878 ;
  assign n3880 = x82 & n1434 ;
  assign n3881 = x81 & n1431 ;
  assign n3882 = n3880 | n3881 ;
  assign n3883 = x80 & n1531 ;
  assign n3884 = n3882 | n3883 ;
  assign n3885 = ( ~x23 & n3878 ) | ( ~x23 & n3884 ) | ( n3878 & n3884 ) ;
  assign n3886 = x23 & ~n3884 ;
  assign n3887 = ( ~n3879 & n3885 ) | ( ~n3879 & n3886 ) | ( n3885 & n3886 ) ;
  assign n3888 = ( n3712 & ~n3877 ) | ( n3712 & n3887 ) | ( ~n3877 & n3887 ) ;
  assign n3889 = ( n3712 & n3877 ) | ( n3712 & n3887 ) | ( n3877 & n3887 ) ;
  assign n3890 = ( n3877 & n3888 ) | ( n3877 & ~n3889 ) | ( n3888 & ~n3889 ) ;
  assign n3891 = ( n3725 & n3807 ) | ( n3725 & n3890 ) | ( n3807 & n3890 ) ;
  assign n3892 = ( ~n3725 & n3807 ) | ( ~n3725 & n3890 ) | ( n3807 & n3890 ) ;
  assign n3893 = ( n3725 & ~n3891 ) | ( n3725 & n3892 ) | ( ~n3891 & n3892 ) ;
  assign n3894 = n874 & n1602 ;
  assign n3895 = x17 & n3894 ;
  assign n3896 = x88 & n881 ;
  assign n3897 = x87 & n878 ;
  assign n3898 = n3896 | n3897 ;
  assign n3899 = x86 & n959 ;
  assign n3900 = n3898 | n3899 ;
  assign n3901 = ( ~x17 & n3894 ) | ( ~x17 & n3900 ) | ( n3894 & n3900 ) ;
  assign n3902 = x17 & ~n3900 ;
  assign n3903 = ( ~n3895 & n3901 ) | ( ~n3895 & n3902 ) | ( n3901 & n3902 ) ;
  assign n3904 = ( n3728 & ~n3893 ) | ( n3728 & n3903 ) | ( ~n3893 & n3903 ) ;
  assign n3905 = ( n3728 & n3893 ) | ( n3728 & n3903 ) | ( n3893 & n3903 ) ;
  assign n3906 = ( n3893 & n3904 ) | ( n3893 & ~n3905 ) | ( n3904 & ~n3905 ) ;
  assign n3907 = ( n3741 & n3797 ) | ( n3741 & n3906 ) | ( n3797 & n3906 ) ;
  assign n3908 = ( ~n3741 & n3797 ) | ( ~n3741 & n3906 ) | ( n3797 & n3906 ) ;
  assign n3909 = ( n3741 & ~n3907 ) | ( n3741 & n3908 ) | ( ~n3907 & n3908 ) ;
  assign n3910 = n449 & n2476 ;
  assign n3911 = x11 & n3910 ;
  assign n3912 = x94 & n456 ;
  assign n3913 = x93 & n453 ;
  assign n3914 = n3912 | n3913 ;
  assign n3915 = x92 & n536 ;
  assign n3916 = n3914 | n3915 ;
  assign n3917 = ( ~x11 & n3910 ) | ( ~x11 & n3916 ) | ( n3910 & n3916 ) ;
  assign n3918 = x11 & ~n3916 ;
  assign n3919 = ( ~n3911 & n3917 ) | ( ~n3911 & n3918 ) | ( n3917 & n3918 ) ;
  assign n3920 = ( n3754 & ~n3909 ) | ( n3754 & n3919 ) | ( ~n3909 & n3919 ) ;
  assign n3921 = ( n3754 & n3909 ) | ( n3754 & n3919 ) | ( n3909 & n3919 ) ;
  assign n3922 = ( n3909 & n3920 ) | ( n3909 & ~n3921 ) | ( n3920 & ~n3921 ) ;
  assign n3923 = ( n3756 & n3787 ) | ( n3756 & n3922 ) | ( n3787 & n3922 ) ;
  assign n3924 = ( ~n3756 & n3787 ) | ( ~n3756 & n3922 ) | ( n3787 & n3922 ) ;
  assign n3925 = ( n3756 & ~n3923 ) | ( n3756 & n3924 ) | ( ~n3923 & n3924 ) ;
  assign n3926 = n206 & n3264 ;
  assign n3927 = x5 & n3926 ;
  assign n3928 = x100 & n205 ;
  assign n3929 = x99 & n201 ;
  assign n3930 = n3928 | n3929 ;
  assign n3931 = x98 & n221 ;
  assign n3932 = n3930 | n3931 ;
  assign n3933 = ( ~x5 & n3926 ) | ( ~x5 & n3932 ) | ( n3926 & n3932 ) ;
  assign n3934 = x5 & ~n3932 ;
  assign n3935 = ( ~n3927 & n3933 ) | ( ~n3927 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3936 = ( ~n3759 & n3925 ) | ( ~n3759 & n3935 ) | ( n3925 & n3935 ) ;
  assign n3937 = ( n3759 & n3925 ) | ( n3759 & n3935 ) | ( n3925 & n3935 ) ;
  assign n3938 = ( n3759 & n3936 ) | ( n3759 & ~n3937 ) | ( n3936 & ~n3937 ) ;
  assign n3939 = ( ~x102 & x103 ) | ( ~x102 & n3763 ) | ( x103 & n3763 ) ;
  assign n3940 = ( x102 & x103 ) | ( x102 & n3763 ) | ( x103 & n3763 ) ;
  assign n3941 = ( x102 & n3939 ) | ( x102 & ~n3940 ) | ( n3939 & ~n3940 ) ;
  assign n3942 = x0 & n3941 ;
  assign n3943 = ( x1 & x2 ) | ( x1 & n3942 ) | ( x2 & n3942 ) ;
  assign n3944 = x102 & n172 ;
  assign n3945 = x103 | n3944 ;
  assign n3946 = ( n147 & n3944 ) | ( n147 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3947 = ( ~x101 & n135 ) | ( ~x101 & n174 ) | ( n135 & n174 ) ;
  assign n3948 = n3946 | n3947 ;
  assign n3949 = n3943 | n3948 ;
  assign n3950 = n3943 & n3948 ;
  assign n3951 = n3949 & ~n3950 ;
  assign n3952 = ( n3775 & ~n3938 ) | ( n3775 & n3951 ) | ( ~n3938 & n3951 ) ;
  assign n3953 = ( n3775 & n3938 ) | ( n3775 & n3951 ) | ( n3938 & n3951 ) ;
  assign n3954 = ( n3938 & n3952 ) | ( n3938 & ~n3953 ) | ( n3952 & ~n3953 ) ;
  assign n3955 = ( ~x103 & x104 ) | ( ~x103 & n3940 ) | ( x104 & n3940 ) ;
  assign n3956 = ( x103 & x104 ) | ( x103 & n3940 ) | ( x104 & n3940 ) ;
  assign n3957 = ( x103 & n3955 ) | ( x103 & ~n3956 ) | ( n3955 & ~n3956 ) ;
  assign n3958 = x0 & n3957 ;
  assign n3959 = ( x1 & x2 ) | ( x1 & n3958 ) | ( x2 & n3958 ) ;
  assign n3960 = x103 & n172 ;
  assign n3961 = ( ~x102 & n135 ) | ( ~x102 & n174 ) | ( n135 & n174 ) ;
  assign n3962 = n3960 | n3961 ;
  assign n3963 = x104 & n147 ;
  assign n3964 = n3962 | n3963 ;
  assign n3965 = n3959 | n3964 ;
  assign n3966 = n3959 & n3964 ;
  assign n3967 = n3965 & ~n3966 ;
  assign n3968 = n301 & n2939 ;
  assign n3969 = x8 & n3968 ;
  assign n3970 = x98 & n309 ;
  assign n3971 = x97 & n306 ;
  assign n3972 = n3970 | n3971 ;
  assign n3973 = x96 & n359 ;
  assign n3974 = n3972 | n3973 ;
  assign n3975 = ( ~x8 & n3968 ) | ( ~x8 & n3974 ) | ( n3968 & n3974 ) ;
  assign n3976 = x8 & ~n3974 ;
  assign n3977 = ( ~n3969 & n3975 ) | ( ~n3969 & n3976 ) | ( n3975 & n3976 ) ;
  assign n3978 = n874 & n1822 ;
  assign n3979 = x17 & n3978 ;
  assign n3980 = x89 & n881 ;
  assign n3981 = x88 & n878 ;
  assign n3982 = n3980 | n3981 ;
  assign n3983 = x87 & n959 ;
  assign n3984 = n3982 | n3983 ;
  assign n3985 = ( ~x17 & n3978 ) | ( ~x17 & n3984 ) | ( n3978 & n3984 ) ;
  assign n3986 = x17 & ~n3984 ;
  assign n3987 = ( ~n3979 & n3985 ) | ( ~n3979 & n3986 ) | ( n3985 & n3986 ) ;
  assign n3988 = n1093 & n1427 ;
  assign n3989 = x23 & n3988 ;
  assign n3990 = x83 & n1434 ;
  assign n3991 = x82 & n1431 ;
  assign n3992 = n3990 | n3991 ;
  assign n3993 = x81 & n1531 ;
  assign n3994 = n3992 | n3993 ;
  assign n3995 = ( ~x23 & n3988 ) | ( ~x23 & n3994 ) | ( n3988 & n3994 ) ;
  assign n3996 = x23 & ~n3994 ;
  assign n3997 = ( ~n3989 & n3995 ) | ( ~n3989 & n3996 ) | ( n3995 & n3996 ) ;
  assign n3998 = n626 & n2137 ;
  assign n3999 = x29 & n3998 ;
  assign n4000 = x77 & n2144 ;
  assign n4001 = x76 & n2141 ;
  assign n4002 = n4000 | n4001 ;
  assign n4003 = x75 & n2267 ;
  assign n4004 = n4002 | n4003 ;
  assign n4005 = ( ~x29 & n3998 ) | ( ~x29 & n4004 ) | ( n3998 & n4004 ) ;
  assign n4006 = x29 & ~n4004 ;
  assign n4007 = ( ~n3999 & n4005 ) | ( ~n3999 & n4006 ) | ( n4005 & n4006 ) ;
  assign n4008 = n322 & n2982 ;
  assign n4009 = x35 & n4008 ;
  assign n4010 = x71 & n2989 ;
  assign n4011 = x70 & n2986 ;
  assign n4012 = n4010 | n4011 ;
  assign n4013 = x69 & n3159 ;
  assign n4014 = n4012 | n4013 ;
  assign n4015 = ( ~x35 & n4008 ) | ( ~x35 & n4014 ) | ( n4008 & n4014 ) ;
  assign n4016 = x35 & ~n4014 ;
  assign n4017 = ( ~n4009 & n4015 ) | ( ~n4009 & n4016 ) | ( n4015 & n4016 ) ;
  assign n4018 = ~x40 & x41 ;
  assign n4019 = x40 & ~x41 ;
  assign n4020 = ( n3849 & n4018 ) | ( n3849 & n4019 ) | ( n4018 & n4019 ) ;
  assign n4021 = n302 & n4020 ;
  assign n4022 = ~x38 & x40 ;
  assign n4023 = x39 & x40 ;
  assign n4024 = ( n3848 & n4022 ) | ( n3848 & ~n4023 ) | ( n4022 & ~n4023 ) ;
  assign n4025 = x64 & n4024 ;
  assign n4026 = n4021 | n4025 ;
  assign n4027 = n3849 & ~n4020 ;
  assign n4028 = x65 & n4027 ;
  assign n4029 = n4026 | n4028 ;
  assign n4030 = x41 & n3850 ;
  assign n4031 = ~n4029 & n4030 ;
  assign n4032 = n4029 & ~n4030 ;
  assign n4033 = n4031 | n4032 ;
  assign n4034 = x68 & n3499 ;
  assign n4035 = x38 & n4034 ;
  assign n4036 = x67 & n3496 ;
  assign n4037 = x66 & n3662 ;
  assign n4038 = n4036 | n4037 ;
  assign n4039 = n193 & n3492 ;
  assign n4040 = n4038 | n4039 ;
  assign n4041 = ( ~x38 & n4034 ) | ( ~x38 & n4040 ) | ( n4034 & n4040 ) ;
  assign n4042 = x38 & ~n4040 ;
  assign n4043 = ( ~n4035 & n4041 ) | ( ~n4035 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4044 = ( n3854 & ~n4033 ) | ( n3854 & n4043 ) | ( ~n4033 & n4043 ) ;
  assign n4045 = ( n3854 & n4033 ) | ( n3854 & n4043 ) | ( n4033 & n4043 ) ;
  assign n4046 = ( n4033 & n4044 ) | ( n4033 & ~n4045 ) | ( n4044 & ~n4045 ) ;
  assign n4047 = ( n3856 & n4017 ) | ( n3856 & n4046 ) | ( n4017 & n4046 ) ;
  assign n4048 = ( ~n3856 & n4017 ) | ( ~n3856 & n4046 ) | ( n4017 & n4046 ) ;
  assign n4049 = ( n3856 & ~n4047 ) | ( n3856 & n4048 ) | ( ~n4047 & n4048 ) ;
  assign n4050 = n436 & n2545 ;
  assign n4051 = x32 & n4050 ;
  assign n4052 = x74 & n2552 ;
  assign n4053 = x73 & n2549 ;
  assign n4054 = n4052 | n4053 ;
  assign n4055 = x72 & n2696 ;
  assign n4056 = n4054 | n4055 ;
  assign n4057 = ( ~x32 & n4050 ) | ( ~x32 & n4056 ) | ( n4050 & n4056 ) ;
  assign n4058 = x32 & ~n4056 ;
  assign n4059 = ( ~n4051 & n4057 ) | ( ~n4051 & n4058 ) | ( n4057 & n4058 ) ;
  assign n4060 = ( n3870 & ~n4049 ) | ( n3870 & n4059 ) | ( ~n4049 & n4059 ) ;
  assign n4061 = ( n3870 & n4049 ) | ( n3870 & n4059 ) | ( n4049 & n4059 ) ;
  assign n4062 = ( n4049 & n4060 ) | ( n4049 & ~n4061 ) | ( n4060 & ~n4061 ) ;
  assign n4063 = ( n3872 & n4007 ) | ( n3872 & n4062 ) | ( n4007 & n4062 ) ;
  assign n4064 = ( ~n3872 & n4007 ) | ( ~n3872 & n4062 ) | ( n4007 & n4062 ) ;
  assign n4065 = ( n3872 & ~n4063 ) | ( n3872 & n4064 ) | ( ~n4063 & n4064 ) ;
  assign n4066 = n840 & n1755 ;
  assign n4067 = x26 & n4066 ;
  assign n4068 = x80 & n1762 ;
  assign n4069 = x79 & n1759 ;
  assign n4070 = n4068 | n4069 ;
  assign n4071 = x78 & n1895 ;
  assign n4072 = n4070 | n4071 ;
  assign n4073 = ( ~x26 & n4066 ) | ( ~x26 & n4072 ) | ( n4066 & n4072 ) ;
  assign n4074 = x26 & ~n4072 ;
  assign n4075 = ( ~n4067 & n4073 ) | ( ~n4067 & n4074 ) | ( n4073 & n4074 ) ;
  assign n4076 = ( n3875 & ~n4065 ) | ( n3875 & n4075 ) | ( ~n4065 & n4075 ) ;
  assign n4077 = ( n3875 & n4065 ) | ( n3875 & n4075 ) | ( n4065 & n4075 ) ;
  assign n4078 = ( n4065 & n4076 ) | ( n4065 & ~n4077 ) | ( n4076 & ~n4077 ) ;
  assign n4079 = ( n3889 & n3997 ) | ( n3889 & n4078 ) | ( n3997 & n4078 ) ;
  assign n4080 = ( ~n3889 & n3997 ) | ( ~n3889 & n4078 ) | ( n3997 & n4078 ) ;
  assign n4081 = ( n3889 & ~n4079 ) | ( n3889 & n4080 ) | ( ~n4079 & n4080 ) ;
  assign n4082 = n1146 & n1384 ;
  assign n4083 = x20 & n4082 ;
  assign n4084 = x86 & n1153 ;
  assign n4085 = x85 & n1150 ;
  assign n4086 = n4084 | n4085 ;
  assign n4087 = x84 & n1217 ;
  assign n4088 = n4086 | n4087 ;
  assign n4089 = ( ~x20 & n4082 ) | ( ~x20 & n4088 ) | ( n4082 & n4088 ) ;
  assign n4090 = x20 & ~n4088 ;
  assign n4091 = ( ~n4083 & n4089 ) | ( ~n4083 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4092 = ( n3891 & ~n4081 ) | ( n3891 & n4091 ) | ( ~n4081 & n4091 ) ;
  assign n4093 = ( n3891 & n4081 ) | ( n3891 & n4091 ) | ( n4081 & n4091 ) ;
  assign n4094 = ( n4081 & n4092 ) | ( n4081 & ~n4093 ) | ( n4092 & ~n4093 ) ;
  assign n4095 = ( n3905 & n3987 ) | ( n3905 & n4094 ) | ( n3987 & n4094 ) ;
  assign n4096 = ( ~n3905 & n3987 ) | ( ~n3905 & n4094 ) | ( n3987 & n4094 ) ;
  assign n4097 = ( n3905 & ~n4095 ) | ( n3905 & n4096 ) | ( ~n4095 & n4096 ) ;
  assign n4098 = n649 & n2083 ;
  assign n4099 = x14 & n4098 ;
  assign n4100 = x92 & n656 ;
  assign n4101 = x91 & n653 ;
  assign n4102 = n4100 | n4101 ;
  assign n4103 = x90 & n744 ;
  assign n4104 = n4102 | n4103 ;
  assign n4105 = ( ~x14 & n4098 ) | ( ~x14 & n4104 ) | ( n4098 & n4104 ) ;
  assign n4106 = x14 & ~n4104 ;
  assign n4107 = ( ~n4099 & n4105 ) | ( ~n4099 & n4106 ) | ( n4105 & n4106 ) ;
  assign n4108 = ( n3907 & ~n4097 ) | ( n3907 & n4107 ) | ( ~n4097 & n4107 ) ;
  assign n4109 = ( n3907 & n4097 ) | ( n3907 & n4107 ) | ( n4097 & n4107 ) ;
  assign n4110 = ( n4097 & n4108 ) | ( n4097 & ~n4109 ) | ( n4108 & ~n4109 ) ;
  assign n4111 = n449 & n2492 ;
  assign n4112 = x11 & n4111 ;
  assign n4113 = x95 & n456 ;
  assign n4114 = x94 & n453 ;
  assign n4115 = n4113 | n4114 ;
  assign n4116 = x93 & n536 ;
  assign n4117 = n4115 | n4116 ;
  assign n4118 = ( ~x11 & n4111 ) | ( ~x11 & n4117 ) | ( n4111 & n4117 ) ;
  assign n4119 = x11 & ~n4117 ;
  assign n4120 = ( ~n4112 & n4118 ) | ( ~n4112 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4121 = ( n3921 & ~n4110 ) | ( n3921 & n4120 ) | ( ~n4110 & n4120 ) ;
  assign n4122 = ( n3921 & n4110 ) | ( n3921 & n4120 ) | ( n4110 & n4120 ) ;
  assign n4123 = ( n4110 & n4121 ) | ( n4110 & ~n4122 ) | ( n4121 & ~n4122 ) ;
  assign n4124 = ( n3923 & n3977 ) | ( n3923 & n4123 ) | ( n3977 & n4123 ) ;
  assign n4125 = ( ~n3923 & n3977 ) | ( ~n3923 & n4123 ) | ( n3977 & n4123 ) ;
  assign n4126 = ( n3923 & ~n4124 ) | ( n3923 & n4125 ) | ( ~n4124 & n4125 ) ;
  assign n4127 = n206 & n3591 ;
  assign n4128 = x5 & n4127 ;
  assign n4129 = x101 & n205 ;
  assign n4130 = x100 & n201 ;
  assign n4131 = n4129 | n4130 ;
  assign n4132 = x99 & n221 ;
  assign n4133 = n4131 | n4132 ;
  assign n4134 = ( ~x5 & n4127 ) | ( ~x5 & n4133 ) | ( n4127 & n4133 ) ;
  assign n4135 = x5 & ~n4133 ;
  assign n4136 = ( ~n4128 & n4134 ) | ( ~n4128 & n4135 ) | ( n4134 & n4135 ) ;
  assign n4137 = ( n3937 & ~n4126 ) | ( n3937 & n4136 ) | ( ~n4126 & n4136 ) ;
  assign n4138 = ( n3937 & n4126 ) | ( n3937 & n4136 ) | ( n4126 & n4136 ) ;
  assign n4139 = ( n4126 & n4137 ) | ( n4126 & ~n4138 ) | ( n4137 & ~n4138 ) ;
  assign n4140 = ( n3953 & n3967 ) | ( n3953 & n4139 ) | ( n3967 & n4139 ) ;
  assign n4141 = ( ~n3953 & n3967 ) | ( ~n3953 & n4139 ) | ( n3967 & n4139 ) ;
  assign n4142 = ( n3953 & ~n4140 ) | ( n3953 & n4141 ) | ( ~n4140 & n4141 ) ;
  assign n4143 = ( ~x104 & x105 ) | ( ~x104 & n3956 ) | ( x105 & n3956 ) ;
  assign n4144 = ( x104 & x105 ) | ( x104 & n3956 ) | ( x105 & n3956 ) ;
  assign n4145 = ( x104 & n4143 ) | ( x104 & ~n4144 ) | ( n4143 & ~n4144 ) ;
  assign n4146 = x0 & n4145 ;
  assign n4147 = ( x1 & x2 ) | ( x1 & n4146 ) | ( x2 & n4146 ) ;
  assign n4148 = x104 & n172 ;
  assign n4149 = ( ~x103 & n135 ) | ( ~x103 & n174 ) | ( n135 & n174 ) ;
  assign n4150 = n4148 | n4149 ;
  assign n4151 = x105 & n147 ;
  assign n4152 = n4150 | n4151 ;
  assign n4153 = n4147 | n4152 ;
  assign n4154 = n4147 & n4152 ;
  assign n4155 = n4153 & ~n4154 ;
  assign n4156 = n206 & n3764 ;
  assign n4157 = x5 & n4156 ;
  assign n4158 = x102 & n205 ;
  assign n4159 = x101 & n201 ;
  assign n4160 = n4158 | n4159 ;
  assign n4161 = x100 & n221 ;
  assign n4162 = n4160 | n4161 ;
  assign n4163 = ( ~x5 & n4156 ) | ( ~x5 & n4162 ) | ( n4156 & n4162 ) ;
  assign n4164 = x5 & ~n4162 ;
  assign n4165 = ( ~n4157 & n4163 ) | ( ~n4157 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4166 = n301 & n3248 ;
  assign n4167 = x8 & n4166 ;
  assign n4168 = x99 & n309 ;
  assign n4169 = x98 & n306 ;
  assign n4170 = n4168 | n4169 ;
  assign n4171 = x97 & n359 ;
  assign n4172 = n4170 | n4171 ;
  assign n4173 = ( ~x8 & n4166 ) | ( ~x8 & n4172 ) | ( n4166 & n4172 ) ;
  assign n4174 = x8 & ~n4172 ;
  assign n4175 = ( ~n4167 & n4173 ) | ( ~n4167 & n4174 ) | ( n4173 & n4174 ) ;
  assign n4176 = n449 & n2772 ;
  assign n4177 = x11 & n4176 ;
  assign n4178 = x96 & n456 ;
  assign n4179 = x95 & n453 ;
  assign n4180 = n4178 | n4179 ;
  assign n4181 = x94 & n536 ;
  assign n4182 = n4180 | n4181 ;
  assign n4183 = ( ~x11 & n4176 ) | ( ~x11 & n4182 ) | ( n4176 & n4182 ) ;
  assign n4184 = x11 & ~n4182 ;
  assign n4185 = ( ~n4177 & n4183 ) | ( ~n4177 & n4184 ) | ( n4183 & n4184 ) ;
  assign n4186 = n1146 & n1494 ;
  assign n4187 = x20 & n4186 ;
  assign n4188 = x87 & n1153 ;
  assign n4189 = x86 & n1150 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = x85 & n1217 ;
  assign n4192 = n4190 | n4191 ;
  assign n4193 = ( ~x20 & n4186 ) | ( ~x20 & n4192 ) | ( n4186 & n4192 ) ;
  assign n4194 = x20 & ~n4192 ;
  assign n4195 = ( ~n4187 & n4193 ) | ( ~n4187 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = n697 & n2137 ;
  assign n4197 = x29 & n4196 ;
  assign n4198 = x78 & n2144 ;
  assign n4199 = x77 & n2141 ;
  assign n4200 = n4198 | n4199 ;
  assign n4201 = x76 & n2267 ;
  assign n4202 = n4200 | n4201 ;
  assign n4203 = ( ~x29 & n4196 ) | ( ~x29 & n4202 ) | ( n4196 & n4202 ) ;
  assign n4204 = x29 & ~n4202 ;
  assign n4205 = ( ~n4197 & n4203 ) | ( ~n4197 & n4204 ) | ( n4203 & n4204 ) ;
  assign n4206 = n508 & n2545 ;
  assign n4207 = x32 & n4206 ;
  assign n4208 = x75 & n2552 ;
  assign n4209 = x74 & n2549 ;
  assign n4210 = n4208 | n4209 ;
  assign n4211 = x73 & n2696 ;
  assign n4212 = n4210 | n4211 ;
  assign n4213 = ( ~x32 & n4206 ) | ( ~x32 & n4212 ) | ( n4206 & n4212 ) ;
  assign n4214 = x32 & ~n4212 ;
  assign n4215 = ( ~n4207 & n4213 ) | ( ~n4207 & n4214 ) | ( n4213 & n4214 ) ;
  assign n4216 = x66 & n4027 ;
  assign n4217 = x65 & n4024 ;
  assign n4218 = n4216 | n4217 ;
  assign n4219 = n226 & n4020 ;
  assign n4220 = n4218 | n4219 ;
  assign n4221 = n3848 & n4019 ;
  assign n4222 = ~n3847 & n4018 ;
  assign n4223 = n4221 | n4222 ;
  assign n4224 = x64 & n4223 ;
  assign n4225 = n4220 | n4224 ;
  assign n4226 = ( x41 & n4029 ) | ( x41 & n4030 ) | ( n4029 & n4030 ) ;
  assign n4227 = ~n4225 & n4226 ;
  assign n4228 = n4225 & ~n4226 ;
  assign n4229 = n4227 | n4228 ;
  assign n4230 = n240 & n3492 ;
  assign n4231 = x38 & n4230 ;
  assign n4232 = x69 & n3499 ;
  assign n4233 = x68 & n3496 ;
  assign n4234 = n4232 | n4233 ;
  assign n4235 = x67 & n3662 ;
  assign n4236 = n4234 | n4235 ;
  assign n4237 = ( ~x38 & n4230 ) | ( ~x38 & n4236 ) | ( n4230 & n4236 ) ;
  assign n4238 = x38 & ~n4236 ;
  assign n4239 = ( ~n4231 & n4237 ) | ( ~n4231 & n4238 ) | ( n4237 & n4238 ) ;
  assign n4240 = ( n4045 & n4229 ) | ( n4045 & n4239 ) | ( n4229 & n4239 ) ;
  assign n4241 = ( ~n4045 & n4229 ) | ( ~n4045 & n4239 ) | ( n4229 & n4239 ) ;
  assign n4242 = ( n4045 & ~n4240 ) | ( n4045 & n4241 ) | ( ~n4240 & n4241 ) ;
  assign n4243 = n372 & n2982 ;
  assign n4244 = x35 & n4243 ;
  assign n4245 = x72 & n2989 ;
  assign n4246 = x71 & n2986 ;
  assign n4247 = n4245 | n4246 ;
  assign n4248 = x70 & n3159 ;
  assign n4249 = n4247 | n4248 ;
  assign n4250 = ( ~x35 & n4243 ) | ( ~x35 & n4249 ) | ( n4243 & n4249 ) ;
  assign n4251 = x35 & ~n4249 ;
  assign n4252 = ( ~n4244 & n4250 ) | ( ~n4244 & n4251 ) | ( n4250 & n4251 ) ;
  assign n4253 = ( n4047 & ~n4242 ) | ( n4047 & n4252 ) | ( ~n4242 & n4252 ) ;
  assign n4254 = ( n4047 & n4242 ) | ( n4047 & n4252 ) | ( n4242 & n4252 ) ;
  assign n4255 = ( n4242 & n4253 ) | ( n4242 & ~n4254 ) | ( n4253 & ~n4254 ) ;
  assign n4256 = ( n4061 & n4215 ) | ( n4061 & n4255 ) | ( n4215 & n4255 ) ;
  assign n4257 = ( ~n4061 & n4215 ) | ( ~n4061 & n4255 ) | ( n4215 & n4255 ) ;
  assign n4258 = ( n4061 & ~n4256 ) | ( n4061 & n4257 ) | ( ~n4256 & n4257 ) ;
  assign n4259 = ( n4063 & n4205 ) | ( n4063 & n4258 ) | ( n4205 & n4258 ) ;
  assign n4260 = ( ~n4063 & n4205 ) | ( ~n4063 & n4258 ) | ( n4205 & n4258 ) ;
  assign n4261 = ( n4063 & ~n4259 ) | ( n4063 & n4260 ) | ( ~n4259 & n4260 ) ;
  assign n4262 = n990 & n1755 ;
  assign n4263 = x26 & n4262 ;
  assign n4264 = x81 & n1762 ;
  assign n4265 = x80 & n1759 ;
  assign n4266 = n4264 | n4265 ;
  assign n4267 = x79 & n1895 ;
  assign n4268 = n4266 | n4267 ;
  assign n4269 = ( ~x26 & n4262 ) | ( ~x26 & n4268 ) | ( n4262 & n4268 ) ;
  assign n4270 = x26 & ~n4268 ;
  assign n4271 = ( ~n4263 & n4269 ) | ( ~n4263 & n4270 ) | ( n4269 & n4270 ) ;
  assign n4272 = ( n4077 & n4261 ) | ( n4077 & n4271 ) | ( n4261 & n4271 ) ;
  assign n4273 = ( ~n4077 & n4261 ) | ( ~n4077 & n4271 ) | ( n4261 & n4271 ) ;
  assign n4274 = ( n4077 & ~n4272 ) | ( n4077 & n4273 ) | ( ~n4272 & n4273 ) ;
  assign n4275 = n1190 & n1427 ;
  assign n4276 = x23 & n4275 ;
  assign n4277 = x84 & n1434 ;
  assign n4278 = x83 & n1431 ;
  assign n4279 = n4277 | n4278 ;
  assign n4280 = x82 & n1531 ;
  assign n4281 = n4279 | n4280 ;
  assign n4282 = ( ~x23 & n4275 ) | ( ~x23 & n4281 ) | ( n4275 & n4281 ) ;
  assign n4283 = x23 & ~n4281 ;
  assign n4284 = ( ~n4276 & n4282 ) | ( ~n4276 & n4283 ) | ( n4282 & n4283 ) ;
  assign n4285 = ( n4079 & ~n4274 ) | ( n4079 & n4284 ) | ( ~n4274 & n4284 ) ;
  assign n4286 = ( n4079 & n4274 ) | ( n4079 & n4284 ) | ( n4274 & n4284 ) ;
  assign n4287 = ( n4274 & n4285 ) | ( n4274 & ~n4286 ) | ( n4285 & ~n4286 ) ;
  assign n4288 = ( n4093 & n4195 ) | ( n4093 & n4287 ) | ( n4195 & n4287 ) ;
  assign n4289 = ( ~n4093 & n4195 ) | ( ~n4093 & n4287 ) | ( n4195 & n4287 ) ;
  assign n4290 = ( n4093 & ~n4288 ) | ( n4093 & n4289 ) | ( ~n4288 & n4289 ) ;
  assign n4291 = n874 & n1838 ;
  assign n4292 = x17 & n4291 ;
  assign n4293 = x90 & n881 ;
  assign n4294 = x89 & n878 ;
  assign n4295 = n4293 | n4294 ;
  assign n4296 = x88 & n959 ;
  assign n4297 = n4295 | n4296 ;
  assign n4298 = ( ~x17 & n4291 ) | ( ~x17 & n4297 ) | ( n4291 & n4297 ) ;
  assign n4299 = x17 & ~n4297 ;
  assign n4300 = ( ~n4292 & n4298 ) | ( ~n4292 & n4299 ) | ( n4298 & n4299 ) ;
  assign n4301 = ( n4095 & n4290 ) | ( n4095 & n4300 ) | ( n4290 & n4300 ) ;
  assign n4302 = ( ~n4095 & n4290 ) | ( ~n4095 & n4300 ) | ( n4290 & n4300 ) ;
  assign n4303 = ( n4095 & ~n4301 ) | ( n4095 & n4302 ) | ( ~n4301 & n4302 ) ;
  assign n4304 = n649 & n2220 ;
  assign n4305 = x14 & n4304 ;
  assign n4306 = x93 & n656 ;
  assign n4307 = x92 & n653 ;
  assign n4308 = n4306 | n4307 ;
  assign n4309 = x91 & n744 ;
  assign n4310 = n4308 | n4309 ;
  assign n4311 = ( ~x14 & n4304 ) | ( ~x14 & n4310 ) | ( n4304 & n4310 ) ;
  assign n4312 = x14 & ~n4310 ;
  assign n4313 = ( ~n4305 & n4311 ) | ( ~n4305 & n4312 ) | ( n4311 & n4312 ) ;
  assign n4314 = ( n4109 & n4303 ) | ( n4109 & n4313 ) | ( n4303 & n4313 ) ;
  assign n4315 = ( ~n4109 & n4303 ) | ( ~n4109 & n4313 ) | ( n4303 & n4313 ) ;
  assign n4316 = ( n4109 & ~n4314 ) | ( n4109 & n4315 ) | ( ~n4314 & n4315 ) ;
  assign n4317 = ( n4122 & ~n4185 ) | ( n4122 & n4316 ) | ( ~n4185 & n4316 ) ;
  assign n4318 = ( n4122 & n4185 ) | ( n4122 & n4316 ) | ( n4185 & n4316 ) ;
  assign n4319 = ( n4185 & n4317 ) | ( n4185 & ~n4318 ) | ( n4317 & ~n4318 ) ;
  assign n4320 = ( n4124 & n4175 ) | ( n4124 & n4319 ) | ( n4175 & n4319 ) ;
  assign n4321 = ( ~n4124 & n4175 ) | ( ~n4124 & n4319 ) | ( n4175 & n4319 ) ;
  assign n4322 = ( n4124 & ~n4320 ) | ( n4124 & n4321 ) | ( ~n4320 & n4321 ) ;
  assign n4323 = ( n4138 & ~n4165 ) | ( n4138 & n4322 ) | ( ~n4165 & n4322 ) ;
  assign n4324 = ( n4138 & n4165 ) | ( n4138 & n4322 ) | ( n4165 & n4322 ) ;
  assign n4325 = ( n4165 & n4323 ) | ( n4165 & ~n4324 ) | ( n4323 & ~n4324 ) ;
  assign n4326 = ( n4140 & n4155 ) | ( n4140 & n4325 ) | ( n4155 & n4325 ) ;
  assign n4327 = ( ~n4140 & n4155 ) | ( ~n4140 & n4325 ) | ( n4155 & n4325 ) ;
  assign n4328 = ( n4140 & ~n4326 ) | ( n4140 & n4327 ) | ( ~n4326 & n4327 ) ;
  assign n4329 = ( ~x105 & x106 ) | ( ~x105 & n4144 ) | ( x106 & n4144 ) ;
  assign n4330 = ( x105 & x106 ) | ( x105 & n4144 ) | ( x106 & n4144 ) ;
  assign n4331 = ( x105 & n4329 ) | ( x105 & ~n4330 ) | ( n4329 & ~n4330 ) ;
  assign n4332 = x0 & n4331 ;
  assign n4333 = ( x1 & x2 ) | ( x1 & n4332 ) | ( x2 & n4332 ) ;
  assign n4334 = x105 & n172 ;
  assign n4335 = x106 | n4334 ;
  assign n4336 = ( n147 & n4334 ) | ( n147 & n4335 ) | ( n4334 & n4335 ) ;
  assign n4337 = ( ~x104 & n135 ) | ( ~x104 & n174 ) | ( n135 & n174 ) ;
  assign n4338 = n4336 | n4337 ;
  assign n4339 = n4333 | n4338 ;
  assign n4340 = n4333 & n4338 ;
  assign n4341 = n4339 & ~n4340 ;
  assign n4342 = n301 & n3264 ;
  assign n4343 = x8 & n4342 ;
  assign n4344 = x100 & n309 ;
  assign n4345 = x99 & n306 ;
  assign n4346 = n4344 | n4345 ;
  assign n4347 = x98 & n359 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = ( ~x8 & n4342 ) | ( ~x8 & n4348 ) | ( n4342 & n4348 ) ;
  assign n4350 = x8 & ~n4348 ;
  assign n4351 = ( ~n4343 & n4349 ) | ( ~n4343 & n4350 ) | ( n4349 & n4350 ) ;
  assign n4352 = n874 & n1959 ;
  assign n4353 = x17 & n4352 ;
  assign n4354 = x91 & n881 ;
  assign n4355 = x90 & n878 ;
  assign n4356 = n4354 | n4355 ;
  assign n4357 = x89 & n959 ;
  assign n4358 = n4356 | n4357 ;
  assign n4359 = ( ~x17 & n4352 ) | ( ~x17 & n4358 ) | ( n4352 & n4358 ) ;
  assign n4360 = x17 & ~n4358 ;
  assign n4361 = ( ~n4353 & n4359 ) | ( ~n4353 & n4360 ) | ( n4359 & n4360 ) ;
  assign n4362 = n1368 & n1427 ;
  assign n4363 = x23 & n4362 ;
  assign n4364 = x85 & n1434 ;
  assign n4365 = x84 & n1431 ;
  assign n4366 = n4364 | n4365 ;
  assign n4367 = x83 & n1531 ;
  assign n4368 = n4366 | n4367 ;
  assign n4369 = ( ~x23 & n4362 ) | ( ~x23 & n4368 ) | ( n4362 & n4368 ) ;
  assign n4370 = x23 & ~n4368 ;
  assign n4371 = ( ~n4363 & n4369 ) | ( ~n4363 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = n1006 & n1755 ;
  assign n4373 = x26 & n4372 ;
  assign n4374 = x82 & n1762 ;
  assign n4375 = x81 & n1759 ;
  assign n4376 = n4374 | n4375 ;
  assign n4377 = x80 & n1895 ;
  assign n4378 = n4376 | n4377 ;
  assign n4379 = ( ~x26 & n4372 ) | ( ~x26 & n4378 ) | ( n4372 & n4378 ) ;
  assign n4380 = x26 & ~n4378 ;
  assign n4381 = ( ~n4373 & n4379 ) | ( ~n4373 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4382 = n565 & n2545 ;
  assign n4383 = x32 & n4382 ;
  assign n4384 = x76 & n2552 ;
  assign n4385 = x75 & n2549 ;
  assign n4386 = n4384 | n4385 ;
  assign n4387 = x74 & n2696 ;
  assign n4388 = n4386 | n4387 ;
  assign n4389 = ( ~x32 & n4382 ) | ( ~x32 & n4388 ) | ( n4382 & n4388 ) ;
  assign n4390 = x32 & ~n4388 ;
  assign n4391 = ( ~n4383 & n4389 ) | ( ~n4383 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4392 = n4225 | n4226 ;
  assign n4393 = ~x42 & x64 ;
  assign n4394 = ( ~x41 & n4392 ) | ( ~x41 & n4393 ) | ( n4392 & n4393 ) ;
  assign n4395 = n4392 | n4393 ;
  assign n4396 = x41 & x42 ;
  assign n4397 = x41 | x42 ;
  assign n4398 = ~n4396 & n4397 ;
  assign n4399 = x64 & n4398 ;
  assign n4400 = ~x41 & n4399 ;
  assign n4401 = ( ~n4394 & n4395 ) | ( ~n4394 & n4400 ) | ( n4395 & n4400 ) ;
  assign n4402 = x67 & n4027 ;
  assign n4403 = x66 & n4024 ;
  assign n4404 = x65 & n4223 ;
  assign n4405 = n4403 | n4404 ;
  assign n4406 = n4402 | n4405 ;
  assign n4407 = n169 & n4020 ;
  assign n4408 = n4406 | n4407 ;
  assign n4409 = n4401 | n4408 ;
  assign n4410 = n4401 & n4408 ;
  assign n4411 = n4409 & ~n4410 ;
  assign n4412 = n276 & n3492 ;
  assign n4413 = x38 & n4412 ;
  assign n4414 = x70 & n3499 ;
  assign n4415 = x69 & n3496 ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = x68 & n3662 ;
  assign n4418 = n4416 | n4417 ;
  assign n4419 = ( ~x38 & n4412 ) | ( ~x38 & n4418 ) | ( n4412 & n4418 ) ;
  assign n4420 = x38 & ~n4418 ;
  assign n4421 = ( ~n4413 & n4419 ) | ( ~n4413 & n4420 ) | ( n4419 & n4420 ) ;
  assign n4422 = ( n4240 & n4411 ) | ( n4240 & n4421 ) | ( n4411 & n4421 ) ;
  assign n4423 = ( ~n4240 & n4411 ) | ( ~n4240 & n4421 ) | ( n4411 & n4421 ) ;
  assign n4424 = ( n4240 & ~n4422 ) | ( n4240 & n4423 ) | ( ~n4422 & n4423 ) ;
  assign n4425 = n388 & n2982 ;
  assign n4426 = x35 & n4425 ;
  assign n4427 = x73 & n2989 ;
  assign n4428 = x72 & n2986 ;
  assign n4429 = n4427 | n4428 ;
  assign n4430 = x71 & n3159 ;
  assign n4431 = n4429 | n4430 ;
  assign n4432 = ( ~x35 & n4425 ) | ( ~x35 & n4431 ) | ( n4425 & n4431 ) ;
  assign n4433 = x35 & ~n4431 ;
  assign n4434 = ( ~n4426 & n4432 ) | ( ~n4426 & n4433 ) | ( n4432 & n4433 ) ;
  assign n4435 = ( n4254 & ~n4424 ) | ( n4254 & n4434 ) | ( ~n4424 & n4434 ) ;
  assign n4436 = ( n4254 & n4424 ) | ( n4254 & n4434 ) | ( n4424 & n4434 ) ;
  assign n4437 = ( n4424 & n4435 ) | ( n4424 & ~n4436 ) | ( n4435 & ~n4436 ) ;
  assign n4438 = ( n4256 & n4391 ) | ( n4256 & n4437 ) | ( n4391 & n4437 ) ;
  assign n4439 = ( ~n4256 & n4391 ) | ( ~n4256 & n4437 ) | ( n4391 & n4437 ) ;
  assign n4440 = ( n4256 & ~n4438 ) | ( n4256 & n4439 ) | ( ~n4438 & n4439 ) ;
  assign n4441 = n823 & n2137 ;
  assign n4442 = x29 & n4441 ;
  assign n4443 = x79 & n2144 ;
  assign n4444 = x78 & n2141 ;
  assign n4445 = n4443 | n4444 ;
  assign n4446 = x77 & n2267 ;
  assign n4447 = n4445 | n4446 ;
  assign n4448 = ( ~x29 & n4441 ) | ( ~x29 & n4447 ) | ( n4441 & n4447 ) ;
  assign n4449 = x29 & ~n4447 ;
  assign n4450 = ( ~n4442 & n4448 ) | ( ~n4442 & n4449 ) | ( n4448 & n4449 ) ;
  assign n4451 = ( n4259 & ~n4440 ) | ( n4259 & n4450 ) | ( ~n4440 & n4450 ) ;
  assign n4452 = ( n4259 & n4440 ) | ( n4259 & n4450 ) | ( n4440 & n4450 ) ;
  assign n4453 = ( n4440 & n4451 ) | ( n4440 & ~n4452 ) | ( n4451 & ~n4452 ) ;
  assign n4454 = ( n4272 & n4381 ) | ( n4272 & n4453 ) | ( n4381 & n4453 ) ;
  assign n4455 = ( ~n4272 & n4381 ) | ( ~n4272 & n4453 ) | ( n4381 & n4453 ) ;
  assign n4456 = ( n4272 & ~n4454 ) | ( n4272 & n4455 ) | ( ~n4454 & n4455 ) ;
  assign n4457 = ( n4286 & n4371 ) | ( n4286 & n4456 ) | ( n4371 & n4456 ) ;
  assign n4458 = ( ~n4286 & n4371 ) | ( ~n4286 & n4456 ) | ( n4371 & n4456 ) ;
  assign n4459 = ( n4286 & ~n4457 ) | ( n4286 & n4458 ) | ( ~n4457 & n4458 ) ;
  assign n4460 = n1146 & n1602 ;
  assign n4461 = x20 & n4460 ;
  assign n4462 = x88 & n1153 ;
  assign n4463 = x87 & n1150 ;
  assign n4464 = n4462 | n4463 ;
  assign n4465 = x86 & n1217 ;
  assign n4466 = n4464 | n4465 ;
  assign n4467 = ( ~x20 & n4460 ) | ( ~x20 & n4466 ) | ( n4460 & n4466 ) ;
  assign n4468 = x20 & ~n4466 ;
  assign n4469 = ( ~n4461 & n4467 ) | ( ~n4461 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4470 = ( n4288 & ~n4459 ) | ( n4288 & n4469 ) | ( ~n4459 & n4469 ) ;
  assign n4471 = ( n4288 & n4459 ) | ( n4288 & n4469 ) | ( n4459 & n4469 ) ;
  assign n4472 = ( n4459 & n4470 ) | ( n4459 & ~n4471 ) | ( n4470 & ~n4471 ) ;
  assign n4473 = ( n4301 & n4361 ) | ( n4301 & n4472 ) | ( n4361 & n4472 ) ;
  assign n4474 = ( ~n4301 & n4361 ) | ( ~n4301 & n4472 ) | ( n4361 & n4472 ) ;
  assign n4475 = ( n4301 & ~n4473 ) | ( n4301 & n4474 ) | ( ~n4473 & n4474 ) ;
  assign n4476 = n649 & n2476 ;
  assign n4477 = x14 & n4476 ;
  assign n4478 = x94 & n656 ;
  assign n4479 = x93 & n653 ;
  assign n4480 = n4478 | n4479 ;
  assign n4481 = x92 & n744 ;
  assign n4482 = n4480 | n4481 ;
  assign n4483 = ( ~x14 & n4476 ) | ( ~x14 & n4482 ) | ( n4476 & n4482 ) ;
  assign n4484 = x14 & ~n4482 ;
  assign n4485 = ( ~n4477 & n4483 ) | ( ~n4477 & n4484 ) | ( n4483 & n4484 ) ;
  assign n4486 = ( n4314 & ~n4475 ) | ( n4314 & n4485 ) | ( ~n4475 & n4485 ) ;
  assign n4487 = ( n4314 & n4475 ) | ( n4314 & n4485 ) | ( n4475 & n4485 ) ;
  assign n4488 = ( n4475 & n4486 ) | ( n4475 & ~n4487 ) | ( n4486 & ~n4487 ) ;
  assign n4489 = n449 & n2788 ;
  assign n4490 = x11 & n4489 ;
  assign n4491 = x97 & n456 ;
  assign n4492 = x96 & n453 ;
  assign n4493 = n4491 | n4492 ;
  assign n4494 = x95 & n536 ;
  assign n4495 = n4493 | n4494 ;
  assign n4496 = ( ~x11 & n4489 ) | ( ~x11 & n4495 ) | ( n4489 & n4495 ) ;
  assign n4497 = x11 & ~n4495 ;
  assign n4498 = ( ~n4490 & n4496 ) | ( ~n4490 & n4497 ) | ( n4496 & n4497 ) ;
  assign n4499 = ( n4318 & ~n4488 ) | ( n4318 & n4498 ) | ( ~n4488 & n4498 ) ;
  assign n4500 = ( n4318 & n4488 ) | ( n4318 & n4498 ) | ( n4488 & n4498 ) ;
  assign n4501 = ( n4488 & n4499 ) | ( n4488 & ~n4500 ) | ( n4499 & ~n4500 ) ;
  assign n4502 = ( n4320 & n4351 ) | ( n4320 & n4501 ) | ( n4351 & n4501 ) ;
  assign n4503 = ( ~n4320 & n4351 ) | ( ~n4320 & n4501 ) | ( n4351 & n4501 ) ;
  assign n4504 = ( n4320 & ~n4502 ) | ( n4320 & n4503 ) | ( ~n4502 & n4503 ) ;
  assign n4505 = n206 & n3941 ;
  assign n4506 = x5 & n4505 ;
  assign n4507 = x103 & n205 ;
  assign n4508 = x102 & n201 ;
  assign n4509 = n4507 | n4508 ;
  assign n4510 = x101 & n221 ;
  assign n4511 = n4509 | n4510 ;
  assign n4512 = ( ~x5 & n4505 ) | ( ~x5 & n4511 ) | ( n4505 & n4511 ) ;
  assign n4513 = x5 & ~n4511 ;
  assign n4514 = ( ~n4506 & n4512 ) | ( ~n4506 & n4513 ) | ( n4512 & n4513 ) ;
  assign n4515 = ( n4324 & ~n4504 ) | ( n4324 & n4514 ) | ( ~n4504 & n4514 ) ;
  assign n4516 = ( n4324 & n4504 ) | ( n4324 & n4514 ) | ( n4504 & n4514 ) ;
  assign n4517 = ( n4504 & n4515 ) | ( n4504 & ~n4516 ) | ( n4515 & ~n4516 ) ;
  assign n4518 = ( n4326 & n4341 ) | ( n4326 & n4517 ) | ( n4341 & n4517 ) ;
  assign n4519 = ( ~n4326 & n4341 ) | ( ~n4326 & n4517 ) | ( n4341 & n4517 ) ;
  assign n4520 = ( n4326 & ~n4518 ) | ( n4326 & n4519 ) | ( ~n4518 & n4519 ) ;
  assign n4521 = ( ~x106 & x107 ) | ( ~x106 & n4330 ) | ( x107 & n4330 ) ;
  assign n4522 = ( x106 & x107 ) | ( x106 & n4330 ) | ( x107 & n4330 ) ;
  assign n4523 = ( x106 & n4521 ) | ( x106 & ~n4522 ) | ( n4521 & ~n4522 ) ;
  assign n4524 = x0 & n4523 ;
  assign n4525 = ( x1 & x2 ) | ( x1 & n4524 ) | ( x2 & n4524 ) ;
  assign n4526 = x106 & n172 ;
  assign n4527 = ( ~x105 & n135 ) | ( ~x105 & n174 ) | ( n135 & n174 ) ;
  assign n4528 = n4526 | n4527 ;
  assign n4529 = x107 & n147 ;
  assign n4530 = n4528 | n4529 ;
  assign n4531 = n4525 | n4530 ;
  assign n4532 = n4525 & n4530 ;
  assign n4533 = n4531 & ~n4532 ;
  assign n4534 = n206 & n3957 ;
  assign n4535 = x5 & n4534 ;
  assign n4536 = x104 & n205 ;
  assign n4537 = x103 & n201 ;
  assign n4538 = n4536 | n4537 ;
  assign n4539 = x102 & n221 ;
  assign n4540 = n4538 | n4539 ;
  assign n4541 = ( ~x5 & n4534 ) | ( ~x5 & n4540 ) | ( n4534 & n4540 ) ;
  assign n4542 = x5 & ~n4540 ;
  assign n4543 = ( ~n4535 & n4541 ) | ( ~n4535 & n4542 ) | ( n4541 & n4542 ) ;
  assign n4544 = n301 & n3591 ;
  assign n4545 = x8 & n4544 ;
  assign n4546 = x101 & n309 ;
  assign n4547 = x100 & n306 ;
  assign n4548 = n4546 | n4547 ;
  assign n4549 = x99 & n359 ;
  assign n4550 = n4548 | n4549 ;
  assign n4551 = ( ~x8 & n4544 ) | ( ~x8 & n4550 ) | ( n4544 & n4550 ) ;
  assign n4552 = x8 & ~n4550 ;
  assign n4553 = ( ~n4545 & n4551 ) | ( ~n4545 & n4552 ) | ( n4551 & n4552 ) ;
  assign n4554 = n649 & n2492 ;
  assign n4555 = x14 & n4554 ;
  assign n4556 = x95 & n656 ;
  assign n4557 = x94 & n653 ;
  assign n4558 = n4556 | n4557 ;
  assign n4559 = x93 & n744 ;
  assign n4560 = n4558 | n4559 ;
  assign n4561 = ( ~x14 & n4554 ) | ( ~x14 & n4560 ) | ( n4554 & n4560 ) ;
  assign n4562 = x14 & ~n4560 ;
  assign n4563 = ( ~n4555 & n4561 ) | ( ~n4555 & n4562 ) | ( n4561 & n4562 ) ;
  assign n4564 = n1146 & n1822 ;
  assign n4565 = x20 & n4564 ;
  assign n4566 = x89 & n1153 ;
  assign n4567 = x88 & n1150 ;
  assign n4568 = n4566 | n4567 ;
  assign n4569 = x87 & n1217 ;
  assign n4570 = n4568 | n4569 ;
  assign n4571 = ( ~x20 & n4564 ) | ( ~x20 & n4570 ) | ( n4564 & n4570 ) ;
  assign n4572 = x20 & ~n4570 ;
  assign n4573 = ( ~n4565 & n4571 ) | ( ~n4565 & n4572 ) | ( n4571 & n4572 ) ;
  assign n4574 = n1093 & n1755 ;
  assign n4575 = x26 & n4574 ;
  assign n4576 = x83 & n1762 ;
  assign n4577 = x82 & n1759 ;
  assign n4578 = n4576 | n4577 ;
  assign n4579 = x81 & n1895 ;
  assign n4580 = n4578 | n4579 ;
  assign n4581 = ( ~x26 & n4574 ) | ( ~x26 & n4580 ) | ( n4574 & n4580 ) ;
  assign n4582 = x26 & ~n4580 ;
  assign n4583 = ( ~n4575 & n4581 ) | ( ~n4575 & n4582 ) | ( n4581 & n4582 ) ;
  assign n4584 = n626 & n2545 ;
  assign n4585 = x32 & n4584 ;
  assign n4586 = x77 & n2552 ;
  assign n4587 = x76 & n2549 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = x75 & n2696 ;
  assign n4590 = n4588 | n4589 ;
  assign n4591 = ( ~x32 & n4584 ) | ( ~x32 & n4590 ) | ( n4584 & n4590 ) ;
  assign n4592 = x32 & ~n4590 ;
  assign n4593 = ( ~n4585 & n4591 ) | ( ~n4585 & n4592 ) | ( n4591 & n4592 ) ;
  assign n4594 = n322 & n3492 ;
  assign n4595 = x38 & n4594 ;
  assign n4596 = x71 & n3499 ;
  assign n4597 = x70 & n3496 ;
  assign n4598 = n4596 | n4597 ;
  assign n4599 = x69 & n3662 ;
  assign n4600 = n4598 | n4599 ;
  assign n4601 = ( ~x38 & n4594 ) | ( ~x38 & n4600 ) | ( n4594 & n4600 ) ;
  assign n4602 = x38 & ~n4600 ;
  assign n4603 = ( ~n4595 & n4601 ) | ( ~n4595 & n4602 ) | ( n4601 & n4602 ) ;
  assign n4604 = x68 & n4027 ;
  assign n4605 = x41 & n4604 ;
  assign n4606 = x67 & n4024 ;
  assign n4607 = x66 & n4223 ;
  assign n4608 = n4606 | n4607 ;
  assign n4609 = n193 & n4020 ;
  assign n4610 = n4608 | n4609 ;
  assign n4611 = ( ~x41 & n4604 ) | ( ~x41 & n4610 ) | ( n4604 & n4610 ) ;
  assign n4612 = x41 & ~n4610 ;
  assign n4613 = ( ~n4605 & n4611 ) | ( ~n4605 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4614 = n4400 & n4408 ;
  assign n4615 = x41 & n4393 ;
  assign n4616 = ( x41 & ~n4392 ) | ( x41 & n4615 ) | ( ~n4392 & n4615 ) ;
  assign n4617 = n4408 & ~n4614 ;
  assign n4618 = ( n4614 & n4616 ) | ( n4614 & ~n4617 ) | ( n4616 & ~n4617 ) ;
  assign n4619 = ~x41 & x43 ;
  assign n4620 = x42 & x43 ;
  assign n4621 = ( n4396 & n4619 ) | ( n4396 & ~n4620 ) | ( n4619 & ~n4620 ) ;
  assign n4622 = x43 & x44 ;
  assign n4623 = x43 | x44 ;
  assign n4624 = ~n4622 & n4623 ;
  assign n4625 = n4398 & n4624 ;
  assign n4626 = x65 & ~n4621 ;
  assign n4627 = ( n4621 & n4625 ) | ( n4621 & ~n4626 ) | ( n4625 & ~n4626 ) ;
  assign n4628 = x64 & n4627 ;
  assign n4629 = ( x65 & n138 ) | ( x65 & ~n4624 ) | ( n138 & ~n4624 ) ;
  assign n4630 = n4398 & n4629 ;
  assign n4631 = n4628 | n4630 ;
  assign n4632 = x44 | n4631 ;
  assign n4633 = ~n4399 & n4631 ;
  assign n4634 = ( x44 & ~n4399 ) | ( x44 & n4631 ) | ( ~n4399 & n4631 ) ;
  assign n4635 = ( n4632 & n4633 ) | ( n4632 & ~n4634 ) | ( n4633 & ~n4634 ) ;
  assign n4636 = ( ~n4613 & n4618 ) | ( ~n4613 & n4635 ) | ( n4618 & n4635 ) ;
  assign n4637 = ( n4613 & n4618 ) | ( n4613 & n4635 ) | ( n4618 & n4635 ) ;
  assign n4638 = ( n4613 & n4636 ) | ( n4613 & ~n4637 ) | ( n4636 & ~n4637 ) ;
  assign n4639 = ( n4422 & n4603 ) | ( n4422 & n4638 ) | ( n4603 & n4638 ) ;
  assign n4640 = ( ~n4422 & n4603 ) | ( ~n4422 & n4638 ) | ( n4603 & n4638 ) ;
  assign n4641 = ( n4422 & ~n4639 ) | ( n4422 & n4640 ) | ( ~n4639 & n4640 ) ;
  assign n4642 = n436 & n2982 ;
  assign n4643 = x35 & n4642 ;
  assign n4644 = x74 & n2989 ;
  assign n4645 = x73 & n2986 ;
  assign n4646 = n4644 | n4645 ;
  assign n4647 = x72 & n3159 ;
  assign n4648 = n4646 | n4647 ;
  assign n4649 = ( ~x35 & n4642 ) | ( ~x35 & n4648 ) | ( n4642 & n4648 ) ;
  assign n4650 = x35 & ~n4648 ;
  assign n4651 = ( ~n4643 & n4649 ) | ( ~n4643 & n4650 ) | ( n4649 & n4650 ) ;
  assign n4652 = ( n4436 & ~n4641 ) | ( n4436 & n4651 ) | ( ~n4641 & n4651 ) ;
  assign n4653 = ( n4436 & n4641 ) | ( n4436 & n4651 ) | ( n4641 & n4651 ) ;
  assign n4654 = ( n4641 & n4652 ) | ( n4641 & ~n4653 ) | ( n4652 & ~n4653 ) ;
  assign n4655 = ( n4438 & n4593 ) | ( n4438 & n4654 ) | ( n4593 & n4654 ) ;
  assign n4656 = ( ~n4438 & n4593 ) | ( ~n4438 & n4654 ) | ( n4593 & n4654 ) ;
  assign n4657 = ( n4438 & ~n4655 ) | ( n4438 & n4656 ) | ( ~n4655 & n4656 ) ;
  assign n4658 = n840 & n2137 ;
  assign n4659 = x29 & n4658 ;
  assign n4660 = x80 & n2144 ;
  assign n4661 = x79 & n2141 ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = x78 & n2267 ;
  assign n4664 = n4662 | n4663 ;
  assign n4665 = ( ~x29 & n4658 ) | ( ~x29 & n4664 ) | ( n4658 & n4664 ) ;
  assign n4666 = x29 & ~n4664 ;
  assign n4667 = ( ~n4659 & n4665 ) | ( ~n4659 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4668 = ( n4452 & ~n4657 ) | ( n4452 & n4667 ) | ( ~n4657 & n4667 ) ;
  assign n4669 = ( n4452 & n4657 ) | ( n4452 & n4667 ) | ( n4657 & n4667 ) ;
  assign n4670 = ( n4657 & n4668 ) | ( n4657 & ~n4669 ) | ( n4668 & ~n4669 ) ;
  assign n4671 = ( n4454 & n4583 ) | ( n4454 & n4670 ) | ( n4583 & n4670 ) ;
  assign n4672 = ( ~n4454 & n4583 ) | ( ~n4454 & n4670 ) | ( n4583 & n4670 ) ;
  assign n4673 = ( n4454 & ~n4671 ) | ( n4454 & n4672 ) | ( ~n4671 & n4672 ) ;
  assign n4674 = n1384 & n1427 ;
  assign n4675 = x23 & n4674 ;
  assign n4676 = x86 & n1434 ;
  assign n4677 = x85 & n1431 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = x84 & n1531 ;
  assign n4680 = n4678 | n4679 ;
  assign n4681 = ( ~x23 & n4674 ) | ( ~x23 & n4680 ) | ( n4674 & n4680 ) ;
  assign n4682 = x23 & ~n4680 ;
  assign n4683 = ( ~n4675 & n4681 ) | ( ~n4675 & n4682 ) | ( n4681 & n4682 ) ;
  assign n4684 = ( n4457 & ~n4673 ) | ( n4457 & n4683 ) | ( ~n4673 & n4683 ) ;
  assign n4685 = ( n4457 & n4673 ) | ( n4457 & n4683 ) | ( n4673 & n4683 ) ;
  assign n4686 = ( n4673 & n4684 ) | ( n4673 & ~n4685 ) | ( n4684 & ~n4685 ) ;
  assign n4687 = ( n4471 & n4573 ) | ( n4471 & n4686 ) | ( n4573 & n4686 ) ;
  assign n4688 = ( ~n4471 & n4573 ) | ( ~n4471 & n4686 ) | ( n4573 & n4686 ) ;
  assign n4689 = ( n4471 & ~n4687 ) | ( n4471 & n4688 ) | ( ~n4687 & n4688 ) ;
  assign n4690 = n874 & n2083 ;
  assign n4691 = x17 & n4690 ;
  assign n4692 = x92 & n881 ;
  assign n4693 = x91 & n878 ;
  assign n4694 = n4692 | n4693 ;
  assign n4695 = x90 & n959 ;
  assign n4696 = n4694 | n4695 ;
  assign n4697 = ( ~x17 & n4690 ) | ( ~x17 & n4696 ) | ( n4690 & n4696 ) ;
  assign n4698 = x17 & ~n4696 ;
  assign n4699 = ( ~n4691 & n4697 ) | ( ~n4691 & n4698 ) | ( n4697 & n4698 ) ;
  assign n4700 = ( n4473 & ~n4689 ) | ( n4473 & n4699 ) | ( ~n4689 & n4699 ) ;
  assign n4701 = ( n4473 & n4689 ) | ( n4473 & n4699 ) | ( n4689 & n4699 ) ;
  assign n4702 = ( n4689 & n4700 ) | ( n4689 & ~n4701 ) | ( n4700 & ~n4701 ) ;
  assign n4703 = ( n4487 & n4563 ) | ( n4487 & n4702 ) | ( n4563 & n4702 ) ;
  assign n4704 = ( ~n4487 & n4563 ) | ( ~n4487 & n4702 ) | ( n4563 & n4702 ) ;
  assign n4705 = ( n4487 & ~n4703 ) | ( n4487 & n4704 ) | ( ~n4703 & n4704 ) ;
  assign n4706 = n449 & n2939 ;
  assign n4707 = x11 & n4706 ;
  assign n4708 = x98 & n456 ;
  assign n4709 = x97 & n453 ;
  assign n4710 = n4708 | n4709 ;
  assign n4711 = x96 & n536 ;
  assign n4712 = n4710 | n4711 ;
  assign n4713 = ( ~x11 & n4706 ) | ( ~x11 & n4712 ) | ( n4706 & n4712 ) ;
  assign n4714 = x11 & ~n4712 ;
  assign n4715 = ( ~n4707 & n4713 ) | ( ~n4707 & n4714 ) | ( n4713 & n4714 ) ;
  assign n4716 = ( n4500 & ~n4705 ) | ( n4500 & n4715 ) | ( ~n4705 & n4715 ) ;
  assign n4717 = ( n4500 & n4705 ) | ( n4500 & n4715 ) | ( n4705 & n4715 ) ;
  assign n4718 = ( n4705 & n4716 ) | ( n4705 & ~n4717 ) | ( n4716 & ~n4717 ) ;
  assign n4719 = ( n4502 & n4553 ) | ( n4502 & n4718 ) | ( n4553 & n4718 ) ;
  assign n4720 = ( ~n4502 & n4553 ) | ( ~n4502 & n4718 ) | ( n4553 & n4718 ) ;
  assign n4721 = ( n4502 & ~n4719 ) | ( n4502 & n4720 ) | ( ~n4719 & n4720 ) ;
  assign n4722 = ( n4516 & ~n4543 ) | ( n4516 & n4721 ) | ( ~n4543 & n4721 ) ;
  assign n4723 = ( n4516 & n4543 ) | ( n4516 & n4721 ) | ( n4543 & n4721 ) ;
  assign n4724 = ( n4543 & n4722 ) | ( n4543 & ~n4723 ) | ( n4722 & ~n4723 ) ;
  assign n4725 = ( n4518 & n4533 ) | ( n4518 & n4724 ) | ( n4533 & n4724 ) ;
  assign n4726 = ( ~n4518 & n4533 ) | ( ~n4518 & n4724 ) | ( n4533 & n4724 ) ;
  assign n4727 = ( n4518 & ~n4725 ) | ( n4518 & n4726 ) | ( ~n4725 & n4726 ) ;
  assign n4728 = n206 & n4145 ;
  assign n4729 = x5 & n4728 ;
  assign n4730 = x105 & n205 ;
  assign n4731 = x104 & n201 ;
  assign n4732 = n4730 | n4731 ;
  assign n4733 = x103 & n221 ;
  assign n4734 = n4732 | n4733 ;
  assign n4735 = ( ~x5 & n4728 ) | ( ~x5 & n4734 ) | ( n4728 & n4734 ) ;
  assign n4736 = x5 & ~n4734 ;
  assign n4737 = ( ~n4729 & n4735 ) | ( ~n4729 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4738 = n301 & n3764 ;
  assign n4739 = x8 & n4738 ;
  assign n4740 = x102 & n309 ;
  assign n4741 = x101 & n306 ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = x100 & n359 ;
  assign n4744 = n4742 | n4743 ;
  assign n4745 = ( ~x8 & n4738 ) | ( ~x8 & n4744 ) | ( n4738 & n4744 ) ;
  assign n4746 = x8 & ~n4744 ;
  assign n4747 = ( ~n4739 & n4745 ) | ( ~n4739 & n4746 ) | ( n4745 & n4746 ) ;
  assign n4748 = n874 & n2220 ;
  assign n4749 = x17 & n4748 ;
  assign n4750 = x93 & n881 ;
  assign n4751 = x92 & n878 ;
  assign n4752 = n4750 | n4751 ;
  assign n4753 = x91 & n959 ;
  assign n4754 = n4752 | n4753 ;
  assign n4755 = ( ~x17 & n4748 ) | ( ~x17 & n4754 ) | ( n4748 & n4754 ) ;
  assign n4756 = x17 & ~n4754 ;
  assign n4757 = ( ~n4749 & n4755 ) | ( ~n4749 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = n1427 & n1494 ;
  assign n4759 = x23 & n4758 ;
  assign n4760 = x87 & n1434 ;
  assign n4761 = x86 & n1431 ;
  assign n4762 = n4760 | n4761 ;
  assign n4763 = x85 & n1531 ;
  assign n4764 = n4762 | n4763 ;
  assign n4765 = ( ~x23 & n4758 ) | ( ~x23 & n4764 ) | ( n4758 & n4764 ) ;
  assign n4766 = x23 & ~n4764 ;
  assign n4767 = ( ~n4759 & n4765 ) | ( ~n4759 & n4766 ) | ( n4765 & n4766 ) ;
  assign n4768 = n990 & n2137 ;
  assign n4769 = x29 & n4768 ;
  assign n4770 = x81 & n2144 ;
  assign n4771 = x80 & n2141 ;
  assign n4772 = n4770 | n4771 ;
  assign n4773 = x79 & n2267 ;
  assign n4774 = n4772 | n4773 ;
  assign n4775 = ( ~x29 & n4768 ) | ( ~x29 & n4774 ) | ( n4768 & n4774 ) ;
  assign n4776 = x29 & ~n4774 ;
  assign n4777 = ( ~n4769 & n4775 ) | ( ~n4769 & n4776 ) | ( n4775 & n4776 ) ;
  assign n4778 = n508 & n2982 ;
  assign n4779 = x35 & n4778 ;
  assign n4780 = x75 & n2989 ;
  assign n4781 = x74 & n2986 ;
  assign n4782 = n4780 | n4781 ;
  assign n4783 = x73 & n3159 ;
  assign n4784 = n4782 | n4783 ;
  assign n4785 = ( ~x35 & n4778 ) | ( ~x35 & n4784 ) | ( n4778 & n4784 ) ;
  assign n4786 = x35 & ~n4784 ;
  assign n4787 = ( ~n4779 & n4785 ) | ( ~n4779 & n4786 ) | ( n4785 & n4786 ) ;
  assign n4788 = x65 & n4621 ;
  assign n4789 = n226 & n4625 ;
  assign n4790 = n4788 | n4789 ;
  assign n4791 = ( n4398 & n4622 ) | ( n4398 & ~n4623 ) | ( n4622 & ~n4623 ) ;
  assign n4792 = x66 & n4791 ;
  assign n4793 = n4790 | n4792 ;
  assign n4794 = ~n4398 & n4624 ;
  assign n4795 = ~n4621 & n4794 ;
  assign n4796 = x64 & n4795 ;
  assign n4797 = n4793 | n4796 ;
  assign n4798 = x44 & n4399 ;
  assign n4799 = ( x44 & n4631 ) | ( x44 & n4798 ) | ( n4631 & n4798 ) ;
  assign n4800 = ~n4797 & n4799 ;
  assign n4801 = n4797 & ~n4799 ;
  assign n4802 = n4800 | n4801 ;
  assign n4803 = n240 & n4020 ;
  assign n4804 = x41 & n4803 ;
  assign n4805 = x69 & n4027 ;
  assign n4806 = x68 & n4024 ;
  assign n4807 = n4805 | n4806 ;
  assign n4808 = x67 & n4223 ;
  assign n4809 = n4807 | n4808 ;
  assign n4810 = ( ~x41 & n4803 ) | ( ~x41 & n4809 ) | ( n4803 & n4809 ) ;
  assign n4811 = x41 & ~n4809 ;
  assign n4812 = ( ~n4804 & n4810 ) | ( ~n4804 & n4811 ) | ( n4810 & n4811 ) ;
  assign n4813 = ( n4637 & n4802 ) | ( n4637 & n4812 ) | ( n4802 & n4812 ) ;
  assign n4814 = ( ~n4637 & n4802 ) | ( ~n4637 & n4812 ) | ( n4802 & n4812 ) ;
  assign n4815 = ( n4637 & ~n4813 ) | ( n4637 & n4814 ) | ( ~n4813 & n4814 ) ;
  assign n4816 = n372 & n3492 ;
  assign n4817 = x38 & n4816 ;
  assign n4818 = x72 & n3499 ;
  assign n4819 = x71 & n3496 ;
  assign n4820 = n4818 | n4819 ;
  assign n4821 = x70 & n3662 ;
  assign n4822 = n4820 | n4821 ;
  assign n4823 = ( ~x38 & n4816 ) | ( ~x38 & n4822 ) | ( n4816 & n4822 ) ;
  assign n4824 = x38 & ~n4822 ;
  assign n4825 = ( ~n4817 & n4823 ) | ( ~n4817 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4826 = ( n4639 & ~n4815 ) | ( n4639 & n4825 ) | ( ~n4815 & n4825 ) ;
  assign n4827 = ( n4639 & n4815 ) | ( n4639 & n4825 ) | ( n4815 & n4825 ) ;
  assign n4828 = ( n4815 & n4826 ) | ( n4815 & ~n4827 ) | ( n4826 & ~n4827 ) ;
  assign n4829 = ( n4653 & n4787 ) | ( n4653 & n4828 ) | ( n4787 & n4828 ) ;
  assign n4830 = ( ~n4653 & n4787 ) | ( ~n4653 & n4828 ) | ( n4787 & n4828 ) ;
  assign n4831 = ( n4653 & ~n4829 ) | ( n4653 & n4830 ) | ( ~n4829 & n4830 ) ;
  assign n4832 = n697 & n2545 ;
  assign n4833 = x32 & n4832 ;
  assign n4834 = x78 & n2552 ;
  assign n4835 = x77 & n2549 ;
  assign n4836 = n4834 | n4835 ;
  assign n4837 = x76 & n2696 ;
  assign n4838 = n4836 | n4837 ;
  assign n4839 = ( ~x32 & n4832 ) | ( ~x32 & n4838 ) | ( n4832 & n4838 ) ;
  assign n4840 = x32 & ~n4838 ;
  assign n4841 = ( ~n4833 & n4839 ) | ( ~n4833 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4842 = ( n4655 & ~n4831 ) | ( n4655 & n4841 ) | ( ~n4831 & n4841 ) ;
  assign n4843 = ( n4655 & n4831 ) | ( n4655 & n4841 ) | ( n4831 & n4841 ) ;
  assign n4844 = ( n4831 & n4842 ) | ( n4831 & ~n4843 ) | ( n4842 & ~n4843 ) ;
  assign n4845 = ( n4669 & n4777 ) | ( n4669 & n4844 ) | ( n4777 & n4844 ) ;
  assign n4846 = ( ~n4669 & n4777 ) | ( ~n4669 & n4844 ) | ( n4777 & n4844 ) ;
  assign n4847 = ( n4669 & ~n4845 ) | ( n4669 & n4846 ) | ( ~n4845 & n4846 ) ;
  assign n4848 = n1190 & n1755 ;
  assign n4849 = x26 & n4848 ;
  assign n4850 = x84 & n1762 ;
  assign n4851 = x83 & n1759 ;
  assign n4852 = n4850 | n4851 ;
  assign n4853 = x82 & n1895 ;
  assign n4854 = n4852 | n4853 ;
  assign n4855 = ( ~x26 & n4848 ) | ( ~x26 & n4854 ) | ( n4848 & n4854 ) ;
  assign n4856 = x26 & ~n4854 ;
  assign n4857 = ( ~n4849 & n4855 ) | ( ~n4849 & n4856 ) | ( n4855 & n4856 ) ;
  assign n4858 = ( n4671 & ~n4847 ) | ( n4671 & n4857 ) | ( ~n4847 & n4857 ) ;
  assign n4859 = ( n4671 & n4847 ) | ( n4671 & n4857 ) | ( n4847 & n4857 ) ;
  assign n4860 = ( n4847 & n4858 ) | ( n4847 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  assign n4861 = ( n4685 & n4767 ) | ( n4685 & n4860 ) | ( n4767 & n4860 ) ;
  assign n4862 = ( ~n4685 & n4767 ) | ( ~n4685 & n4860 ) | ( n4767 & n4860 ) ;
  assign n4863 = ( n4685 & ~n4861 ) | ( n4685 & n4862 ) | ( ~n4861 & n4862 ) ;
  assign n4864 = n1146 & n1838 ;
  assign n4865 = x20 & n4864 ;
  assign n4866 = x90 & n1153 ;
  assign n4867 = x89 & n1150 ;
  assign n4868 = n4866 | n4867 ;
  assign n4869 = x88 & n1217 ;
  assign n4870 = n4868 | n4869 ;
  assign n4871 = ( ~x20 & n4864 ) | ( ~x20 & n4870 ) | ( n4864 & n4870 ) ;
  assign n4872 = x20 & ~n4870 ;
  assign n4873 = ( ~n4865 & n4871 ) | ( ~n4865 & n4872 ) | ( n4871 & n4872 ) ;
  assign n4874 = ( n4687 & ~n4863 ) | ( n4687 & n4873 ) | ( ~n4863 & n4873 ) ;
  assign n4875 = ( n4687 & n4863 ) | ( n4687 & n4873 ) | ( n4863 & n4873 ) ;
  assign n4876 = ( n4863 & n4874 ) | ( n4863 & ~n4875 ) | ( n4874 & ~n4875 ) ;
  assign n4877 = ( n4701 & n4757 ) | ( n4701 & n4876 ) | ( n4757 & n4876 ) ;
  assign n4878 = ( ~n4701 & n4757 ) | ( ~n4701 & n4876 ) | ( n4757 & n4876 ) ;
  assign n4879 = ( n4701 & ~n4877 ) | ( n4701 & n4878 ) | ( ~n4877 & n4878 ) ;
  assign n4880 = n649 & n2772 ;
  assign n4881 = x14 & n4880 ;
  assign n4882 = x96 & n656 ;
  assign n4883 = x95 & n653 ;
  assign n4884 = n4882 | n4883 ;
  assign n4885 = x94 & n744 ;
  assign n4886 = n4884 | n4885 ;
  assign n4887 = ( ~x14 & n4880 ) | ( ~x14 & n4886 ) | ( n4880 & n4886 ) ;
  assign n4888 = x14 & ~n4886 ;
  assign n4889 = ( ~n4881 & n4887 ) | ( ~n4881 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4890 = ( n4703 & ~n4879 ) | ( n4703 & n4889 ) | ( ~n4879 & n4889 ) ;
  assign n4891 = ( n4703 & n4879 ) | ( n4703 & n4889 ) | ( n4879 & n4889 ) ;
  assign n4892 = ( n4879 & n4890 ) | ( n4879 & ~n4891 ) | ( n4890 & ~n4891 ) ;
  assign n4893 = n449 & n3248 ;
  assign n4894 = x11 & n4893 ;
  assign n4895 = x99 & n456 ;
  assign n4896 = x98 & n453 ;
  assign n4897 = n4895 | n4896 ;
  assign n4898 = x97 & n536 ;
  assign n4899 = n4897 | n4898 ;
  assign n4900 = ( ~x11 & n4893 ) | ( ~x11 & n4899 ) | ( n4893 & n4899 ) ;
  assign n4901 = x11 & ~n4899 ;
  assign n4902 = ( ~n4894 & n4900 ) | ( ~n4894 & n4901 ) | ( n4900 & n4901 ) ;
  assign n4903 = ( n4717 & ~n4892 ) | ( n4717 & n4902 ) | ( ~n4892 & n4902 ) ;
  assign n4904 = ( n4717 & n4892 ) | ( n4717 & n4902 ) | ( n4892 & n4902 ) ;
  assign n4905 = ( n4892 & n4903 ) | ( n4892 & ~n4904 ) | ( n4903 & ~n4904 ) ;
  assign n4906 = ( n4719 & n4747 ) | ( n4719 & n4905 ) | ( n4747 & n4905 ) ;
  assign n4907 = ( ~n4719 & n4747 ) | ( ~n4719 & n4905 ) | ( n4747 & n4905 ) ;
  assign n4908 = ( n4719 & ~n4906 ) | ( n4719 & n4907 ) | ( ~n4906 & n4907 ) ;
  assign n4909 = ( n4723 & n4737 ) | ( n4723 & n4908 ) | ( n4737 & n4908 ) ;
  assign n4910 = ( ~n4723 & n4737 ) | ( ~n4723 & n4908 ) | ( n4737 & n4908 ) ;
  assign n4911 = ( n4723 & ~n4909 ) | ( n4723 & n4910 ) | ( ~n4909 & n4910 ) ;
  assign n4912 = ( ~x107 & x108 ) | ( ~x107 & n4522 ) | ( x108 & n4522 ) ;
  assign n4913 = ( x107 & x108 ) | ( x107 & n4522 ) | ( x108 & n4522 ) ;
  assign n4914 = ( x107 & n4912 ) | ( x107 & ~n4913 ) | ( n4912 & ~n4913 ) ;
  assign n4915 = x0 & n4914 ;
  assign n4916 = ( x1 & x2 ) | ( x1 & n4915 ) | ( x2 & n4915 ) ;
  assign n4917 = x107 & n172 ;
  assign n4918 = ( ~x106 & n135 ) | ( ~x106 & n174 ) | ( n135 & n174 ) ;
  assign n4919 = n4917 | n4918 ;
  assign n4920 = x108 & n147 ;
  assign n4921 = n4919 | n4920 ;
  assign n4922 = n4916 | n4921 ;
  assign n4923 = n4916 & n4921 ;
  assign n4924 = n4922 & ~n4923 ;
  assign n4925 = ( n4725 & ~n4911 ) | ( n4725 & n4924 ) | ( ~n4911 & n4924 ) ;
  assign n4926 = ( n4725 & n4911 ) | ( n4725 & n4924 ) | ( n4911 & n4924 ) ;
  assign n4927 = ( n4911 & n4925 ) | ( n4911 & ~n4926 ) | ( n4925 & ~n4926 ) ;
  assign n4928 = ( ~x108 & x109 ) | ( ~x108 & n4913 ) | ( x109 & n4913 ) ;
  assign n4929 = ( x108 & x109 ) | ( x108 & n4913 ) | ( x109 & n4913 ) ;
  assign n4930 = ( x108 & n4928 ) | ( x108 & ~n4929 ) | ( n4928 & ~n4929 ) ;
  assign n4931 = x0 & n4930 ;
  assign n4932 = ( x1 & x2 ) | ( x1 & n4931 ) | ( x2 & n4931 ) ;
  assign n4933 = x108 & n172 ;
  assign n4934 = x109 | n4933 ;
  assign n4935 = ( n147 & n4933 ) | ( n147 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4936 = ( ~x107 & n135 ) | ( ~x107 & n174 ) | ( n135 & n174 ) ;
  assign n4937 = n4935 | n4936 ;
  assign n4938 = n4932 | n4937 ;
  assign n4939 = n4932 & n4937 ;
  assign n4940 = n4938 & ~n4939 ;
  assign n4941 = n449 & n3264 ;
  assign n4942 = x11 & n4941 ;
  assign n4943 = x100 & n456 ;
  assign n4944 = x99 & n453 ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = x98 & n536 ;
  assign n4947 = n4945 | n4946 ;
  assign n4948 = ( ~x11 & n4941 ) | ( ~x11 & n4947 ) | ( n4941 & n4947 ) ;
  assign n4949 = x11 & ~n4947 ;
  assign n4950 = ( ~n4942 & n4948 ) | ( ~n4942 & n4949 ) | ( n4948 & n4949 ) ;
  assign n4951 = n874 & n2476 ;
  assign n4952 = x17 & n4951 ;
  assign n4953 = x94 & n881 ;
  assign n4954 = x93 & n878 ;
  assign n4955 = n4953 | n4954 ;
  assign n4956 = x92 & n959 ;
  assign n4957 = n4955 | n4956 ;
  assign n4958 = ( ~x17 & n4951 ) | ( ~x17 & n4957 ) | ( n4951 & n4957 ) ;
  assign n4959 = x17 & ~n4957 ;
  assign n4960 = ( ~n4952 & n4958 ) | ( ~n4952 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4961 = n1427 & n1602 ;
  assign n4962 = x23 & n4961 ;
  assign n4963 = x88 & n1434 ;
  assign n4964 = x87 & n1431 ;
  assign n4965 = n4963 | n4964 ;
  assign n4966 = x86 & n1531 ;
  assign n4967 = n4965 | n4966 ;
  assign n4968 = ( ~x23 & n4961 ) | ( ~x23 & n4967 ) | ( n4961 & n4967 ) ;
  assign n4969 = x23 & ~n4967 ;
  assign n4970 = ( ~n4962 & n4968 ) | ( ~n4962 & n4969 ) | ( n4968 & n4969 ) ;
  assign n4971 = n1006 & n2137 ;
  assign n4972 = x29 & n4971 ;
  assign n4973 = x82 & n2144 ;
  assign n4974 = x81 & n2141 ;
  assign n4975 = n4973 | n4974 ;
  assign n4976 = x80 & n2267 ;
  assign n4977 = n4975 | n4976 ;
  assign n4978 = ( ~x29 & n4971 ) | ( ~x29 & n4977 ) | ( n4971 & n4977 ) ;
  assign n4979 = x29 & ~n4977 ;
  assign n4980 = ( ~n4972 & n4978 ) | ( ~n4972 & n4979 ) | ( n4978 & n4979 ) ;
  assign n4981 = n565 & n2982 ;
  assign n4982 = x35 & n4981 ;
  assign n4983 = x76 & n2989 ;
  assign n4984 = x75 & n2986 ;
  assign n4985 = n4983 | n4984 ;
  assign n4986 = x74 & n3159 ;
  assign n4987 = n4985 | n4986 ;
  assign n4988 = ( ~x35 & n4981 ) | ( ~x35 & n4987 ) | ( n4981 & n4987 ) ;
  assign n4989 = x35 & ~n4987 ;
  assign n4990 = ( ~n4982 & n4988 ) | ( ~n4982 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4991 = n276 & n4020 ;
  assign n4992 = x41 & n4991 ;
  assign n4993 = x70 & n4027 ;
  assign n4994 = x69 & n4024 ;
  assign n4995 = n4993 | n4994 ;
  assign n4996 = x68 & n4223 ;
  assign n4997 = n4995 | n4996 ;
  assign n4998 = ( ~x41 & n4991 ) | ( ~x41 & n4997 ) | ( n4991 & n4997 ) ;
  assign n4999 = x41 & ~n4997 ;
  assign n5000 = ( ~n4992 & n4998 ) | ( ~n4992 & n4999 ) | ( n4998 & n4999 ) ;
  assign n5001 = x67 & n4791 ;
  assign n5002 = x66 & n4621 ;
  assign n5003 = n5001 | n5002 ;
  assign n5004 = x65 & n4795 ;
  assign n5005 = n5003 | n5004 ;
  assign n5006 = n169 & n4625 ;
  assign n5007 = n5005 | n5006 ;
  assign n5008 = x44 & x45 ;
  assign n5009 = x44 | x45 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = x64 & n5010 ;
  assign n5012 = ( x44 & n4797 ) | ( x44 & n4799 ) | ( n4797 & n4799 ) ;
  assign n5013 = ( ~n5007 & n5011 ) | ( ~n5007 & n5012 ) | ( n5011 & n5012 ) ;
  assign n5014 = x44 & ~n5007 ;
  assign n5015 = ( n5007 & ~n5012 ) | ( n5007 & n5014 ) | ( ~n5012 & n5014 ) ;
  assign n5016 = ( n5011 & n5014 ) | ( n5011 & n5015 ) | ( n5014 & n5015 ) ;
  assign n5017 = ( n5013 & n5015 ) | ( n5013 & ~n5016 ) | ( n5015 & ~n5016 ) ;
  assign n5018 = ( n4813 & n5000 ) | ( n4813 & n5017 ) | ( n5000 & n5017 ) ;
  assign n5019 = ( ~n4813 & n5000 ) | ( ~n4813 & n5017 ) | ( n5000 & n5017 ) ;
  assign n5020 = ( n4813 & ~n5018 ) | ( n4813 & n5019 ) | ( ~n5018 & n5019 ) ;
  assign n5021 = n388 & n3492 ;
  assign n5022 = x38 & n5021 ;
  assign n5023 = x73 & n3499 ;
  assign n5024 = x72 & n3496 ;
  assign n5025 = n5023 | n5024 ;
  assign n5026 = x71 & n3662 ;
  assign n5027 = n5025 | n5026 ;
  assign n5028 = ( ~x38 & n5021 ) | ( ~x38 & n5027 ) | ( n5021 & n5027 ) ;
  assign n5029 = x38 & ~n5027 ;
  assign n5030 = ( ~n5022 & n5028 ) | ( ~n5022 & n5029 ) | ( n5028 & n5029 ) ;
  assign n5031 = ( n4827 & ~n5020 ) | ( n4827 & n5030 ) | ( ~n5020 & n5030 ) ;
  assign n5032 = ( n4827 & n5020 ) | ( n4827 & n5030 ) | ( n5020 & n5030 ) ;
  assign n5033 = ( n5020 & n5031 ) | ( n5020 & ~n5032 ) | ( n5031 & ~n5032 ) ;
  assign n5034 = ( n4829 & n4990 ) | ( n4829 & n5033 ) | ( n4990 & n5033 ) ;
  assign n5035 = ( ~n4829 & n4990 ) | ( ~n4829 & n5033 ) | ( n4990 & n5033 ) ;
  assign n5036 = ( n4829 & ~n5034 ) | ( n4829 & n5035 ) | ( ~n5034 & n5035 ) ;
  assign n5037 = n823 & n2545 ;
  assign n5038 = x32 & n5037 ;
  assign n5039 = x79 & n2552 ;
  assign n5040 = x78 & n2549 ;
  assign n5041 = n5039 | n5040 ;
  assign n5042 = x77 & n2696 ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = ( ~x32 & n5037 ) | ( ~x32 & n5043 ) | ( n5037 & n5043 ) ;
  assign n5045 = x32 & ~n5043 ;
  assign n5046 = ( ~n5038 & n5044 ) | ( ~n5038 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5047 = ( n4843 & ~n5036 ) | ( n4843 & n5046 ) | ( ~n5036 & n5046 ) ;
  assign n5048 = ( n4843 & n5036 ) | ( n4843 & n5046 ) | ( n5036 & n5046 ) ;
  assign n5049 = ( n5036 & n5047 ) | ( n5036 & ~n5048 ) | ( n5047 & ~n5048 ) ;
  assign n5050 = ( n4845 & n4980 ) | ( n4845 & n5049 ) | ( n4980 & n5049 ) ;
  assign n5051 = ( ~n4845 & n4980 ) | ( ~n4845 & n5049 ) | ( n4980 & n5049 ) ;
  assign n5052 = ( n4845 & ~n5050 ) | ( n4845 & n5051 ) | ( ~n5050 & n5051 ) ;
  assign n5053 = n1368 & n1755 ;
  assign n5054 = x26 & n5053 ;
  assign n5055 = x85 & n1762 ;
  assign n5056 = x84 & n1759 ;
  assign n5057 = n5055 | n5056 ;
  assign n5058 = x83 & n1895 ;
  assign n5059 = n5057 | n5058 ;
  assign n5060 = ( ~x26 & n5053 ) | ( ~x26 & n5059 ) | ( n5053 & n5059 ) ;
  assign n5061 = x26 & ~n5059 ;
  assign n5062 = ( ~n5054 & n5060 ) | ( ~n5054 & n5061 ) | ( n5060 & n5061 ) ;
  assign n5063 = ( n4859 & ~n5052 ) | ( n4859 & n5062 ) | ( ~n5052 & n5062 ) ;
  assign n5064 = ( n4859 & n5052 ) | ( n4859 & n5062 ) | ( n5052 & n5062 ) ;
  assign n5065 = ( n5052 & n5063 ) | ( n5052 & ~n5064 ) | ( n5063 & ~n5064 ) ;
  assign n5066 = ( n4861 & n4970 ) | ( n4861 & n5065 ) | ( n4970 & n5065 ) ;
  assign n5067 = ( ~n4861 & n4970 ) | ( ~n4861 & n5065 ) | ( n4970 & n5065 ) ;
  assign n5068 = ( n4861 & ~n5066 ) | ( n4861 & n5067 ) | ( ~n5066 & n5067 ) ;
  assign n5069 = n1146 & n1959 ;
  assign n5070 = x20 & n5069 ;
  assign n5071 = x91 & n1153 ;
  assign n5072 = x90 & n1150 ;
  assign n5073 = n5071 | n5072 ;
  assign n5074 = x89 & n1217 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = ( ~x20 & n5069 ) | ( ~x20 & n5075 ) | ( n5069 & n5075 ) ;
  assign n5077 = x20 & ~n5075 ;
  assign n5078 = ( ~n5070 & n5076 ) | ( ~n5070 & n5077 ) | ( n5076 & n5077 ) ;
  assign n5079 = ( n4875 & ~n5068 ) | ( n4875 & n5078 ) | ( ~n5068 & n5078 ) ;
  assign n5080 = ( n4875 & n5068 ) | ( n4875 & n5078 ) | ( n5068 & n5078 ) ;
  assign n5081 = ( n5068 & n5079 ) | ( n5068 & ~n5080 ) | ( n5079 & ~n5080 ) ;
  assign n5082 = ( ~n4877 & n4960 ) | ( ~n4877 & n5081 ) | ( n4960 & n5081 ) ;
  assign n5083 = ( n4877 & n4960 ) | ( n4877 & n5081 ) | ( n4960 & n5081 ) ;
  assign n5084 = ( n4877 & n5082 ) | ( n4877 & ~n5083 ) | ( n5082 & ~n5083 ) ;
  assign n5085 = x97 & n656 ;
  assign n5086 = x95 & n744 ;
  assign n5087 = n5085 | n5086 ;
  assign n5088 = n649 | n5087 ;
  assign n5089 = ( n2788 & n5087 ) | ( n2788 & n5088 ) | ( n5087 & n5088 ) ;
  assign n5090 = x96 & n653 ;
  assign n5091 = ( ~x14 & n5089 ) | ( ~x14 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5092 = ( x14 & ~n5089 ) | ( x14 & n5090 ) | ( ~n5089 & n5090 ) ;
  assign n5093 = ~n5090 & n5092 ;
  assign n5094 = n5091 | n5093 ;
  assign n5095 = ( n4891 & ~n5084 ) | ( n4891 & n5094 ) | ( ~n5084 & n5094 ) ;
  assign n5096 = ( n4891 & n5084 ) | ( n4891 & n5094 ) | ( n5084 & n5094 ) ;
  assign n5097 = ( n5084 & n5095 ) | ( n5084 & ~n5096 ) | ( n5095 & ~n5096 ) ;
  assign n5098 = ( ~n4904 & n4950 ) | ( ~n4904 & n5097 ) | ( n4950 & n5097 ) ;
  assign n5099 = ( n4904 & n4950 ) | ( n4904 & n5097 ) | ( n4950 & n5097 ) ;
  assign n5100 = ( n4904 & n5098 ) | ( n4904 & ~n5099 ) | ( n5098 & ~n5099 ) ;
  assign n5101 = n301 & n3941 ;
  assign n5102 = x8 & n5101 ;
  assign n5103 = x103 & n309 ;
  assign n5104 = x102 & n306 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = x101 & n359 ;
  assign n5107 = n5105 | n5106 ;
  assign n5108 = ( ~x8 & n5101 ) | ( ~x8 & n5107 ) | ( n5101 & n5107 ) ;
  assign n5109 = x8 & ~n5107 ;
  assign n5110 = ( ~n5102 & n5108 ) | ( ~n5102 & n5109 ) | ( n5108 & n5109 ) ;
  assign n5111 = ( n4906 & ~n5100 ) | ( n4906 & n5110 ) | ( ~n5100 & n5110 ) ;
  assign n5112 = ( n4906 & n5100 ) | ( n4906 & n5110 ) | ( n5100 & n5110 ) ;
  assign n5113 = ( n5100 & n5111 ) | ( n5100 & ~n5112 ) | ( n5111 & ~n5112 ) ;
  assign n5114 = n206 & n4331 ;
  assign n5115 = x5 & n5114 ;
  assign n5116 = x106 & n205 ;
  assign n5117 = x105 & n201 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = x104 & n221 ;
  assign n5120 = n5118 | n5119 ;
  assign n5121 = ( ~x5 & n5114 ) | ( ~x5 & n5120 ) | ( n5114 & n5120 ) ;
  assign n5122 = x5 & ~n5120 ;
  assign n5123 = ( ~n5115 & n5121 ) | ( ~n5115 & n5122 ) | ( n5121 & n5122 ) ;
  assign n5124 = ( n4909 & ~n5113 ) | ( n4909 & n5123 ) | ( ~n5113 & n5123 ) ;
  assign n5125 = ( n4909 & n5113 ) | ( n4909 & n5123 ) | ( n5113 & n5123 ) ;
  assign n5126 = ( n5113 & n5124 ) | ( n5113 & ~n5125 ) | ( n5124 & ~n5125 ) ;
  assign n5127 = ( n4926 & n4940 ) | ( n4926 & n5126 ) | ( n4940 & n5126 ) ;
  assign n5128 = ( ~n4926 & n4940 ) | ( ~n4926 & n5126 ) | ( n4940 & n5126 ) ;
  assign n5129 = ( n4926 & ~n5127 ) | ( n4926 & n5128 ) | ( ~n5127 & n5128 ) ;
  assign n5130 = n206 & n4523 ;
  assign n5131 = x5 & n5130 ;
  assign n5132 = x107 & n205 ;
  assign n5133 = x106 & n201 ;
  assign n5134 = n5132 | n5133 ;
  assign n5135 = x105 & n221 ;
  assign n5136 = n5134 | n5135 ;
  assign n5137 = ( ~x5 & n5130 ) | ( ~x5 & n5136 ) | ( n5130 & n5136 ) ;
  assign n5138 = x5 & ~n5136 ;
  assign n5139 = ( ~n5131 & n5137 ) | ( ~n5131 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5140 = n301 & n3957 ;
  assign n5141 = x8 & n5140 ;
  assign n5142 = x104 & n309 ;
  assign n5143 = x103 & n306 ;
  assign n5144 = n5142 | n5143 ;
  assign n5145 = x102 & n359 ;
  assign n5146 = n5144 | n5145 ;
  assign n5147 = ( ~x8 & n5140 ) | ( ~x8 & n5146 ) | ( n5140 & n5146 ) ;
  assign n5148 = x8 & ~n5146 ;
  assign n5149 = ( ~n5141 & n5147 ) | ( ~n5141 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5150 = n449 & n3591 ;
  assign n5151 = x11 & n5150 ;
  assign n5152 = x101 & n456 ;
  assign n5153 = x100 & n453 ;
  assign n5154 = n5152 | n5153 ;
  assign n5155 = x99 & n536 ;
  assign n5156 = n5154 | n5155 ;
  assign n5157 = ( ~x11 & n5150 ) | ( ~x11 & n5156 ) | ( n5150 & n5156 ) ;
  assign n5158 = x11 & ~n5156 ;
  assign n5159 = ( ~n5151 & n5157 ) | ( ~n5151 & n5158 ) | ( n5157 & n5158 ) ;
  assign n5160 = n649 & n2939 ;
  assign n5161 = x14 & n5160 ;
  assign n5162 = x98 & n656 ;
  assign n5163 = x97 & n653 ;
  assign n5164 = n5162 | n5163 ;
  assign n5165 = x96 & n744 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = ( ~x14 & n5160 ) | ( ~x14 & n5166 ) | ( n5160 & n5166 ) ;
  assign n5168 = x14 & ~n5166 ;
  assign n5169 = ( ~n5161 & n5167 ) | ( ~n5161 & n5168 ) | ( n5167 & n5168 ) ;
  assign n5170 = n874 & n2492 ;
  assign n5171 = x17 & n5170 ;
  assign n5172 = x95 & n881 ;
  assign n5173 = x94 & n878 ;
  assign n5174 = n5172 | n5173 ;
  assign n5175 = x93 & n959 ;
  assign n5176 = n5174 | n5175 ;
  assign n5177 = ( ~x17 & n5170 ) | ( ~x17 & n5176 ) | ( n5170 & n5176 ) ;
  assign n5178 = x17 & ~n5176 ;
  assign n5179 = ( ~n5171 & n5177 ) | ( ~n5171 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5180 = n1427 & n1822 ;
  assign n5181 = x23 & n5180 ;
  assign n5182 = x89 & n1434 ;
  assign n5183 = x88 & n1431 ;
  assign n5184 = n5182 | n5183 ;
  assign n5185 = x87 & n1531 ;
  assign n5186 = n5184 | n5185 ;
  assign n5187 = ( ~x23 & n5180 ) | ( ~x23 & n5186 ) | ( n5180 & n5186 ) ;
  assign n5188 = x23 & ~n5186 ;
  assign n5189 = ( ~n5181 & n5187 ) | ( ~n5181 & n5188 ) | ( n5187 & n5188 ) ;
  assign n5190 = n1093 & n2137 ;
  assign n5191 = x29 & n5190 ;
  assign n5192 = x83 & n2144 ;
  assign n5193 = x82 & n2141 ;
  assign n5194 = n5192 | n5193 ;
  assign n5195 = x81 & n2267 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = ( ~x29 & n5190 ) | ( ~x29 & n5196 ) | ( n5190 & n5196 ) ;
  assign n5198 = x29 & ~n5196 ;
  assign n5199 = ( ~n5191 & n5197 ) | ( ~n5191 & n5198 ) | ( n5197 & n5198 ) ;
  assign n5200 = n626 & n2982 ;
  assign n5201 = x35 & n5200 ;
  assign n5202 = x77 & n2989 ;
  assign n5203 = x76 & n2986 ;
  assign n5204 = n5202 | n5203 ;
  assign n5205 = x75 & n3159 ;
  assign n5206 = n5204 | n5205 ;
  assign n5207 = ( ~x35 & n5200 ) | ( ~x35 & n5206 ) | ( n5200 & n5206 ) ;
  assign n5208 = x35 & ~n5206 ;
  assign n5209 = ( ~n5201 & n5207 ) | ( ~n5201 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5210 = n193 & n4625 ;
  assign n5211 = x44 & n5210 ;
  assign n5212 = x68 & n4791 ;
  assign n5213 = x67 & n4621 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = x66 & n4795 ;
  assign n5216 = n5214 | n5215 ;
  assign n5217 = ( ~x44 & n5210 ) | ( ~x44 & n5216 ) | ( n5210 & n5216 ) ;
  assign n5218 = x44 & ~n5216 ;
  assign n5219 = ( ~n5211 & n5217 ) | ( ~n5211 & n5218 ) | ( n5217 & n5218 ) ;
  assign n5220 = x46 & x47 ;
  assign n5221 = x46 | x47 ;
  assign n5222 = ~n5220 & n5221 ;
  assign n5223 = n5010 & n5222 ;
  assign n5224 = n302 & n5223 ;
  assign n5225 = ~x44 & x46 ;
  assign n5226 = x45 & x46 ;
  assign n5227 = ( n5008 & n5225 ) | ( n5008 & ~n5226 ) | ( n5225 & ~n5226 ) ;
  assign n5228 = x64 & n5227 ;
  assign n5229 = n5224 | n5228 ;
  assign n5230 = ( n5010 & n5220 ) | ( n5010 & ~n5221 ) | ( n5220 & ~n5221 ) ;
  assign n5231 = x65 & n5230 ;
  assign n5232 = n5229 | n5231 ;
  assign n5233 = n5011 | n5232 ;
  assign n5234 = ( x47 & n5011 ) | ( x47 & ~n5232 ) | ( n5011 & ~n5232 ) ;
  assign n5235 = x47 & ~n5232 ;
  assign n5236 = ( n5233 & ~n5234 ) | ( n5233 & n5235 ) | ( ~n5234 & n5235 ) ;
  assign n5237 = ( ~n5016 & n5219 ) | ( ~n5016 & n5236 ) | ( n5219 & n5236 ) ;
  assign n5238 = ( n5016 & n5219 ) | ( n5016 & n5236 ) | ( n5219 & n5236 ) ;
  assign n5239 = ( n5016 & n5237 ) | ( n5016 & ~n5238 ) | ( n5237 & ~n5238 ) ;
  assign n5240 = n322 & n4020 ;
  assign n5241 = x41 & n5240 ;
  assign n5242 = x71 & n4027 ;
  assign n5243 = x70 & n4024 ;
  assign n5244 = n5242 | n5243 ;
  assign n5245 = x69 & n4223 ;
  assign n5246 = n5244 | n5245 ;
  assign n5247 = ( ~x41 & n5240 ) | ( ~x41 & n5246 ) | ( n5240 & n5246 ) ;
  assign n5248 = x41 & ~n5246 ;
  assign n5249 = ( ~n5241 & n5247 ) | ( ~n5241 & n5248 ) | ( n5247 & n5248 ) ;
  assign n5250 = ( n5018 & n5239 ) | ( n5018 & n5249 ) | ( n5239 & n5249 ) ;
  assign n5251 = ( ~n5018 & n5239 ) | ( ~n5018 & n5249 ) | ( n5239 & n5249 ) ;
  assign n5252 = ( n5018 & ~n5250 ) | ( n5018 & n5251 ) | ( ~n5250 & n5251 ) ;
  assign n5253 = n436 & n3492 ;
  assign n5254 = x38 & n5253 ;
  assign n5255 = x74 & n3499 ;
  assign n5256 = x73 & n3496 ;
  assign n5257 = n5255 | n5256 ;
  assign n5258 = x72 & n3662 ;
  assign n5259 = n5257 | n5258 ;
  assign n5260 = ( ~x38 & n5253 ) | ( ~x38 & n5259 ) | ( n5253 & n5259 ) ;
  assign n5261 = x38 & ~n5259 ;
  assign n5262 = ( ~n5254 & n5260 ) | ( ~n5254 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = ( n5032 & ~n5252 ) | ( n5032 & n5262 ) | ( ~n5252 & n5262 ) ;
  assign n5264 = ( n5032 & n5252 ) | ( n5032 & n5262 ) | ( n5252 & n5262 ) ;
  assign n5265 = ( n5252 & n5263 ) | ( n5252 & ~n5264 ) | ( n5263 & ~n5264 ) ;
  assign n5266 = ( n5034 & n5209 ) | ( n5034 & n5265 ) | ( n5209 & n5265 ) ;
  assign n5267 = ( ~n5034 & n5209 ) | ( ~n5034 & n5265 ) | ( n5209 & n5265 ) ;
  assign n5268 = ( n5034 & ~n5266 ) | ( n5034 & n5267 ) | ( ~n5266 & n5267 ) ;
  assign n5269 = n840 & n2545 ;
  assign n5270 = x32 & n5269 ;
  assign n5271 = x80 & n2552 ;
  assign n5272 = x79 & n2549 ;
  assign n5273 = n5271 | n5272 ;
  assign n5274 = x78 & n2696 ;
  assign n5275 = n5273 | n5274 ;
  assign n5276 = ( ~x32 & n5269 ) | ( ~x32 & n5275 ) | ( n5269 & n5275 ) ;
  assign n5277 = x32 & ~n5275 ;
  assign n5278 = ( ~n5270 & n5276 ) | ( ~n5270 & n5277 ) | ( n5276 & n5277 ) ;
  assign n5279 = ( n5048 & ~n5268 ) | ( n5048 & n5278 ) | ( ~n5268 & n5278 ) ;
  assign n5280 = ( n5048 & n5268 ) | ( n5048 & n5278 ) | ( n5268 & n5278 ) ;
  assign n5281 = ( n5268 & n5279 ) | ( n5268 & ~n5280 ) | ( n5279 & ~n5280 ) ;
  assign n5282 = ( n5050 & n5199 ) | ( n5050 & n5281 ) | ( n5199 & n5281 ) ;
  assign n5283 = ( ~n5050 & n5199 ) | ( ~n5050 & n5281 ) | ( n5199 & n5281 ) ;
  assign n5284 = ( n5050 & ~n5282 ) | ( n5050 & n5283 ) | ( ~n5282 & n5283 ) ;
  assign n5285 = n1384 & n1755 ;
  assign n5286 = x26 & n5285 ;
  assign n5287 = x86 & n1762 ;
  assign n5288 = x85 & n1759 ;
  assign n5289 = n5287 | n5288 ;
  assign n5290 = x84 & n1895 ;
  assign n5291 = n5289 | n5290 ;
  assign n5292 = ( ~x26 & n5285 ) | ( ~x26 & n5291 ) | ( n5285 & n5291 ) ;
  assign n5293 = x26 & ~n5291 ;
  assign n5294 = ( ~n5286 & n5292 ) | ( ~n5286 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5295 = ( n5064 & ~n5284 ) | ( n5064 & n5294 ) | ( ~n5284 & n5294 ) ;
  assign n5296 = ( n5064 & n5284 ) | ( n5064 & n5294 ) | ( n5284 & n5294 ) ;
  assign n5297 = ( n5284 & n5295 ) | ( n5284 & ~n5296 ) | ( n5295 & ~n5296 ) ;
  assign n5298 = ( n5066 & n5189 ) | ( n5066 & n5297 ) | ( n5189 & n5297 ) ;
  assign n5299 = ( ~n5066 & n5189 ) | ( ~n5066 & n5297 ) | ( n5189 & n5297 ) ;
  assign n5300 = ( n5066 & ~n5298 ) | ( n5066 & n5299 ) | ( ~n5298 & n5299 ) ;
  assign n5301 = n1146 & n2083 ;
  assign n5302 = x20 & n5301 ;
  assign n5303 = x92 & n1153 ;
  assign n5304 = x91 & n1150 ;
  assign n5305 = n5303 | n5304 ;
  assign n5306 = x90 & n1217 ;
  assign n5307 = n5305 | n5306 ;
  assign n5308 = ( ~x20 & n5301 ) | ( ~x20 & n5307 ) | ( n5301 & n5307 ) ;
  assign n5309 = x20 & ~n5307 ;
  assign n5310 = ( ~n5302 & n5308 ) | ( ~n5302 & n5309 ) | ( n5308 & n5309 ) ;
  assign n5311 = ( n5080 & ~n5300 ) | ( n5080 & n5310 ) | ( ~n5300 & n5310 ) ;
  assign n5312 = ( n5080 & n5300 ) | ( n5080 & n5310 ) | ( n5300 & n5310 ) ;
  assign n5313 = ( n5300 & n5311 ) | ( n5300 & ~n5312 ) | ( n5311 & ~n5312 ) ;
  assign n5314 = ( n5083 & n5179 ) | ( n5083 & n5313 ) | ( n5179 & n5313 ) ;
  assign n5315 = ( ~n5083 & n5179 ) | ( ~n5083 & n5313 ) | ( n5179 & n5313 ) ;
  assign n5316 = ( n5083 & ~n5314 ) | ( n5083 & n5315 ) | ( ~n5314 & n5315 ) ;
  assign n5317 = ( n5096 & n5169 ) | ( n5096 & n5316 ) | ( n5169 & n5316 ) ;
  assign n5318 = ( ~n5096 & n5169 ) | ( ~n5096 & n5316 ) | ( n5169 & n5316 ) ;
  assign n5319 = ( n5096 & ~n5317 ) | ( n5096 & n5318 ) | ( ~n5317 & n5318 ) ;
  assign n5320 = ( n5099 & ~n5159 ) | ( n5099 & n5319 ) | ( ~n5159 & n5319 ) ;
  assign n5321 = ( n5099 & n5159 ) | ( n5099 & n5319 ) | ( n5159 & n5319 ) ;
  assign n5322 = ( n5159 & n5320 ) | ( n5159 & ~n5321 ) | ( n5320 & ~n5321 ) ;
  assign n5323 = ( n5112 & n5149 ) | ( n5112 & n5322 ) | ( n5149 & n5322 ) ;
  assign n5324 = ( ~n5112 & n5149 ) | ( ~n5112 & n5322 ) | ( n5149 & n5322 ) ;
  assign n5325 = ( n5112 & ~n5323 ) | ( n5112 & n5324 ) | ( ~n5323 & n5324 ) ;
  assign n5326 = ( n5125 & n5139 ) | ( n5125 & n5325 ) | ( n5139 & n5325 ) ;
  assign n5327 = ( ~n5125 & n5139 ) | ( ~n5125 & n5325 ) | ( n5139 & n5325 ) ;
  assign n5328 = ( n5125 & ~n5326 ) | ( n5125 & n5327 ) | ( ~n5326 & n5327 ) ;
  assign n5329 = ( ~x109 & x110 ) | ( ~x109 & n4929 ) | ( x110 & n4929 ) ;
  assign n5330 = ( x109 & x110 ) | ( x109 & n4929 ) | ( x110 & n4929 ) ;
  assign n5331 = ( x109 & n5329 ) | ( x109 & ~n5330 ) | ( n5329 & ~n5330 ) ;
  assign n5332 = x0 & n5331 ;
  assign n5333 = ( x1 & x2 ) | ( x1 & n5332 ) | ( x2 & n5332 ) ;
  assign n5334 = x109 & n172 ;
  assign n5335 = ( ~x108 & n135 ) | ( ~x108 & n174 ) | ( n135 & n174 ) ;
  assign n5336 = n5334 | n5335 ;
  assign n5337 = x110 & n147 ;
  assign n5338 = n5336 | n5337 ;
  assign n5339 = n5333 | n5338 ;
  assign n5340 = n5333 & n5338 ;
  assign n5341 = n5339 & ~n5340 ;
  assign n5342 = ( n5127 & ~n5328 ) | ( n5127 & n5341 ) | ( ~n5328 & n5341 ) ;
  assign n5343 = ( n5127 & n5328 ) | ( n5127 & n5341 ) | ( n5328 & n5341 ) ;
  assign n5344 = ( n5328 & n5342 ) | ( n5328 & ~n5343 ) | ( n5342 & ~n5343 ) ;
  assign n5345 = ( ~x110 & x111 ) | ( ~x110 & n5330 ) | ( x111 & n5330 ) ;
  assign n5346 = ( x110 & x111 ) | ( x110 & n5330 ) | ( x111 & n5330 ) ;
  assign n5347 = ( x110 & n5345 ) | ( x110 & ~n5346 ) | ( n5345 & ~n5346 ) ;
  assign n5348 = x0 & n5347 ;
  assign n5349 = ( x1 & x2 ) | ( x1 & n5348 ) | ( x2 & n5348 ) ;
  assign n5350 = x110 & n172 ;
  assign n5351 = x111 | n5350 ;
  assign n5352 = ( n147 & n5350 ) | ( n147 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5353 = ( ~x109 & n135 ) | ( ~x109 & n174 ) | ( n135 & n174 ) ;
  assign n5354 = n5352 | n5353 ;
  assign n5355 = n5349 | n5354 ;
  assign n5356 = n5349 & n5354 ;
  assign n5357 = n5355 & ~n5356 ;
  assign n5358 = n301 & n4145 ;
  assign n5359 = x8 & n5358 ;
  assign n5360 = x105 & n309 ;
  assign n5361 = x104 & n306 ;
  assign n5362 = n5360 | n5361 ;
  assign n5363 = x103 & n359 ;
  assign n5364 = n5362 | n5363 ;
  assign n5365 = ( ~x8 & n5358 ) | ( ~x8 & n5364 ) | ( n5358 & n5364 ) ;
  assign n5366 = x8 & ~n5364 ;
  assign n5367 = ( ~n5359 & n5365 ) | ( ~n5359 & n5366 ) | ( n5365 & n5366 ) ;
  assign n5368 = n649 & n3248 ;
  assign n5369 = x14 & n5368 ;
  assign n5370 = x99 & n656 ;
  assign n5371 = x98 & n653 ;
  assign n5372 = n5370 | n5371 ;
  assign n5373 = x97 & n744 ;
  assign n5374 = n5372 | n5373 ;
  assign n5375 = ( ~x14 & n5368 ) | ( ~x14 & n5374 ) | ( n5368 & n5374 ) ;
  assign n5376 = x14 & ~n5374 ;
  assign n5377 = ( ~n5369 & n5375 ) | ( ~n5369 & n5376 ) | ( n5375 & n5376 ) ;
  assign n5378 = n1427 & n1838 ;
  assign n5379 = x23 & n5378 ;
  assign n5380 = x90 & n1434 ;
  assign n5381 = x89 & n1431 ;
  assign n5382 = n5380 | n5381 ;
  assign n5383 = x88 & n1531 ;
  assign n5384 = n5382 | n5383 ;
  assign n5385 = ( ~x23 & n5378 ) | ( ~x23 & n5384 ) | ( n5378 & n5384 ) ;
  assign n5386 = x23 & ~n5384 ;
  assign n5387 = ( ~n5379 & n5385 ) | ( ~n5379 & n5386 ) | ( n5385 & n5386 ) ;
  assign n5388 = n1494 & n1755 ;
  assign n5389 = x26 & n5388 ;
  assign n5390 = x87 & n1762 ;
  assign n5391 = x86 & n1759 ;
  assign n5392 = n5390 | n5391 ;
  assign n5393 = x85 & n1895 ;
  assign n5394 = n5392 | n5393 ;
  assign n5395 = ( ~x26 & n5388 ) | ( ~x26 & n5394 ) | ( n5388 & n5394 ) ;
  assign n5396 = x26 & ~n5394 ;
  assign n5397 = ( ~n5389 & n5395 ) | ( ~n5389 & n5396 ) | ( n5395 & n5396 ) ;
  assign n5398 = n990 & n2545 ;
  assign n5399 = x32 & n5398 ;
  assign n5400 = x81 & n2552 ;
  assign n5401 = x80 & n2549 ;
  assign n5402 = n5400 | n5401 ;
  assign n5403 = x79 & n2696 ;
  assign n5404 = n5402 | n5403 ;
  assign n5405 = ( ~x32 & n5398 ) | ( ~x32 & n5404 ) | ( n5398 & n5404 ) ;
  assign n5406 = x32 & ~n5404 ;
  assign n5407 = ( ~n5399 & n5405 ) | ( ~n5399 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5408 = n508 & n3492 ;
  assign n5409 = x38 & n5408 ;
  assign n5410 = x75 & n3499 ;
  assign n5411 = x74 & n3496 ;
  assign n5412 = n5410 | n5411 ;
  assign n5413 = x73 & n3662 ;
  assign n5414 = n5412 | n5413 ;
  assign n5415 = ( ~x38 & n5408 ) | ( ~x38 & n5414 ) | ( n5408 & n5414 ) ;
  assign n5416 = x38 & ~n5414 ;
  assign n5417 = ( ~n5409 & n5415 ) | ( ~n5409 & n5416 ) | ( n5415 & n5416 ) ;
  assign n5418 = n240 & n4625 ;
  assign n5419 = x44 & n5418 ;
  assign n5420 = x69 & n4791 ;
  assign n5421 = x68 & n4621 ;
  assign n5422 = n5420 | n5421 ;
  assign n5423 = x67 & n4795 ;
  assign n5424 = n5422 | n5423 ;
  assign n5425 = ( ~x44 & n5418 ) | ( ~x44 & n5424 ) | ( n5418 & n5424 ) ;
  assign n5426 = x44 & ~n5424 ;
  assign n5427 = ( ~n5419 & n5425 ) | ( ~n5419 & n5426 ) | ( n5425 & n5426 ) ;
  assign n5428 = x65 & n5227 ;
  assign n5429 = n226 & n5223 ;
  assign n5430 = n5428 | n5429 ;
  assign n5431 = x66 & n5230 ;
  assign n5432 = n5430 | n5431 ;
  assign n5433 = ~n5010 & n5222 ;
  assign n5434 = ~n5227 & n5433 ;
  assign n5435 = x64 & n5434 ;
  assign n5436 = n5432 | n5435 ;
  assign n5437 = ~x47 & n5436 ;
  assign n5438 = ( x47 & n5233 ) | ( x47 & n5436 ) | ( n5233 & n5436 ) ;
  assign n5439 = n5233 & n5436 ;
  assign n5440 = ( n5437 & n5438 ) | ( n5437 & ~n5439 ) | ( n5438 & ~n5439 ) ;
  assign n5441 = ( n5238 & n5427 ) | ( n5238 & n5440 ) | ( n5427 & n5440 ) ;
  assign n5442 = ( ~n5238 & n5427 ) | ( ~n5238 & n5440 ) | ( n5427 & n5440 ) ;
  assign n5443 = ( n5238 & ~n5441 ) | ( n5238 & n5442 ) | ( ~n5441 & n5442 ) ;
  assign n5444 = n372 & n4020 ;
  assign n5445 = x41 & n5444 ;
  assign n5446 = x72 & n4027 ;
  assign n5447 = x71 & n4024 ;
  assign n5448 = n5446 | n5447 ;
  assign n5449 = x70 & n4223 ;
  assign n5450 = n5448 | n5449 ;
  assign n5451 = ( ~x41 & n5444 ) | ( ~x41 & n5450 ) | ( n5444 & n5450 ) ;
  assign n5452 = x41 & ~n5450 ;
  assign n5453 = ( ~n5445 & n5451 ) | ( ~n5445 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5454 = ( ~n5250 & n5443 ) | ( ~n5250 & n5453 ) | ( n5443 & n5453 ) ;
  assign n5455 = ( n5250 & n5443 ) | ( n5250 & n5453 ) | ( n5443 & n5453 ) ;
  assign n5456 = ( n5250 & n5454 ) | ( n5250 & ~n5455 ) | ( n5454 & ~n5455 ) ;
  assign n5457 = ( n5264 & n5417 ) | ( n5264 & n5456 ) | ( n5417 & n5456 ) ;
  assign n5458 = ( ~n5264 & n5417 ) | ( ~n5264 & n5456 ) | ( n5417 & n5456 ) ;
  assign n5459 = ( n5264 & ~n5457 ) | ( n5264 & n5458 ) | ( ~n5457 & n5458 ) ;
  assign n5460 = n697 & n2982 ;
  assign n5461 = x35 & n5460 ;
  assign n5462 = x78 & n2989 ;
  assign n5463 = x77 & n2986 ;
  assign n5464 = n5462 | n5463 ;
  assign n5465 = x76 & n3159 ;
  assign n5466 = n5464 | n5465 ;
  assign n5467 = ( ~x35 & n5460 ) | ( ~x35 & n5466 ) | ( n5460 & n5466 ) ;
  assign n5468 = x35 & ~n5466 ;
  assign n5469 = ( ~n5461 & n5467 ) | ( ~n5461 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5470 = ( n5266 & ~n5459 ) | ( n5266 & n5469 ) | ( ~n5459 & n5469 ) ;
  assign n5471 = ( n5266 & n5459 ) | ( n5266 & n5469 ) | ( n5459 & n5469 ) ;
  assign n5472 = ( n5459 & n5470 ) | ( n5459 & ~n5471 ) | ( n5470 & ~n5471 ) ;
  assign n5473 = ( n5280 & n5407 ) | ( n5280 & n5472 ) | ( n5407 & n5472 ) ;
  assign n5474 = ( ~n5280 & n5407 ) | ( ~n5280 & n5472 ) | ( n5407 & n5472 ) ;
  assign n5475 = ( n5280 & ~n5473 ) | ( n5280 & n5474 ) | ( ~n5473 & n5474 ) ;
  assign n5476 = n1190 & n2137 ;
  assign n5477 = x29 & n5476 ;
  assign n5478 = x84 & n2144 ;
  assign n5479 = x83 & n2141 ;
  assign n5480 = n5478 | n5479 ;
  assign n5481 = x82 & n2267 ;
  assign n5482 = n5480 | n5481 ;
  assign n5483 = ( ~x29 & n5476 ) | ( ~x29 & n5482 ) | ( n5476 & n5482 ) ;
  assign n5484 = x29 & ~n5482 ;
  assign n5485 = ( ~n5477 & n5483 ) | ( ~n5477 & n5484 ) | ( n5483 & n5484 ) ;
  assign n5486 = ( n5282 & ~n5475 ) | ( n5282 & n5485 ) | ( ~n5475 & n5485 ) ;
  assign n5487 = ( n5282 & n5475 ) | ( n5282 & n5485 ) | ( n5475 & n5485 ) ;
  assign n5488 = ( n5475 & n5486 ) | ( n5475 & ~n5487 ) | ( n5486 & ~n5487 ) ;
  assign n5489 = ( n5296 & n5397 ) | ( n5296 & n5488 ) | ( n5397 & n5488 ) ;
  assign n5490 = ( ~n5296 & n5397 ) | ( ~n5296 & n5488 ) | ( n5397 & n5488 ) ;
  assign n5491 = ( n5296 & ~n5489 ) | ( n5296 & n5490 ) | ( ~n5489 & n5490 ) ;
  assign n5492 = ( n5298 & n5387 ) | ( n5298 & n5491 ) | ( n5387 & n5491 ) ;
  assign n5493 = ( ~n5298 & n5387 ) | ( ~n5298 & n5491 ) | ( n5387 & n5491 ) ;
  assign n5494 = ( n5298 & ~n5492 ) | ( n5298 & n5493 ) | ( ~n5492 & n5493 ) ;
  assign n5495 = n1146 & n2220 ;
  assign n5496 = x20 & n5495 ;
  assign n5497 = x93 & n1153 ;
  assign n5498 = x92 & n1150 ;
  assign n5499 = n5497 | n5498 ;
  assign n5500 = x91 & n1217 ;
  assign n5501 = n5499 | n5500 ;
  assign n5502 = ( ~x20 & n5495 ) | ( ~x20 & n5501 ) | ( n5495 & n5501 ) ;
  assign n5503 = x20 & ~n5501 ;
  assign n5504 = ( ~n5496 & n5502 ) | ( ~n5496 & n5503 ) | ( n5502 & n5503 ) ;
  assign n5505 = ( n5312 & n5494 ) | ( n5312 & n5504 ) | ( n5494 & n5504 ) ;
  assign n5506 = ( ~n5312 & n5494 ) | ( ~n5312 & n5504 ) | ( n5494 & n5504 ) ;
  assign n5507 = ( n5312 & ~n5505 ) | ( n5312 & n5506 ) | ( ~n5505 & n5506 ) ;
  assign n5508 = n874 & n2772 ;
  assign n5509 = x17 & n5508 ;
  assign n5510 = x96 & n881 ;
  assign n5511 = x95 & n878 ;
  assign n5512 = n5510 | n5511 ;
  assign n5513 = x94 & n959 ;
  assign n5514 = n5512 | n5513 ;
  assign n5515 = ( ~x17 & n5508 ) | ( ~x17 & n5514 ) | ( n5508 & n5514 ) ;
  assign n5516 = x17 & ~n5514 ;
  assign n5517 = ( ~n5509 & n5515 ) | ( ~n5509 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5518 = ( n5314 & ~n5507 ) | ( n5314 & n5517 ) | ( ~n5507 & n5517 ) ;
  assign n5519 = ( n5314 & n5507 ) | ( n5314 & n5517 ) | ( n5507 & n5517 ) ;
  assign n5520 = ( n5507 & n5518 ) | ( n5507 & ~n5519 ) | ( n5518 & ~n5519 ) ;
  assign n5521 = ( n5317 & n5377 ) | ( n5317 & n5520 ) | ( n5377 & n5520 ) ;
  assign n5522 = ( ~n5317 & n5377 ) | ( ~n5317 & n5520 ) | ( n5377 & n5520 ) ;
  assign n5523 = ( n5317 & ~n5521 ) | ( n5317 & n5522 ) | ( ~n5521 & n5522 ) ;
  assign n5524 = n449 & n3764 ;
  assign n5525 = x11 & n5524 ;
  assign n5526 = x101 & n453 ;
  assign n5527 = x100 & n536 ;
  assign n5528 = n5526 | n5527 ;
  assign n5529 = x102 & n456 ;
  assign n5530 = n5528 | n5529 ;
  assign n5531 = ( ~x11 & n5524 ) | ( ~x11 & n5530 ) | ( n5524 & n5530 ) ;
  assign n5532 = x11 & ~n5530 ;
  assign n5533 = ( ~n5525 & n5531 ) | ( ~n5525 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5534 = ( n5321 & ~n5523 ) | ( n5321 & n5533 ) | ( ~n5523 & n5533 ) ;
  assign n5535 = ( n5321 & n5523 ) | ( n5321 & n5533 ) | ( n5523 & n5533 ) ;
  assign n5536 = ( n5523 & n5534 ) | ( n5523 & ~n5535 ) | ( n5534 & ~n5535 ) ;
  assign n5537 = ( n5323 & n5367 ) | ( n5323 & n5536 ) | ( n5367 & n5536 ) ;
  assign n5538 = ( ~n5323 & n5367 ) | ( ~n5323 & n5536 ) | ( n5367 & n5536 ) ;
  assign n5539 = ( n5323 & ~n5537 ) | ( n5323 & n5538 ) | ( ~n5537 & n5538 ) ;
  assign n5540 = n206 & n4914 ;
  assign n5541 = x5 & n5540 ;
  assign n5542 = x108 & n205 ;
  assign n5543 = x107 & n201 ;
  assign n5544 = n5542 | n5543 ;
  assign n5545 = x106 & n221 ;
  assign n5546 = n5544 | n5545 ;
  assign n5547 = ( ~x5 & n5540 ) | ( ~x5 & n5546 ) | ( n5540 & n5546 ) ;
  assign n5548 = x5 & ~n5546 ;
  assign n5549 = ( ~n5541 & n5547 ) | ( ~n5541 & n5548 ) | ( n5547 & n5548 ) ;
  assign n5550 = ( n5326 & ~n5539 ) | ( n5326 & n5549 ) | ( ~n5539 & n5549 ) ;
  assign n5551 = ( n5326 & n5539 ) | ( n5326 & n5549 ) | ( n5539 & n5549 ) ;
  assign n5552 = ( n5539 & n5550 ) | ( n5539 & ~n5551 ) | ( n5550 & ~n5551 ) ;
  assign n5553 = ( n5343 & n5357 ) | ( n5343 & n5552 ) | ( n5357 & n5552 ) ;
  assign n5554 = ( ~n5343 & n5357 ) | ( ~n5343 & n5552 ) | ( n5357 & n5552 ) ;
  assign n5555 = ( n5343 & ~n5553 ) | ( n5343 & n5554 ) | ( ~n5553 & n5554 ) ;
  assign n5556 = ( ~x111 & x112 ) | ( ~x111 & n5346 ) | ( x112 & n5346 ) ;
  assign n5557 = ( x111 & x112 ) | ( x111 & n5346 ) | ( x112 & n5346 ) ;
  assign n5558 = ( x111 & n5556 ) | ( x111 & ~n5557 ) | ( n5556 & ~n5557 ) ;
  assign n5559 = x0 & n5558 ;
  assign n5560 = ( x1 & x2 ) | ( x1 & n5559 ) | ( x2 & n5559 ) ;
  assign n5561 = x111 & n172 ;
  assign n5562 = x112 | n5561 ;
  assign n5563 = ( n147 & n5561 ) | ( n147 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = ( ~x110 & n135 ) | ( ~x110 & n174 ) | ( n135 & n174 ) ;
  assign n5565 = n5563 | n5564 ;
  assign n5566 = n5560 | n5565 ;
  assign n5567 = n5560 & n5565 ;
  assign n5568 = n5566 & ~n5567 ;
  assign n5569 = n301 & n4331 ;
  assign n5570 = x8 & n5569 ;
  assign n5571 = x106 & n309 ;
  assign n5572 = x105 & n306 ;
  assign n5573 = n5571 | n5572 ;
  assign n5574 = x104 & n359 ;
  assign n5575 = n5573 | n5574 ;
  assign n5576 = ( ~x8 & n5569 ) | ( ~x8 & n5575 ) | ( n5569 & n5575 ) ;
  assign n5577 = x8 & ~n5575 ;
  assign n5578 = ( ~n5570 & n5576 ) | ( ~n5570 & n5577 ) | ( n5576 & n5577 ) ;
  assign n5579 = n449 & n3941 ;
  assign n5580 = x11 & n5579 ;
  assign n5581 = x103 & n456 ;
  assign n5582 = x102 & n453 ;
  assign n5583 = n5581 | n5582 ;
  assign n5584 = x101 & n536 ;
  assign n5585 = n5583 | n5584 ;
  assign n5586 = ( ~x11 & n5579 ) | ( ~x11 & n5585 ) | ( n5579 & n5585 ) ;
  assign n5587 = x11 & ~n5585 ;
  assign n5588 = ( ~n5580 & n5586 ) | ( ~n5580 & n5587 ) | ( n5586 & n5587 ) ;
  assign n5589 = n649 & n3264 ;
  assign n5590 = x14 & n5589 ;
  assign n5591 = x100 & n656 ;
  assign n5592 = x99 & n653 ;
  assign n5593 = n5591 | n5592 ;
  assign n5594 = x98 & n744 ;
  assign n5595 = n5593 | n5594 ;
  assign n5596 = ( ~x14 & n5589 ) | ( ~x14 & n5595 ) | ( n5589 & n5595 ) ;
  assign n5597 = x14 & ~n5595 ;
  assign n5598 = ( ~n5590 & n5596 ) | ( ~n5590 & n5597 ) | ( n5596 & n5597 ) ;
  assign n5599 = n1146 & n2476 ;
  assign n5600 = x20 & n5599 ;
  assign n5601 = x94 & n1153 ;
  assign n5602 = x93 & n1150 ;
  assign n5603 = n5601 | n5602 ;
  assign n5604 = x92 & n1217 ;
  assign n5605 = n5603 | n5604 ;
  assign n5606 = ( ~x20 & n5599 ) | ( ~x20 & n5605 ) | ( n5599 & n5605 ) ;
  assign n5607 = x20 & ~n5605 ;
  assign n5608 = ( ~n5600 & n5606 ) | ( ~n5600 & n5607 ) | ( n5606 & n5607 ) ;
  assign n5609 = n1602 & n1755 ;
  assign n5610 = x26 & n5609 ;
  assign n5611 = x88 & n1762 ;
  assign n5612 = x87 & n1759 ;
  assign n5613 = n5611 | n5612 ;
  assign n5614 = x86 & n1895 ;
  assign n5615 = n5613 | n5614 ;
  assign n5616 = ( ~x26 & n5609 ) | ( ~x26 & n5615 ) | ( n5609 & n5615 ) ;
  assign n5617 = x26 & ~n5615 ;
  assign n5618 = ( ~n5610 & n5616 ) | ( ~n5610 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5619 = n1368 & n2137 ;
  assign n5620 = x29 & n5619 ;
  assign n5621 = x85 & n2144 ;
  assign n5622 = x84 & n2141 ;
  assign n5623 = n5621 | n5622 ;
  assign n5624 = x83 & n2267 ;
  assign n5625 = n5623 | n5624 ;
  assign n5626 = ( ~x29 & n5619 ) | ( ~x29 & n5625 ) | ( n5619 & n5625 ) ;
  assign n5627 = x29 & ~n5625 ;
  assign n5628 = ( ~n5620 & n5626 ) | ( ~n5620 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5629 = n276 & n4625 ;
  assign n5630 = x44 & n5629 ;
  assign n5631 = x70 & n4791 ;
  assign n5632 = x69 & n4621 ;
  assign n5633 = n5631 | n5632 ;
  assign n5634 = x68 & n4795 ;
  assign n5635 = n5633 | n5634 ;
  assign n5636 = ( ~x44 & n5629 ) | ( ~x44 & n5635 ) | ( n5629 & n5635 ) ;
  assign n5637 = x44 & ~n5635 ;
  assign n5638 = ( ~n5630 & n5636 ) | ( ~n5630 & n5637 ) | ( n5636 & n5637 ) ;
  assign n5639 = n5233 | n5436 ;
  assign n5640 = x47 & n5639 ;
  assign n5641 = x67 & n5230 ;
  assign n5642 = x66 & n5227 ;
  assign n5643 = n5641 | n5642 ;
  assign n5644 = x65 & n5434 ;
  assign n5645 = n5643 | n5644 ;
  assign n5646 = n169 & n5223 ;
  assign n5647 = n5645 | n5646 ;
  assign n5648 = x47 & x48 ;
  assign n5649 = x47 | x48 ;
  assign n5650 = ~n5648 & n5649 ;
  assign n5651 = x64 & n5650 ;
  assign n5652 = ( n5640 & ~n5647 ) | ( n5640 & n5651 ) | ( ~n5647 & n5651 ) ;
  assign n5653 = x47 & ~n5647 ;
  assign n5654 = ( ~n5640 & n5647 ) | ( ~n5640 & n5653 ) | ( n5647 & n5653 ) ;
  assign n5655 = ( n5651 & n5653 ) | ( n5651 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5656 = ( n5652 & n5654 ) | ( n5652 & ~n5655 ) | ( n5654 & ~n5655 ) ;
  assign n5657 = ( n5441 & n5638 ) | ( n5441 & n5656 ) | ( n5638 & n5656 ) ;
  assign n5658 = ( ~n5441 & n5638 ) | ( ~n5441 & n5656 ) | ( n5638 & n5656 ) ;
  assign n5659 = ( n5441 & ~n5657 ) | ( n5441 & n5658 ) | ( ~n5657 & n5658 ) ;
  assign n5660 = n388 & n4020 ;
  assign n5661 = x41 & n5660 ;
  assign n5662 = x73 & n4027 ;
  assign n5663 = x72 & n4024 ;
  assign n5664 = n5662 | n5663 ;
  assign n5665 = x71 & n4223 ;
  assign n5666 = n5664 | n5665 ;
  assign n5667 = ( ~x41 & n5660 ) | ( ~x41 & n5666 ) | ( n5660 & n5666 ) ;
  assign n5668 = x41 & ~n5666 ;
  assign n5669 = ( ~n5661 & n5667 ) | ( ~n5661 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5670 = ( n5455 & n5659 ) | ( n5455 & n5669 ) | ( n5659 & n5669 ) ;
  assign n5671 = ( n5455 & ~n5659 ) | ( n5455 & n5669 ) | ( ~n5659 & n5669 ) ;
  assign n5672 = ( n5659 & ~n5670 ) | ( n5659 & n5671 ) | ( ~n5670 & n5671 ) ;
  assign n5673 = n565 & n3492 ;
  assign n5674 = x38 & n5673 ;
  assign n5675 = x76 & n3499 ;
  assign n5676 = x75 & n3496 ;
  assign n5677 = n5675 | n5676 ;
  assign n5678 = x74 & n3662 ;
  assign n5679 = n5677 | n5678 ;
  assign n5680 = ( ~x38 & n5673 ) | ( ~x38 & n5679 ) | ( n5673 & n5679 ) ;
  assign n5681 = x38 & ~n5679 ;
  assign n5682 = ( ~n5674 & n5680 ) | ( ~n5674 & n5681 ) | ( n5680 & n5681 ) ;
  assign n5683 = ( n5457 & ~n5672 ) | ( n5457 & n5682 ) | ( ~n5672 & n5682 ) ;
  assign n5684 = ( n5457 & n5672 ) | ( n5457 & n5682 ) | ( n5672 & n5682 ) ;
  assign n5685 = ( n5672 & n5683 ) | ( n5672 & ~n5684 ) | ( n5683 & ~n5684 ) ;
  assign n5686 = n823 & n2982 ;
  assign n5687 = x35 & n5686 ;
  assign n5688 = x79 & n2989 ;
  assign n5689 = x78 & n2986 ;
  assign n5690 = n5688 | n5689 ;
  assign n5691 = x77 & n3159 ;
  assign n5692 = n5690 | n5691 ;
  assign n5693 = ( ~x35 & n5686 ) | ( ~x35 & n5692 ) | ( n5686 & n5692 ) ;
  assign n5694 = x35 & ~n5692 ;
  assign n5695 = ( ~n5687 & n5693 ) | ( ~n5687 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5696 = ( n5471 & n5685 ) | ( n5471 & n5695 ) | ( n5685 & n5695 ) ;
  assign n5697 = ( ~n5471 & n5685 ) | ( ~n5471 & n5695 ) | ( n5685 & n5695 ) ;
  assign n5698 = ( n5471 & ~n5696 ) | ( n5471 & n5697 ) | ( ~n5696 & n5697 ) ;
  assign n5699 = n1006 & n2545 ;
  assign n5700 = x32 & n5699 ;
  assign n5701 = x82 & n2552 ;
  assign n5702 = x81 & n2549 ;
  assign n5703 = n5701 | n5702 ;
  assign n5704 = x80 & n2696 ;
  assign n5705 = n5703 | n5704 ;
  assign n5706 = ( ~x32 & n5699 ) | ( ~x32 & n5705 ) | ( n5699 & n5705 ) ;
  assign n5707 = x32 & ~n5705 ;
  assign n5708 = ( ~n5700 & n5706 ) | ( ~n5700 & n5707 ) | ( n5706 & n5707 ) ;
  assign n5709 = ( n5473 & ~n5698 ) | ( n5473 & n5708 ) | ( ~n5698 & n5708 ) ;
  assign n5710 = ( n5473 & n5698 ) | ( n5473 & n5708 ) | ( n5698 & n5708 ) ;
  assign n5711 = ( n5698 & n5709 ) | ( n5698 & ~n5710 ) | ( n5709 & ~n5710 ) ;
  assign n5712 = ( n5487 & n5628 ) | ( n5487 & n5711 ) | ( n5628 & n5711 ) ;
  assign n5713 = ( ~n5487 & n5628 ) | ( ~n5487 & n5711 ) | ( n5628 & n5711 ) ;
  assign n5714 = ( n5487 & ~n5712 ) | ( n5487 & n5713 ) | ( ~n5712 & n5713 ) ;
  assign n5715 = ( n5489 & n5618 ) | ( n5489 & n5714 ) | ( n5618 & n5714 ) ;
  assign n5716 = ( ~n5489 & n5618 ) | ( ~n5489 & n5714 ) | ( n5618 & n5714 ) ;
  assign n5717 = ( n5489 & ~n5715 ) | ( n5489 & n5716 ) | ( ~n5715 & n5716 ) ;
  assign n5718 = n1427 & n1959 ;
  assign n5719 = x23 & n5718 ;
  assign n5720 = x91 & n1434 ;
  assign n5721 = x90 & n1431 ;
  assign n5722 = n5720 | n5721 ;
  assign n5723 = x89 & n1531 ;
  assign n5724 = n5722 | n5723 ;
  assign n5725 = ( ~x23 & n5718 ) | ( ~x23 & n5724 ) | ( n5718 & n5724 ) ;
  assign n5726 = x23 & ~n5724 ;
  assign n5727 = ( ~n5719 & n5725 ) | ( ~n5719 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = ( n5492 & ~n5717 ) | ( n5492 & n5727 ) | ( ~n5717 & n5727 ) ;
  assign n5729 = ( n5492 & n5717 ) | ( n5492 & n5727 ) | ( n5717 & n5727 ) ;
  assign n5730 = ( n5717 & n5728 ) | ( n5717 & ~n5729 ) | ( n5728 & ~n5729 ) ;
  assign n5731 = ( n5505 & n5608 ) | ( n5505 & n5730 ) | ( n5608 & n5730 ) ;
  assign n5732 = ( ~n5505 & n5608 ) | ( ~n5505 & n5730 ) | ( n5608 & n5730 ) ;
  assign n5733 = ( n5505 & ~n5731 ) | ( n5505 & n5732 ) | ( ~n5731 & n5732 ) ;
  assign n5734 = n874 & n2788 ;
  assign n5735 = x17 & n5734 ;
  assign n5736 = x97 & n881 ;
  assign n5737 = x96 & n878 ;
  assign n5738 = n5736 | n5737 ;
  assign n5739 = x95 & n959 ;
  assign n5740 = n5738 | n5739 ;
  assign n5741 = ( ~x17 & n5734 ) | ( ~x17 & n5740 ) | ( n5734 & n5740 ) ;
  assign n5742 = x17 & ~n5740 ;
  assign n5743 = ( ~n5735 & n5741 ) | ( ~n5735 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5744 = ( n5519 & ~n5733 ) | ( n5519 & n5743 ) | ( ~n5733 & n5743 ) ;
  assign n5745 = ( n5519 & n5733 ) | ( n5519 & n5743 ) | ( n5733 & n5743 ) ;
  assign n5746 = ( n5733 & n5744 ) | ( n5733 & ~n5745 ) | ( n5744 & ~n5745 ) ;
  assign n5747 = ( n5521 & n5598 ) | ( n5521 & n5746 ) | ( n5598 & n5746 ) ;
  assign n5748 = ( ~n5521 & n5598 ) | ( ~n5521 & n5746 ) | ( n5598 & n5746 ) ;
  assign n5749 = ( n5521 & ~n5747 ) | ( n5521 & n5748 ) | ( ~n5747 & n5748 ) ;
  assign n5750 = ( n5535 & ~n5588 ) | ( n5535 & n5749 ) | ( ~n5588 & n5749 ) ;
  assign n5751 = ( n5535 & n5588 ) | ( n5535 & n5749 ) | ( n5588 & n5749 ) ;
  assign n5752 = ( n5588 & n5750 ) | ( n5588 & ~n5751 ) | ( n5750 & ~n5751 ) ;
  assign n5753 = ( n5537 & n5578 ) | ( n5537 & n5752 ) | ( n5578 & n5752 ) ;
  assign n5754 = ( ~n5537 & n5578 ) | ( ~n5537 & n5752 ) | ( n5578 & n5752 ) ;
  assign n5755 = ( n5537 & ~n5753 ) | ( n5537 & n5754 ) | ( ~n5753 & n5754 ) ;
  assign n5756 = n206 & n4930 ;
  assign n5757 = x5 & n5756 ;
  assign n5758 = x109 & n205 ;
  assign n5759 = x108 & n201 ;
  assign n5760 = n5758 | n5759 ;
  assign n5761 = x107 & n221 ;
  assign n5762 = n5760 | n5761 ;
  assign n5763 = ( ~x5 & n5756 ) | ( ~x5 & n5762 ) | ( n5756 & n5762 ) ;
  assign n5764 = x5 & ~n5762 ;
  assign n5765 = ( ~n5757 & n5763 ) | ( ~n5757 & n5764 ) | ( n5763 & n5764 ) ;
  assign n5766 = ( n5551 & ~n5755 ) | ( n5551 & n5765 ) | ( ~n5755 & n5765 ) ;
  assign n5767 = ( n5551 & n5755 ) | ( n5551 & n5765 ) | ( n5755 & n5765 ) ;
  assign n5768 = ( n5755 & n5766 ) | ( n5755 & ~n5767 ) | ( n5766 & ~n5767 ) ;
  assign n5769 = ( n5553 & n5568 ) | ( n5553 & n5768 ) | ( n5568 & n5768 ) ;
  assign n5770 = ( ~n5553 & n5568 ) | ( ~n5553 & n5768 ) | ( n5568 & n5768 ) ;
  assign n5771 = ( n5553 & ~n5769 ) | ( n5553 & n5770 ) | ( ~n5769 & n5770 ) ;
  assign n5772 = ( ~x112 & x113 ) | ( ~x112 & n5557 ) | ( x113 & n5557 ) ;
  assign n5773 = ( x112 & x113 ) | ( x112 & n5557 ) | ( x113 & n5557 ) ;
  assign n5774 = ( x112 & n5772 ) | ( x112 & ~n5773 ) | ( n5772 & ~n5773 ) ;
  assign n5775 = x0 & n5774 ;
  assign n5776 = ( x1 & x2 ) | ( x1 & n5775 ) | ( x2 & n5775 ) ;
  assign n5777 = x112 & n172 ;
  assign n5778 = x113 | n5777 ;
  assign n5779 = ( n147 & n5777 ) | ( n147 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = ( ~x111 & n135 ) | ( ~x111 & n174 ) | ( n135 & n174 ) ;
  assign n5781 = n5779 | n5780 ;
  assign n5782 = n5776 | n5781 ;
  assign n5783 = n5776 & n5781 ;
  assign n5784 = n5782 & ~n5783 ;
  assign n5785 = n301 & n4523 ;
  assign n5786 = x8 & n5785 ;
  assign n5787 = x107 & n309 ;
  assign n5788 = x106 & n306 ;
  assign n5789 = n5787 | n5788 ;
  assign n5790 = x105 & n359 ;
  assign n5791 = n5789 | n5790 ;
  assign n5792 = ( ~x8 & n5785 ) | ( ~x8 & n5791 ) | ( n5785 & n5791 ) ;
  assign n5793 = x8 & ~n5791 ;
  assign n5794 = ( ~n5786 & n5792 ) | ( ~n5786 & n5793 ) | ( n5792 & n5793 ) ;
  assign n5795 = n649 & n3591 ;
  assign n5796 = x14 & n5795 ;
  assign n5797 = x101 & n656 ;
  assign n5798 = x100 & n653 ;
  assign n5799 = n5797 | n5798 ;
  assign n5800 = x99 & n744 ;
  assign n5801 = n5799 | n5800 ;
  assign n5802 = ( ~x14 & n5795 ) | ( ~x14 & n5801 ) | ( n5795 & n5801 ) ;
  assign n5803 = x14 & ~n5801 ;
  assign n5804 = ( ~n5796 & n5802 ) | ( ~n5796 & n5803 ) | ( n5802 & n5803 ) ;
  assign n5805 = n1146 & n2492 ;
  assign n5806 = x20 & n5805 ;
  assign n5807 = x95 & n1153 ;
  assign n5808 = x94 & n1150 ;
  assign n5809 = n5807 | n5808 ;
  assign n5810 = x93 & n1217 ;
  assign n5811 = n5809 | n5810 ;
  assign n5812 = ( ~x20 & n5805 ) | ( ~x20 & n5811 ) | ( n5805 & n5811 ) ;
  assign n5813 = x20 & ~n5811 ;
  assign n5814 = ( ~n5806 & n5812 ) | ( ~n5806 & n5813 ) | ( n5812 & n5813 ) ;
  assign n5815 = n1755 & n1822 ;
  assign n5816 = x26 & n5815 ;
  assign n5817 = x89 & n1762 ;
  assign n5818 = x88 & n1759 ;
  assign n5819 = n5817 | n5818 ;
  assign n5820 = x87 & n1895 ;
  assign n5821 = n5819 | n5820 ;
  assign n5822 = ( ~x26 & n5815 ) | ( ~x26 & n5821 ) | ( n5815 & n5821 ) ;
  assign n5823 = x26 & ~n5821 ;
  assign n5824 = ( ~n5816 & n5822 ) | ( ~n5816 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5825 = n1093 & n2545 ;
  assign n5826 = x32 & n5825 ;
  assign n5827 = x83 & n2552 ;
  assign n5828 = x82 & n2549 ;
  assign n5829 = n5827 | n5828 ;
  assign n5830 = x81 & n2696 ;
  assign n5831 = n5829 | n5830 ;
  assign n5832 = ( ~x32 & n5825 ) | ( ~x32 & n5831 ) | ( n5825 & n5831 ) ;
  assign n5833 = x32 & ~n5831 ;
  assign n5834 = ( ~n5826 & n5832 ) | ( ~n5826 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5835 = n626 & n3492 ;
  assign n5836 = x38 & n5835 ;
  assign n5837 = x77 & n3499 ;
  assign n5838 = x76 & n3496 ;
  assign n5839 = n5837 | n5838 ;
  assign n5840 = x75 & n3662 ;
  assign n5841 = n5839 | n5840 ;
  assign n5842 = ( ~x38 & n5835 ) | ( ~x38 & n5841 ) | ( n5835 & n5841 ) ;
  assign n5843 = x38 & ~n5841 ;
  assign n5844 = ( ~n5836 & n5842 ) | ( ~n5836 & n5843 ) | ( n5842 & n5843 ) ;
  assign n5845 = n193 & n5223 ;
  assign n5846 = x47 & n5845 ;
  assign n5847 = x68 & n5230 ;
  assign n5848 = x67 & n5227 ;
  assign n5849 = n5847 | n5848 ;
  assign n5850 = x66 & n5434 ;
  assign n5851 = n5849 | n5850 ;
  assign n5852 = ( ~x47 & n5845 ) | ( ~x47 & n5851 ) | ( n5845 & n5851 ) ;
  assign n5853 = x47 & ~n5851 ;
  assign n5854 = ( ~n5846 & n5852 ) | ( ~n5846 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5855 = x49 & x50 ;
  assign n5856 = x49 | x50 ;
  assign n5857 = ~n5855 & n5856 ;
  assign n5858 = n5650 & n5857 ;
  assign n5859 = n302 & n5858 ;
  assign n5860 = ~x47 & x49 ;
  assign n5861 = x48 & x49 ;
  assign n5862 = ( n5648 & n5860 ) | ( n5648 & ~n5861 ) | ( n5860 & ~n5861 ) ;
  assign n5863 = x64 & n5862 ;
  assign n5864 = n5859 | n5863 ;
  assign n5865 = ( n5650 & n5855 ) | ( n5650 & ~n5856 ) | ( n5855 & ~n5856 ) ;
  assign n5866 = x65 & n5865 ;
  assign n5867 = n5864 | n5866 ;
  assign n5868 = n5651 | n5867 ;
  assign n5869 = ( x50 & n5651 ) | ( x50 & ~n5867 ) | ( n5651 & ~n5867 ) ;
  assign n5870 = x50 & ~n5867 ;
  assign n5871 = ( n5868 & ~n5869 ) | ( n5868 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = ( ~n5655 & n5854 ) | ( ~n5655 & n5871 ) | ( n5854 & n5871 ) ;
  assign n5873 = ( n5655 & n5854 ) | ( n5655 & n5871 ) | ( n5854 & n5871 ) ;
  assign n5874 = ( n5655 & n5872 ) | ( n5655 & ~n5873 ) | ( n5872 & ~n5873 ) ;
  assign n5875 = n322 & n4625 ;
  assign n5876 = x44 & n5875 ;
  assign n5877 = x71 & n4791 ;
  assign n5878 = x70 & n4621 ;
  assign n5879 = n5877 | n5878 ;
  assign n5880 = x69 & n4795 ;
  assign n5881 = n5879 | n5880 ;
  assign n5882 = ( ~x44 & n5875 ) | ( ~x44 & n5881 ) | ( n5875 & n5881 ) ;
  assign n5883 = x44 & ~n5881 ;
  assign n5884 = ( ~n5876 & n5882 ) | ( ~n5876 & n5883 ) | ( n5882 & n5883 ) ;
  assign n5885 = ( n5657 & n5874 ) | ( n5657 & n5884 ) | ( n5874 & n5884 ) ;
  assign n5886 = ( ~n5657 & n5874 ) | ( ~n5657 & n5884 ) | ( n5874 & n5884 ) ;
  assign n5887 = ( n5657 & ~n5885 ) | ( n5657 & n5886 ) | ( ~n5885 & n5886 ) ;
  assign n5888 = n436 & n4020 ;
  assign n5889 = x41 & n5888 ;
  assign n5890 = x74 & n4027 ;
  assign n5891 = x73 & n4024 ;
  assign n5892 = n5890 | n5891 ;
  assign n5893 = x72 & n4223 ;
  assign n5894 = n5892 | n5893 ;
  assign n5895 = ( ~x41 & n5888 ) | ( ~x41 & n5894 ) | ( n5888 & n5894 ) ;
  assign n5896 = x41 & ~n5894 ;
  assign n5897 = ( ~n5889 & n5895 ) | ( ~n5889 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5898 = ( n5670 & ~n5887 ) | ( n5670 & n5897 ) | ( ~n5887 & n5897 ) ;
  assign n5899 = ( n5670 & n5887 ) | ( n5670 & n5897 ) | ( n5887 & n5897 ) ;
  assign n5900 = ( n5887 & n5898 ) | ( n5887 & ~n5899 ) | ( n5898 & ~n5899 ) ;
  assign n5901 = ( n5684 & n5844 ) | ( n5684 & n5900 ) | ( n5844 & n5900 ) ;
  assign n5902 = ( ~n5684 & n5844 ) | ( ~n5684 & n5900 ) | ( n5844 & n5900 ) ;
  assign n5903 = ( n5684 & ~n5901 ) | ( n5684 & n5902 ) | ( ~n5901 & n5902 ) ;
  assign n5904 = n840 & n2982 ;
  assign n5905 = x35 & n5904 ;
  assign n5906 = x80 & n2989 ;
  assign n5907 = x79 & n2986 ;
  assign n5908 = n5906 | n5907 ;
  assign n5909 = x78 & n3159 ;
  assign n5910 = n5908 | n5909 ;
  assign n5911 = ( ~x35 & n5904 ) | ( ~x35 & n5910 ) | ( n5904 & n5910 ) ;
  assign n5912 = x35 & ~n5910 ;
  assign n5913 = ( ~n5905 & n5911 ) | ( ~n5905 & n5912 ) | ( n5911 & n5912 ) ;
  assign n5914 = ( n5696 & ~n5903 ) | ( n5696 & n5913 ) | ( ~n5903 & n5913 ) ;
  assign n5915 = ( n5696 & n5903 ) | ( n5696 & n5913 ) | ( n5903 & n5913 ) ;
  assign n5916 = ( n5903 & n5914 ) | ( n5903 & ~n5915 ) | ( n5914 & ~n5915 ) ;
  assign n5917 = ( n5710 & n5834 ) | ( n5710 & n5916 ) | ( n5834 & n5916 ) ;
  assign n5918 = ( ~n5710 & n5834 ) | ( ~n5710 & n5916 ) | ( n5834 & n5916 ) ;
  assign n5919 = ( n5710 & ~n5917 ) | ( n5710 & n5918 ) | ( ~n5917 & n5918 ) ;
  assign n5920 = n1384 & n2137 ;
  assign n5921 = x29 & n5920 ;
  assign n5922 = x86 & n2144 ;
  assign n5923 = x85 & n2141 ;
  assign n5924 = n5922 | n5923 ;
  assign n5925 = x84 & n2267 ;
  assign n5926 = n5924 | n5925 ;
  assign n5927 = ( ~x29 & n5920 ) | ( ~x29 & n5926 ) | ( n5920 & n5926 ) ;
  assign n5928 = x29 & ~n5926 ;
  assign n5929 = ( ~n5921 & n5927 ) | ( ~n5921 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5930 = ( n5712 & ~n5919 ) | ( n5712 & n5929 ) | ( ~n5919 & n5929 ) ;
  assign n5931 = ( n5712 & n5919 ) | ( n5712 & n5929 ) | ( n5919 & n5929 ) ;
  assign n5932 = ( n5919 & n5930 ) | ( n5919 & ~n5931 ) | ( n5930 & ~n5931 ) ;
  assign n5933 = ( n5715 & n5824 ) | ( n5715 & n5932 ) | ( n5824 & n5932 ) ;
  assign n5934 = ( ~n5715 & n5824 ) | ( ~n5715 & n5932 ) | ( n5824 & n5932 ) ;
  assign n5935 = ( n5715 & ~n5933 ) | ( n5715 & n5934 ) | ( ~n5933 & n5934 ) ;
  assign n5936 = n1427 & n2083 ;
  assign n5937 = x23 & n5936 ;
  assign n5938 = x92 & n1434 ;
  assign n5939 = x91 & n1431 ;
  assign n5940 = n5938 | n5939 ;
  assign n5941 = x90 & n1531 ;
  assign n5942 = n5940 | n5941 ;
  assign n5943 = ( ~x23 & n5936 ) | ( ~x23 & n5942 ) | ( n5936 & n5942 ) ;
  assign n5944 = x23 & ~n5942 ;
  assign n5945 = ( ~n5937 & n5943 ) | ( ~n5937 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5946 = ( n5729 & ~n5935 ) | ( n5729 & n5945 ) | ( ~n5935 & n5945 ) ;
  assign n5947 = ( n5729 & n5935 ) | ( n5729 & n5945 ) | ( n5935 & n5945 ) ;
  assign n5948 = ( n5935 & n5946 ) | ( n5935 & ~n5947 ) | ( n5946 & ~n5947 ) ;
  assign n5949 = ( n5731 & n5814 ) | ( n5731 & n5948 ) | ( n5814 & n5948 ) ;
  assign n5950 = ( ~n5731 & n5814 ) | ( ~n5731 & n5948 ) | ( n5814 & n5948 ) ;
  assign n5951 = ( n5731 & ~n5949 ) | ( n5731 & n5950 ) | ( ~n5949 & n5950 ) ;
  assign n5952 = n874 & n2939 ;
  assign n5953 = x17 & n5952 ;
  assign n5954 = x98 & n881 ;
  assign n5955 = x97 & n878 ;
  assign n5956 = n5954 | n5955 ;
  assign n5957 = x96 & n959 ;
  assign n5958 = n5956 | n5957 ;
  assign n5959 = ( ~x17 & n5952 ) | ( ~x17 & n5958 ) | ( n5952 & n5958 ) ;
  assign n5960 = x17 & ~n5958 ;
  assign n5961 = ( ~n5953 & n5959 ) | ( ~n5953 & n5960 ) | ( n5959 & n5960 ) ;
  assign n5962 = ( n5745 & ~n5951 ) | ( n5745 & n5961 ) | ( ~n5951 & n5961 ) ;
  assign n5963 = ( n5745 & n5951 ) | ( n5745 & n5961 ) | ( n5951 & n5961 ) ;
  assign n5964 = ( n5951 & n5962 ) | ( n5951 & ~n5963 ) | ( n5962 & ~n5963 ) ;
  assign n5965 = ( n5747 & n5804 ) | ( n5747 & n5964 ) | ( n5804 & n5964 ) ;
  assign n5966 = ( ~n5747 & n5804 ) | ( ~n5747 & n5964 ) | ( n5804 & n5964 ) ;
  assign n5967 = ( n5747 & ~n5965 ) | ( n5747 & n5966 ) | ( ~n5965 & n5966 ) ;
  assign n5968 = n449 & n3957 ;
  assign n5969 = x11 & n5968 ;
  assign n5970 = x104 & n456 ;
  assign n5971 = x103 & n453 ;
  assign n5972 = n5970 | n5971 ;
  assign n5973 = x102 & n536 ;
  assign n5974 = n5972 | n5973 ;
  assign n5975 = ( ~x11 & n5968 ) | ( ~x11 & n5974 ) | ( n5968 & n5974 ) ;
  assign n5976 = x11 & ~n5974 ;
  assign n5977 = ( ~n5969 & n5975 ) | ( ~n5969 & n5976 ) | ( n5975 & n5976 ) ;
  assign n5978 = ( n5751 & ~n5967 ) | ( n5751 & n5977 ) | ( ~n5967 & n5977 ) ;
  assign n5979 = ( n5751 & n5967 ) | ( n5751 & n5977 ) | ( n5967 & n5977 ) ;
  assign n5980 = ( n5967 & n5978 ) | ( n5967 & ~n5979 ) | ( n5978 & ~n5979 ) ;
  assign n5981 = ( n5753 & n5794 ) | ( n5753 & n5980 ) | ( n5794 & n5980 ) ;
  assign n5982 = ( ~n5753 & n5794 ) | ( ~n5753 & n5980 ) | ( n5794 & n5980 ) ;
  assign n5983 = ( n5753 & ~n5981 ) | ( n5753 & n5982 ) | ( ~n5981 & n5982 ) ;
  assign n5984 = n206 & n5331 ;
  assign n5985 = x5 & n5984 ;
  assign n5986 = x110 & n205 ;
  assign n5987 = x109 & n201 ;
  assign n5988 = n5986 | n5987 ;
  assign n5989 = x108 & n221 ;
  assign n5990 = n5988 | n5989 ;
  assign n5991 = ( ~x5 & n5984 ) | ( ~x5 & n5990 ) | ( n5984 & n5990 ) ;
  assign n5992 = x5 & ~n5990 ;
  assign n5993 = ( ~n5985 & n5991 ) | ( ~n5985 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5994 = ( n5767 & ~n5983 ) | ( n5767 & n5993 ) | ( ~n5983 & n5993 ) ;
  assign n5995 = ( n5767 & n5983 ) | ( n5767 & n5993 ) | ( n5983 & n5993 ) ;
  assign n5996 = ( n5983 & n5994 ) | ( n5983 & ~n5995 ) | ( n5994 & ~n5995 ) ;
  assign n5997 = ( n5769 & n5784 ) | ( n5769 & n5996 ) | ( n5784 & n5996 ) ;
  assign n5998 = ( ~n5769 & n5784 ) | ( ~n5769 & n5996 ) | ( n5784 & n5996 ) ;
  assign n5999 = ( n5769 & ~n5997 ) | ( n5769 & n5998 ) | ( ~n5997 & n5998 ) ;
  assign n6000 = ( ~x113 & x114 ) | ( ~x113 & n5773 ) | ( x114 & n5773 ) ;
  assign n6001 = ( x113 & x114 ) | ( x113 & n5773 ) | ( x114 & n5773 ) ;
  assign n6002 = ( x113 & n6000 ) | ( x113 & ~n6001 ) | ( n6000 & ~n6001 ) ;
  assign n6003 = x0 & n6002 ;
  assign n6004 = ( x1 & x2 ) | ( x1 & n6003 ) | ( x2 & n6003 ) ;
  assign n6005 = x113 & n172 ;
  assign n6006 = ( ~x112 & n135 ) | ( ~x112 & n174 ) | ( n135 & n174 ) ;
  assign n6007 = n6005 | n6006 ;
  assign n6008 = x114 & n147 ;
  assign n6009 = n6007 | n6008 ;
  assign n6010 = n6004 | n6009 ;
  assign n6011 = n6004 & n6009 ;
  assign n6012 = n6010 & ~n6011 ;
  assign n6013 = n206 & n5347 ;
  assign n6014 = x5 & n6013 ;
  assign n6015 = x111 & n205 ;
  assign n6016 = x110 & n201 ;
  assign n6017 = n6015 | n6016 ;
  assign n6018 = x109 & n221 ;
  assign n6019 = n6017 | n6018 ;
  assign n6020 = ( ~x5 & n6013 ) | ( ~x5 & n6019 ) | ( n6013 & n6019 ) ;
  assign n6021 = x5 & ~n6019 ;
  assign n6022 = ( ~n6014 & n6020 ) | ( ~n6014 & n6021 ) | ( n6020 & n6021 ) ;
  assign n6023 = n449 & n4145 ;
  assign n6024 = x11 & n6023 ;
  assign n6025 = x105 & n456 ;
  assign n6026 = x104 & n453 ;
  assign n6027 = n6025 | n6026 ;
  assign n6028 = x103 & n536 ;
  assign n6029 = n6027 | n6028 ;
  assign n6030 = ( ~x11 & n6023 ) | ( ~x11 & n6029 ) | ( n6023 & n6029 ) ;
  assign n6031 = x11 & ~n6029 ;
  assign n6032 = ( ~n6024 & n6030 ) | ( ~n6024 & n6031 ) | ( n6030 & n6031 ) ;
  assign n6033 = n649 & n3764 ;
  assign n6034 = x14 & n6033 ;
  assign n6035 = x102 & n656 ;
  assign n6036 = x101 & n653 ;
  assign n6037 = n6035 | n6036 ;
  assign n6038 = x100 & n744 ;
  assign n6039 = n6037 | n6038 ;
  assign n6040 = ( ~x14 & n6033 ) | ( ~x14 & n6039 ) | ( n6033 & n6039 ) ;
  assign n6041 = x14 & ~n6039 ;
  assign n6042 = ( ~n6034 & n6040 ) | ( ~n6034 & n6041 ) | ( n6040 & n6041 ) ;
  assign n6043 = ~n6032 & n6042 ;
  assign n6044 = n6032 & ~n6042 ;
  assign n6045 = n6043 | n6044 ;
  assign n6046 = n1146 & n2772 ;
  assign n6047 = x20 & n6046 ;
  assign n6048 = x96 & n1153 ;
  assign n6049 = x95 & n1150 ;
  assign n6050 = n6048 | n6049 ;
  assign n6051 = x94 & n1217 ;
  assign n6052 = n6050 | n6051 ;
  assign n6053 = ( ~x20 & n6046 ) | ( ~x20 & n6052 ) | ( n6046 & n6052 ) ;
  assign n6054 = x20 & ~n6052 ;
  assign n6055 = ( ~n6047 & n6053 ) | ( ~n6047 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6056 = n1755 & n1838 ;
  assign n6057 = x26 & n6056 ;
  assign n6058 = x90 & n1762 ;
  assign n6059 = x89 & n1759 ;
  assign n6060 = n6058 | n6059 ;
  assign n6061 = x88 & n1895 ;
  assign n6062 = n6060 | n6061 ;
  assign n6063 = ( ~x26 & n6056 ) | ( ~x26 & n6062 ) | ( n6056 & n6062 ) ;
  assign n6064 = x26 & ~n6062 ;
  assign n6065 = ( ~n6057 & n6063 ) | ( ~n6057 & n6064 ) | ( n6063 & n6064 ) ;
  assign n6066 = n1190 & n2545 ;
  assign n6067 = x32 & n6066 ;
  assign n6068 = x84 & n2552 ;
  assign n6069 = x83 & n2549 ;
  assign n6070 = n6068 | n6069 ;
  assign n6071 = x82 & n2696 ;
  assign n6072 = n6070 | n6071 ;
  assign n6073 = ( ~x32 & n6066 ) | ( ~x32 & n6072 ) | ( n6066 & n6072 ) ;
  assign n6074 = x32 & ~n6072 ;
  assign n6075 = ( ~n6067 & n6073 ) | ( ~n6067 & n6074 ) | ( n6073 & n6074 ) ;
  assign n6076 = n508 & n4020 ;
  assign n6077 = x41 & n6076 ;
  assign n6078 = x75 & n4027 ;
  assign n6079 = x74 & n4024 ;
  assign n6080 = n6078 | n6079 ;
  assign n6081 = x73 & n4223 ;
  assign n6082 = n6080 | n6081 ;
  assign n6083 = ( ~x41 & n6076 ) | ( ~x41 & n6082 ) | ( n6076 & n6082 ) ;
  assign n6084 = x41 & ~n6082 ;
  assign n6085 = ( ~n6077 & n6083 ) | ( ~n6077 & n6084 ) | ( n6083 & n6084 ) ;
  assign n6086 = x66 & n5865 ;
  assign n6087 = x65 & n5862 ;
  assign n6088 = n6086 | n6087 ;
  assign n6089 = n226 & n5858 ;
  assign n6090 = n6088 | n6089 ;
  assign n6091 = ~n5650 & n5857 ;
  assign n6092 = ~n5862 & n6091 ;
  assign n6093 = x64 & n6092 ;
  assign n6094 = n6090 | n6093 ;
  assign n6095 = ~x50 & n6094 ;
  assign n6096 = ( x50 & n5868 ) | ( x50 & n6094 ) | ( n5868 & n6094 ) ;
  assign n6097 = n5868 & n6094 ;
  assign n6098 = ( n6095 & n6096 ) | ( n6095 & ~n6097 ) | ( n6096 & ~n6097 ) ;
  assign n6099 = n240 & n5223 ;
  assign n6100 = x47 & n6099 ;
  assign n6101 = x69 & n5230 ;
  assign n6102 = x68 & n5227 ;
  assign n6103 = n6101 | n6102 ;
  assign n6104 = x67 & n5434 ;
  assign n6105 = n6103 | n6104 ;
  assign n6106 = ( ~x47 & n6099 ) | ( ~x47 & n6105 ) | ( n6099 & n6105 ) ;
  assign n6107 = x47 & ~n6105 ;
  assign n6108 = ( ~n6100 & n6106 ) | ( ~n6100 & n6107 ) | ( n6106 & n6107 ) ;
  assign n6109 = ( n5873 & n6098 ) | ( n5873 & n6108 ) | ( n6098 & n6108 ) ;
  assign n6110 = ( ~n5873 & n6098 ) | ( ~n5873 & n6108 ) | ( n6098 & n6108 ) ;
  assign n6111 = ( n5873 & ~n6109 ) | ( n5873 & n6110 ) | ( ~n6109 & n6110 ) ;
  assign n6112 = n372 & n4625 ;
  assign n6113 = x44 & n6112 ;
  assign n6114 = x72 & n4791 ;
  assign n6115 = x71 & n4621 ;
  assign n6116 = n6114 | n6115 ;
  assign n6117 = x70 & n4795 ;
  assign n6118 = n6116 | n6117 ;
  assign n6119 = ( ~x44 & n6112 ) | ( ~x44 & n6118 ) | ( n6112 & n6118 ) ;
  assign n6120 = x44 & ~n6118 ;
  assign n6121 = ( ~n6113 & n6119 ) | ( ~n6113 & n6120 ) | ( n6119 & n6120 ) ;
  assign n6122 = ( n5885 & ~n6111 ) | ( n5885 & n6121 ) | ( ~n6111 & n6121 ) ;
  assign n6123 = ( n5885 & n6111 ) | ( n5885 & n6121 ) | ( n6111 & n6121 ) ;
  assign n6124 = ( n6111 & n6122 ) | ( n6111 & ~n6123 ) | ( n6122 & ~n6123 ) ;
  assign n6125 = ( n5899 & n6085 ) | ( n5899 & n6124 ) | ( n6085 & n6124 ) ;
  assign n6126 = ( ~n5899 & n6085 ) | ( ~n5899 & n6124 ) | ( n6085 & n6124 ) ;
  assign n6127 = ( n5899 & ~n6125 ) | ( n5899 & n6126 ) | ( ~n6125 & n6126 ) ;
  assign n6128 = n697 & n3492 ;
  assign n6129 = x38 & n6128 ;
  assign n6130 = x78 & n3499 ;
  assign n6131 = x77 & n3496 ;
  assign n6132 = n6130 | n6131 ;
  assign n6133 = x76 & n3662 ;
  assign n6134 = n6132 | n6133 ;
  assign n6135 = ( ~x38 & n6128 ) | ( ~x38 & n6134 ) | ( n6128 & n6134 ) ;
  assign n6136 = x38 & ~n6134 ;
  assign n6137 = ( ~n6129 & n6135 ) | ( ~n6129 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = ( ~n5901 & n6127 ) | ( ~n5901 & n6137 ) | ( n6127 & n6137 ) ;
  assign n6139 = ( n5901 & n6127 ) | ( n5901 & n6137 ) | ( n6127 & n6137 ) ;
  assign n6140 = ( n5901 & n6138 ) | ( n5901 & ~n6139 ) | ( n6138 & ~n6139 ) ;
  assign n6141 = n990 & n2982 ;
  assign n6142 = x35 & n6141 ;
  assign n6143 = x81 & n2989 ;
  assign n6144 = x80 & n2986 ;
  assign n6145 = n6143 | n6144 ;
  assign n6146 = x79 & n3159 ;
  assign n6147 = n6145 | n6146 ;
  assign n6148 = ( ~x35 & n6141 ) | ( ~x35 & n6147 ) | ( n6141 & n6147 ) ;
  assign n6149 = x35 & ~n6147 ;
  assign n6150 = ( ~n6142 & n6148 ) | ( ~n6142 & n6149 ) | ( n6148 & n6149 ) ;
  assign n6151 = ( n5915 & ~n6140 ) | ( n5915 & n6150 ) | ( ~n6140 & n6150 ) ;
  assign n6152 = ( n5915 & n6140 ) | ( n5915 & n6150 ) | ( n6140 & n6150 ) ;
  assign n6153 = ( n6140 & n6151 ) | ( n6140 & ~n6152 ) | ( n6151 & ~n6152 ) ;
  assign n6154 = ( n5917 & n6075 ) | ( n5917 & n6153 ) | ( n6075 & n6153 ) ;
  assign n6155 = ( ~n5917 & n6075 ) | ( ~n5917 & n6153 ) | ( n6075 & n6153 ) ;
  assign n6156 = ( n5917 & ~n6154 ) | ( n5917 & n6155 ) | ( ~n6154 & n6155 ) ;
  assign n6157 = n1494 & n2137 ;
  assign n6158 = x29 & n6157 ;
  assign n6159 = x87 & n2144 ;
  assign n6160 = x86 & n2141 ;
  assign n6161 = n6159 | n6160 ;
  assign n6162 = x85 & n2267 ;
  assign n6163 = n6161 | n6162 ;
  assign n6164 = ( ~x29 & n6157 ) | ( ~x29 & n6163 ) | ( n6157 & n6163 ) ;
  assign n6165 = x29 & ~n6163 ;
  assign n6166 = ( ~n6158 & n6164 ) | ( ~n6158 & n6165 ) | ( n6164 & n6165 ) ;
  assign n6167 = ( n5931 & ~n6156 ) | ( n5931 & n6166 ) | ( ~n6156 & n6166 ) ;
  assign n6168 = ( n5931 & n6156 ) | ( n5931 & n6166 ) | ( n6156 & n6166 ) ;
  assign n6169 = ( n6156 & n6167 ) | ( n6156 & ~n6168 ) | ( n6167 & ~n6168 ) ;
  assign n6170 = ( n5933 & n6065 ) | ( n5933 & n6169 ) | ( n6065 & n6169 ) ;
  assign n6171 = ( ~n5933 & n6065 ) | ( ~n5933 & n6169 ) | ( n6065 & n6169 ) ;
  assign n6172 = ( n5933 & ~n6170 ) | ( n5933 & n6171 ) | ( ~n6170 & n6171 ) ;
  assign n6173 = n1427 & n2220 ;
  assign n6174 = x23 & n6173 ;
  assign n6175 = x93 & n1434 ;
  assign n6176 = x92 & n1431 ;
  assign n6177 = n6175 | n6176 ;
  assign n6178 = x91 & n1531 ;
  assign n6179 = n6177 | n6178 ;
  assign n6180 = ( ~x23 & n6173 ) | ( ~x23 & n6179 ) | ( n6173 & n6179 ) ;
  assign n6181 = x23 & ~n6179 ;
  assign n6182 = ( ~n6174 & n6180 ) | ( ~n6174 & n6181 ) | ( n6180 & n6181 ) ;
  assign n6183 = ( n5947 & ~n6172 ) | ( n5947 & n6182 ) | ( ~n6172 & n6182 ) ;
  assign n6184 = ( n5947 & n6172 ) | ( n5947 & n6182 ) | ( n6172 & n6182 ) ;
  assign n6185 = ( n6172 & n6183 ) | ( n6172 & ~n6184 ) | ( n6183 & ~n6184 ) ;
  assign n6186 = ( n5949 & n6055 ) | ( n5949 & n6185 ) | ( n6055 & n6185 ) ;
  assign n6187 = ( ~n5949 & n6055 ) | ( ~n5949 & n6185 ) | ( n6055 & n6185 ) ;
  assign n6188 = ( n5949 & ~n6186 ) | ( n5949 & n6187 ) | ( ~n6186 & n6187 ) ;
  assign n6189 = n874 & n3248 ;
  assign n6190 = x17 & n6189 ;
  assign n6191 = x99 & n881 ;
  assign n6192 = x98 & n878 ;
  assign n6193 = n6191 | n6192 ;
  assign n6194 = x97 & n959 ;
  assign n6195 = n6193 | n6194 ;
  assign n6196 = ( ~x17 & n6189 ) | ( ~x17 & n6195 ) | ( n6189 & n6195 ) ;
  assign n6197 = x17 & ~n6195 ;
  assign n6198 = ( ~n6190 & n6196 ) | ( ~n6190 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = ( n5963 & ~n6188 ) | ( n5963 & n6198 ) | ( ~n6188 & n6198 ) ;
  assign n6200 = ( n5963 & n6188 ) | ( n5963 & n6198 ) | ( n6188 & n6198 ) ;
  assign n6201 = ( n6188 & n6199 ) | ( n6188 & ~n6200 ) | ( n6199 & ~n6200 ) ;
  assign n6202 = n5965 & n6201 ;
  assign n6203 = n5965 | n6201 ;
  assign n6204 = ~n6202 & n6203 ;
  assign n6205 = ( n5979 & n6045 ) | ( n5979 & n6204 ) | ( n6045 & n6204 ) ;
  assign n6206 = ( n5979 & ~n6045 ) | ( n5979 & n6204 ) | ( ~n6045 & n6204 ) ;
  assign n6207 = ( n6045 & ~n6205 ) | ( n6045 & n6206 ) | ( ~n6205 & n6206 ) ;
  assign n6208 = n301 & n4914 ;
  assign n6209 = x8 & n6208 ;
  assign n6210 = x108 & n309 ;
  assign n6211 = x107 & n306 ;
  assign n6212 = n6210 | n6211 ;
  assign n6213 = x106 & n359 ;
  assign n6214 = n6212 | n6213 ;
  assign n6215 = ( ~x8 & n6208 ) | ( ~x8 & n6214 ) | ( n6208 & n6214 ) ;
  assign n6216 = x8 & ~n6214 ;
  assign n6217 = ( ~n6209 & n6215 ) | ( ~n6209 & n6216 ) | ( n6215 & n6216 ) ;
  assign n6218 = ( n5981 & n6207 ) | ( n5981 & n6217 ) | ( n6207 & n6217 ) ;
  assign n6219 = ( ~n5981 & n6207 ) | ( ~n5981 & n6217 ) | ( n6207 & n6217 ) ;
  assign n6220 = ( n5981 & ~n6218 ) | ( n5981 & n6219 ) | ( ~n6218 & n6219 ) ;
  assign n6221 = ( n5995 & ~n6022 ) | ( n5995 & n6220 ) | ( ~n6022 & n6220 ) ;
  assign n6222 = ( n5995 & n6022 ) | ( n5995 & n6220 ) | ( n6022 & n6220 ) ;
  assign n6223 = ( n6022 & n6221 ) | ( n6022 & ~n6222 ) | ( n6221 & ~n6222 ) ;
  assign n6224 = ( n5997 & n6012 ) | ( n5997 & n6223 ) | ( n6012 & n6223 ) ;
  assign n6225 = ( ~n5997 & n6012 ) | ( ~n5997 & n6223 ) | ( n6012 & n6223 ) ;
  assign n6226 = ( n5997 & ~n6224 ) | ( n5997 & n6225 ) | ( ~n6224 & n6225 ) ;
  assign n6227 = n301 & n4930 ;
  assign n6228 = x8 & n6227 ;
  assign n6229 = x109 & n309 ;
  assign n6230 = x108 & n306 ;
  assign n6231 = n6229 | n6230 ;
  assign n6232 = x107 & n359 ;
  assign n6233 = n6231 | n6232 ;
  assign n6234 = ( ~x8 & n6227 ) | ( ~x8 & n6233 ) | ( n6227 & n6233 ) ;
  assign n6235 = x8 & ~n6233 ;
  assign n6236 = ( ~n6228 & n6234 ) | ( ~n6228 & n6235 ) | ( n6234 & n6235 ) ;
  assign n6237 = ( n5965 & n6042 ) | ( n5965 & n6201 ) | ( n6042 & n6201 ) ;
  assign n6238 = n649 & n3941 ;
  assign n6239 = x14 & n6238 ;
  assign n6240 = x103 & n656 ;
  assign n6241 = x102 & n653 ;
  assign n6242 = n6240 | n6241 ;
  assign n6243 = x101 & n744 ;
  assign n6244 = n6242 | n6243 ;
  assign n6245 = ( ~x14 & n6238 ) | ( ~x14 & n6244 ) | ( n6238 & n6244 ) ;
  assign n6246 = x14 & ~n6244 ;
  assign n6247 = ( ~n6239 & n6245 ) | ( ~n6239 & n6246 ) | ( n6245 & n6246 ) ;
  assign n6248 = n1602 & n2137 ;
  assign n6249 = x29 & n6248 ;
  assign n6250 = x88 & n2144 ;
  assign n6251 = x87 & n2141 ;
  assign n6252 = n6250 | n6251 ;
  assign n6253 = x86 & n2267 ;
  assign n6254 = n6252 | n6253 ;
  assign n6255 = ( ~x29 & n6248 ) | ( ~x29 & n6254 ) | ( n6248 & n6254 ) ;
  assign n6256 = x29 & ~n6254 ;
  assign n6257 = ( ~n6249 & n6255 ) | ( ~n6249 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6258 = n1368 & n2545 ;
  assign n6259 = x32 & n6258 ;
  assign n6260 = x85 & n2552 ;
  assign n6261 = x84 & n2549 ;
  assign n6262 = n6260 | n6261 ;
  assign n6263 = x83 & n2696 ;
  assign n6264 = n6262 | n6263 ;
  assign n6265 = ( ~x32 & n6258 ) | ( ~x32 & n6264 ) | ( n6258 & n6264 ) ;
  assign n6266 = x32 & ~n6264 ;
  assign n6267 = ( ~n6259 & n6265 ) | ( ~n6259 & n6266 ) | ( n6265 & n6266 ) ;
  assign n6268 = n823 & n3492 ;
  assign n6269 = x38 & n6268 ;
  assign n6270 = x79 & n3499 ;
  assign n6271 = x78 & n3496 ;
  assign n6272 = n6270 | n6271 ;
  assign n6273 = x77 & n3662 ;
  assign n6274 = n6272 | n6273 ;
  assign n6275 = ( ~x38 & n6268 ) | ( ~x38 & n6274 ) | ( n6268 & n6274 ) ;
  assign n6276 = x38 & ~n6274 ;
  assign n6277 = ( ~n6269 & n6275 ) | ( ~n6269 & n6276 ) | ( n6275 & n6276 ) ;
  assign n6278 = n565 & n4020 ;
  assign n6279 = x41 & n6278 ;
  assign n6280 = x76 & n4027 ;
  assign n6281 = x75 & n4024 ;
  assign n6282 = n6280 | n6281 ;
  assign n6283 = x74 & n4223 ;
  assign n6284 = n6282 | n6283 ;
  assign n6285 = ( ~x41 & n6278 ) | ( ~x41 & n6284 ) | ( n6278 & n6284 ) ;
  assign n6286 = x41 & ~n6284 ;
  assign n6287 = ( ~n6279 & n6285 ) | ( ~n6279 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = n276 & n5223 ;
  assign n6289 = x47 & n6288 ;
  assign n6290 = x70 & n5230 ;
  assign n6291 = x69 & n5227 ;
  assign n6292 = n6290 | n6291 ;
  assign n6293 = x68 & n5434 ;
  assign n6294 = n6292 | n6293 ;
  assign n6295 = ( ~x47 & n6288 ) | ( ~x47 & n6294 ) | ( n6288 & n6294 ) ;
  assign n6296 = x47 & ~n6294 ;
  assign n6297 = ( ~n6289 & n6295 ) | ( ~n6289 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6298 = n5868 | n6094 ;
  assign n6299 = x50 & n6298 ;
  assign n6300 = x67 & n5865 ;
  assign n6301 = x66 & n5862 ;
  assign n6302 = n6300 | n6301 ;
  assign n6303 = x65 & n6092 ;
  assign n6304 = n6302 | n6303 ;
  assign n6305 = n169 & n5858 ;
  assign n6306 = n6304 | n6305 ;
  assign n6307 = x50 & x51 ;
  assign n6308 = x50 | x51 ;
  assign n6309 = ~n6307 & n6308 ;
  assign n6310 = x64 & n6309 ;
  assign n6311 = ( n6299 & ~n6306 ) | ( n6299 & n6310 ) | ( ~n6306 & n6310 ) ;
  assign n6312 = x50 & ~n6306 ;
  assign n6313 = ( ~n6299 & n6306 ) | ( ~n6299 & n6312 ) | ( n6306 & n6312 ) ;
  assign n6314 = ( n6310 & n6312 ) | ( n6310 & n6313 ) | ( n6312 & n6313 ) ;
  assign n6315 = ( n6311 & n6313 ) | ( n6311 & ~n6314 ) | ( n6313 & ~n6314 ) ;
  assign n6316 = ( n6109 & n6297 ) | ( n6109 & n6315 ) | ( n6297 & n6315 ) ;
  assign n6317 = ( ~n6109 & n6297 ) | ( ~n6109 & n6315 ) | ( n6297 & n6315 ) ;
  assign n6318 = ( n6109 & ~n6316 ) | ( n6109 & n6317 ) | ( ~n6316 & n6317 ) ;
  assign n6319 = n388 & n4625 ;
  assign n6320 = x44 & n6319 ;
  assign n6321 = x73 & n4791 ;
  assign n6322 = x72 & n4621 ;
  assign n6323 = n6321 | n6322 ;
  assign n6324 = x71 & n4795 ;
  assign n6325 = n6323 | n6324 ;
  assign n6326 = ( ~x44 & n6319 ) | ( ~x44 & n6325 ) | ( n6319 & n6325 ) ;
  assign n6327 = x44 & ~n6325 ;
  assign n6328 = ( ~n6320 & n6326 ) | ( ~n6320 & n6327 ) | ( n6326 & n6327 ) ;
  assign n6329 = ( n6123 & ~n6318 ) | ( n6123 & n6328 ) | ( ~n6318 & n6328 ) ;
  assign n6330 = ( n6123 & n6318 ) | ( n6123 & n6328 ) | ( n6318 & n6328 ) ;
  assign n6331 = ( n6318 & n6329 ) | ( n6318 & ~n6330 ) | ( n6329 & ~n6330 ) ;
  assign n6332 = ( n6125 & n6287 ) | ( n6125 & n6331 ) | ( n6287 & n6331 ) ;
  assign n6333 = ( ~n6125 & n6287 ) | ( ~n6125 & n6331 ) | ( n6287 & n6331 ) ;
  assign n6334 = ( n6125 & ~n6332 ) | ( n6125 & n6333 ) | ( ~n6332 & n6333 ) ;
  assign n6335 = ( n6139 & n6277 ) | ( n6139 & n6334 ) | ( n6277 & n6334 ) ;
  assign n6336 = ( ~n6139 & n6277 ) | ( ~n6139 & n6334 ) | ( n6277 & n6334 ) ;
  assign n6337 = ( n6139 & ~n6335 ) | ( n6139 & n6336 ) | ( ~n6335 & n6336 ) ;
  assign n6338 = n1006 & n2982 ;
  assign n6339 = x35 & n6338 ;
  assign n6340 = x82 & n2989 ;
  assign n6341 = x81 & n2986 ;
  assign n6342 = n6340 | n6341 ;
  assign n6343 = x80 & n3159 ;
  assign n6344 = n6342 | n6343 ;
  assign n6345 = ( ~x35 & n6338 ) | ( ~x35 & n6344 ) | ( n6338 & n6344 ) ;
  assign n6346 = x35 & ~n6344 ;
  assign n6347 = ( ~n6339 & n6345 ) | ( ~n6339 & n6346 ) | ( n6345 & n6346 ) ;
  assign n6348 = ( n6152 & ~n6337 ) | ( n6152 & n6347 ) | ( ~n6337 & n6347 ) ;
  assign n6349 = ( n6152 & n6337 ) | ( n6152 & n6347 ) | ( n6337 & n6347 ) ;
  assign n6350 = ( n6337 & n6348 ) | ( n6337 & ~n6349 ) | ( n6348 & ~n6349 ) ;
  assign n6351 = ( n6154 & n6267 ) | ( n6154 & n6350 ) | ( n6267 & n6350 ) ;
  assign n6352 = ( ~n6154 & n6267 ) | ( ~n6154 & n6350 ) | ( n6267 & n6350 ) ;
  assign n6353 = ( n6154 & ~n6351 ) | ( n6154 & n6352 ) | ( ~n6351 & n6352 ) ;
  assign n6354 = ( n6168 & n6257 ) | ( n6168 & n6353 ) | ( n6257 & n6353 ) ;
  assign n6355 = ( ~n6168 & n6257 ) | ( ~n6168 & n6353 ) | ( n6257 & n6353 ) ;
  assign n6356 = ( n6168 & ~n6354 ) | ( n6168 & n6355 ) | ( ~n6354 & n6355 ) ;
  assign n6357 = n1755 & n1959 ;
  assign n6358 = x26 & n6357 ;
  assign n6359 = x91 & n1762 ;
  assign n6360 = x90 & n1759 ;
  assign n6361 = n6359 | n6360 ;
  assign n6362 = x89 & n1895 ;
  assign n6363 = n6361 | n6362 ;
  assign n6364 = ( ~x26 & n6357 ) | ( ~x26 & n6363 ) | ( n6357 & n6363 ) ;
  assign n6365 = x26 & ~n6363 ;
  assign n6366 = ( ~n6358 & n6364 ) | ( ~n6358 & n6365 ) | ( n6364 & n6365 ) ;
  assign n6367 = ( n6170 & n6356 ) | ( n6170 & n6366 ) | ( n6356 & n6366 ) ;
  assign n6368 = ( ~n6170 & n6356 ) | ( ~n6170 & n6366 ) | ( n6356 & n6366 ) ;
  assign n6369 = ( n6170 & ~n6367 ) | ( n6170 & n6368 ) | ( ~n6367 & n6368 ) ;
  assign n6370 = n1427 & n2476 ;
  assign n6371 = x23 & n6370 ;
  assign n6372 = x94 & n1434 ;
  assign n6373 = x93 & n1431 ;
  assign n6374 = n6372 | n6373 ;
  assign n6375 = x92 & n1531 ;
  assign n6376 = n6374 | n6375 ;
  assign n6377 = ( ~x23 & n6370 ) | ( ~x23 & n6376 ) | ( n6370 & n6376 ) ;
  assign n6378 = x23 & ~n6376 ;
  assign n6379 = ( ~n6371 & n6377 ) | ( ~n6371 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6380 = ( n6184 & n6369 ) | ( n6184 & n6379 ) | ( n6369 & n6379 ) ;
  assign n6381 = ( ~n6184 & n6369 ) | ( ~n6184 & n6379 ) | ( n6369 & n6379 ) ;
  assign n6382 = ( n6184 & ~n6380 ) | ( n6184 & n6381 ) | ( ~n6380 & n6381 ) ;
  assign n6383 = n1146 & n2788 ;
  assign n6384 = x20 & n6383 ;
  assign n6385 = x97 & n1153 ;
  assign n6386 = x96 & n1150 ;
  assign n6387 = n6385 | n6386 ;
  assign n6388 = x95 & n1217 ;
  assign n6389 = n6387 | n6388 ;
  assign n6390 = ( ~x20 & n6383 ) | ( ~x20 & n6389 ) | ( n6383 & n6389 ) ;
  assign n6391 = x20 & ~n6389 ;
  assign n6392 = ( ~n6384 & n6390 ) | ( ~n6384 & n6391 ) | ( n6390 & n6391 ) ;
  assign n6393 = ( n6186 & n6382 ) | ( n6186 & n6392 ) | ( n6382 & n6392 ) ;
  assign n6394 = ( ~n6186 & n6382 ) | ( ~n6186 & n6392 ) | ( n6382 & n6392 ) ;
  assign n6395 = ( n6186 & ~n6393 ) | ( n6186 & n6394 ) | ( ~n6393 & n6394 ) ;
  assign n6396 = n874 & n3264 ;
  assign n6397 = x17 & n6396 ;
  assign n6398 = x100 & n881 ;
  assign n6399 = x99 & n878 ;
  assign n6400 = n6398 | n6399 ;
  assign n6401 = x98 & n959 ;
  assign n6402 = n6400 | n6401 ;
  assign n6403 = ( ~x17 & n6396 ) | ( ~x17 & n6402 ) | ( n6396 & n6402 ) ;
  assign n6404 = x17 & ~n6402 ;
  assign n6405 = ( ~n6397 & n6403 ) | ( ~n6397 & n6404 ) | ( n6403 & n6404 ) ;
  assign n6406 = ( n6200 & ~n6395 ) | ( n6200 & n6405 ) | ( ~n6395 & n6405 ) ;
  assign n6407 = ( n6200 & n6395 ) | ( n6200 & n6405 ) | ( n6395 & n6405 ) ;
  assign n6408 = ( n6395 & n6406 ) | ( n6395 & ~n6407 ) | ( n6406 & ~n6407 ) ;
  assign n6409 = ( n6237 & n6247 ) | ( n6237 & n6408 ) | ( n6247 & n6408 ) ;
  assign n6410 = ( ~n6237 & n6247 ) | ( ~n6237 & n6408 ) | ( n6247 & n6408 ) ;
  assign n6411 = ( n6237 & ~n6409 ) | ( n6237 & n6410 ) | ( ~n6409 & n6410 ) ;
  assign n6412 = ( n5965 & ~n6042 ) | ( n5965 & n6201 ) | ( ~n6042 & n6201 ) ;
  assign n6413 = ( n6042 & ~n6237 ) | ( n6042 & n6412 ) | ( ~n6237 & n6412 ) ;
  assign n6414 = ( n5979 & n6032 ) | ( n5979 & n6413 ) | ( n6032 & n6413 ) ;
  assign n6415 = n449 & n4331 ;
  assign n6416 = x11 & n6415 ;
  assign n6417 = x106 & n456 ;
  assign n6418 = x105 & n453 ;
  assign n6419 = n6417 | n6418 ;
  assign n6420 = x104 & n536 ;
  assign n6421 = n6419 | n6420 ;
  assign n6422 = ( ~x11 & n6415 ) | ( ~x11 & n6421 ) | ( n6415 & n6421 ) ;
  assign n6423 = x11 & ~n6421 ;
  assign n6424 = ( ~n6416 & n6422 ) | ( ~n6416 & n6423 ) | ( n6422 & n6423 ) ;
  assign n6425 = ( ~n6411 & n6414 ) | ( ~n6411 & n6424 ) | ( n6414 & n6424 ) ;
  assign n6426 = ( n6411 & n6414 ) | ( n6411 & n6424 ) | ( n6414 & n6424 ) ;
  assign n6427 = ( n6411 & n6425 ) | ( n6411 & ~n6426 ) | ( n6425 & ~n6426 ) ;
  assign n6428 = ( n6218 & n6236 ) | ( n6218 & n6427 ) | ( n6236 & n6427 ) ;
  assign n6429 = ( ~n6218 & n6236 ) | ( ~n6218 & n6427 ) | ( n6236 & n6427 ) ;
  assign n6430 = ( n6218 & ~n6428 ) | ( n6218 & n6429 ) | ( ~n6428 & n6429 ) ;
  assign n6431 = n206 & n5558 ;
  assign n6432 = x5 & n6431 ;
  assign n6433 = x112 & n205 ;
  assign n6434 = x111 & n201 ;
  assign n6435 = n6433 | n6434 ;
  assign n6436 = x110 & n221 ;
  assign n6437 = n6435 | n6436 ;
  assign n6438 = ( ~x5 & n6431 ) | ( ~x5 & n6437 ) | ( n6431 & n6437 ) ;
  assign n6439 = x5 & ~n6437 ;
  assign n6440 = ( ~n6432 & n6438 ) | ( ~n6432 & n6439 ) | ( n6438 & n6439 ) ;
  assign n6441 = ( n6222 & n6430 ) | ( n6222 & n6440 ) | ( n6430 & n6440 ) ;
  assign n6442 = ( ~n6222 & n6430 ) | ( ~n6222 & n6440 ) | ( n6430 & n6440 ) ;
  assign n6443 = ( n6222 & ~n6441 ) | ( n6222 & n6442 ) | ( ~n6441 & n6442 ) ;
  assign n6444 = ( ~x114 & x115 ) | ( ~x114 & n6001 ) | ( x115 & n6001 ) ;
  assign n6445 = ( x114 & x115 ) | ( x114 & n6001 ) | ( x115 & n6001 ) ;
  assign n6446 = ( x114 & n6444 ) | ( x114 & ~n6445 ) | ( n6444 & ~n6445 ) ;
  assign n6447 = x0 & n6446 ;
  assign n6448 = ( x1 & x2 ) | ( x1 & n6447 ) | ( x2 & n6447 ) ;
  assign n6449 = x114 & n172 ;
  assign n6450 = ( ~x113 & n135 ) | ( ~x113 & n174 ) | ( n135 & n174 ) ;
  assign n6451 = n6449 | n6450 ;
  assign n6452 = x115 & n147 ;
  assign n6453 = n6451 | n6452 ;
  assign n6454 = n6448 | n6453 ;
  assign n6455 = n6448 & n6453 ;
  assign n6456 = n6454 & ~n6455 ;
  assign n6457 = ( n6224 & ~n6443 ) | ( n6224 & n6456 ) | ( ~n6443 & n6456 ) ;
  assign n6458 = ( n6224 & n6443 ) | ( n6224 & n6456 ) | ( n6443 & n6456 ) ;
  assign n6459 = ( n6443 & n6457 ) | ( n6443 & ~n6458 ) | ( n6457 & ~n6458 ) ;
  assign n6460 = ( ~x115 & x116 ) | ( ~x115 & n6445 ) | ( x116 & n6445 ) ;
  assign n6461 = ( x115 & x116 ) | ( x115 & n6445 ) | ( x116 & n6445 ) ;
  assign n6462 = ( x115 & n6460 ) | ( x115 & ~n6461 ) | ( n6460 & ~n6461 ) ;
  assign n6463 = x0 & n6462 ;
  assign n6464 = ( x1 & x2 ) | ( x1 & n6463 ) | ( x2 & n6463 ) ;
  assign n6465 = x115 & n172 ;
  assign n6466 = x116 | n6465 ;
  assign n6467 = ( n147 & n6465 ) | ( n147 & n6466 ) | ( n6465 & n6466 ) ;
  assign n6468 = ( ~x114 & n135 ) | ( ~x114 & n174 ) | ( n135 & n174 ) ;
  assign n6469 = n6467 | n6468 ;
  assign n6470 = n6464 | n6469 ;
  assign n6471 = n6464 & n6469 ;
  assign n6472 = n6470 & ~n6471 ;
  assign n6473 = n301 & n5331 ;
  assign n6474 = x8 & n6473 ;
  assign n6475 = x110 & n309 ;
  assign n6476 = x109 & n306 ;
  assign n6477 = n6475 | n6476 ;
  assign n6478 = x108 & n359 ;
  assign n6479 = n6477 | n6478 ;
  assign n6480 = ( ~x8 & n6473 ) | ( ~x8 & n6479 ) | ( n6473 & n6479 ) ;
  assign n6481 = x8 & ~n6479 ;
  assign n6482 = ( ~n6474 & n6480 ) | ( ~n6474 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6483 = n874 & n3591 ;
  assign n6484 = x17 & n6483 ;
  assign n6485 = x101 & n881 ;
  assign n6486 = x100 & n878 ;
  assign n6487 = n6485 | n6486 ;
  assign n6488 = x99 & n959 ;
  assign n6489 = n6487 | n6488 ;
  assign n6490 = ( ~x17 & n6483 ) | ( ~x17 & n6489 ) | ( n6483 & n6489 ) ;
  assign n6491 = x17 & ~n6489 ;
  assign n6492 = ( ~n6484 & n6490 ) | ( ~n6484 & n6491 ) | ( n6490 & n6491 ) ;
  assign n6493 = n1427 & n2492 ;
  assign n6494 = x23 & n6493 ;
  assign n6495 = x95 & n1434 ;
  assign n6496 = x94 & n1431 ;
  assign n6497 = n6495 | n6496 ;
  assign n6498 = x93 & n1531 ;
  assign n6499 = n6497 | n6498 ;
  assign n6500 = ( ~x23 & n6493 ) | ( ~x23 & n6499 ) | ( n6493 & n6499 ) ;
  assign n6501 = x23 & ~n6499 ;
  assign n6502 = ( ~n6494 & n6500 ) | ( ~n6494 & n6501 ) | ( n6500 & n6501 ) ;
  assign n6503 = n1822 & n2137 ;
  assign n6504 = x29 & n6503 ;
  assign n6505 = x89 & n2144 ;
  assign n6506 = x88 & n2141 ;
  assign n6507 = n6505 | n6506 ;
  assign n6508 = x87 & n2267 ;
  assign n6509 = n6507 | n6508 ;
  assign n6510 = ( ~x29 & n6503 ) | ( ~x29 & n6509 ) | ( n6503 & n6509 ) ;
  assign n6511 = x29 & ~n6509 ;
  assign n6512 = ( ~n6504 & n6510 ) | ( ~n6504 & n6511 ) | ( n6510 & n6511 ) ;
  assign n6513 = n1384 & n2545 ;
  assign n6514 = x32 & n6513 ;
  assign n6515 = x86 & n2552 ;
  assign n6516 = x85 & n2549 ;
  assign n6517 = n6515 | n6516 ;
  assign n6518 = x84 & n2696 ;
  assign n6519 = n6517 | n6518 ;
  assign n6520 = ( ~x32 & n6513 ) | ( ~x32 & n6519 ) | ( n6513 & n6519 ) ;
  assign n6521 = x32 & ~n6519 ;
  assign n6522 = ( ~n6514 & n6520 ) | ( ~n6514 & n6521 ) | ( n6520 & n6521 ) ;
  assign n6523 = n436 & n4625 ;
  assign n6524 = x44 & n6523 ;
  assign n6525 = x74 & n4791 ;
  assign n6526 = x73 & n4621 ;
  assign n6527 = n6525 | n6526 ;
  assign n6528 = x72 & n4795 ;
  assign n6529 = n6527 | n6528 ;
  assign n6530 = ( ~x44 & n6523 ) | ( ~x44 & n6529 ) | ( n6523 & n6529 ) ;
  assign n6531 = x44 & ~n6529 ;
  assign n6532 = ( ~n6524 & n6530 ) | ( ~n6524 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6533 = n193 & n5858 ;
  assign n6534 = x50 & n6533 ;
  assign n6535 = x68 & n5865 ;
  assign n6536 = x67 & n5862 ;
  assign n6537 = n6535 | n6536 ;
  assign n6538 = x66 & n6092 ;
  assign n6539 = n6537 | n6538 ;
  assign n6540 = ( ~x50 & n6533 ) | ( ~x50 & n6539 ) | ( n6533 & n6539 ) ;
  assign n6541 = x50 & ~n6539 ;
  assign n6542 = ( ~n6534 & n6540 ) | ( ~n6534 & n6541 ) | ( n6540 & n6541 ) ;
  assign n6543 = x52 & x53 ;
  assign n6544 = x52 | x53 ;
  assign n6545 = ~n6543 & n6544 ;
  assign n6546 = n6309 & n6545 ;
  assign n6547 = n302 & n6546 ;
  assign n6548 = ~x50 & x52 ;
  assign n6549 = x51 & x52 ;
  assign n6550 = ( n6307 & n6548 ) | ( n6307 & ~n6549 ) | ( n6548 & ~n6549 ) ;
  assign n6551 = x64 & n6550 ;
  assign n6552 = n6547 | n6551 ;
  assign n6553 = ( n6309 & n6543 ) | ( n6309 & ~n6544 ) | ( n6543 & ~n6544 ) ;
  assign n6554 = x65 & n6553 ;
  assign n6555 = n6552 | n6554 ;
  assign n6556 = n6310 | n6555 ;
  assign n6557 = ( x53 & n6310 ) | ( x53 & ~n6555 ) | ( n6310 & ~n6555 ) ;
  assign n6558 = x53 & ~n6555 ;
  assign n6559 = ( n6556 & ~n6557 ) | ( n6556 & n6558 ) | ( ~n6557 & n6558 ) ;
  assign n6560 = ( ~n6314 & n6542 ) | ( ~n6314 & n6559 ) | ( n6542 & n6559 ) ;
  assign n6561 = ( n6314 & n6542 ) | ( n6314 & n6559 ) | ( n6542 & n6559 ) ;
  assign n6562 = ( n6314 & n6560 ) | ( n6314 & ~n6561 ) | ( n6560 & ~n6561 ) ;
  assign n6563 = n322 & n5223 ;
  assign n6564 = x47 & n6563 ;
  assign n6565 = x71 & n5230 ;
  assign n6566 = x70 & n5227 ;
  assign n6567 = n6565 | n6566 ;
  assign n6568 = x69 & n5434 ;
  assign n6569 = n6567 | n6568 ;
  assign n6570 = ( ~x47 & n6563 ) | ( ~x47 & n6569 ) | ( n6563 & n6569 ) ;
  assign n6571 = x47 & ~n6569 ;
  assign n6572 = ( ~n6564 & n6570 ) | ( ~n6564 & n6571 ) | ( n6570 & n6571 ) ;
  assign n6573 = ( n6316 & ~n6562 ) | ( n6316 & n6572 ) | ( ~n6562 & n6572 ) ;
  assign n6574 = ( n6316 & n6562 ) | ( n6316 & n6572 ) | ( n6562 & n6572 ) ;
  assign n6575 = ( n6562 & n6573 ) | ( n6562 & ~n6574 ) | ( n6573 & ~n6574 ) ;
  assign n6576 = ( n6330 & n6532 ) | ( n6330 & n6575 ) | ( n6532 & n6575 ) ;
  assign n6577 = ( ~n6330 & n6532 ) | ( ~n6330 & n6575 ) | ( n6532 & n6575 ) ;
  assign n6578 = ( n6330 & ~n6576 ) | ( n6330 & n6577 ) | ( ~n6576 & n6577 ) ;
  assign n6579 = n626 & n4020 ;
  assign n6580 = x41 & n6579 ;
  assign n6581 = x77 & n4027 ;
  assign n6582 = x76 & n4024 ;
  assign n6583 = n6581 | n6582 ;
  assign n6584 = x75 & n4223 ;
  assign n6585 = n6583 | n6584 ;
  assign n6586 = ( ~x41 & n6579 ) | ( ~x41 & n6585 ) | ( n6579 & n6585 ) ;
  assign n6587 = x41 & ~n6585 ;
  assign n6588 = ( ~n6580 & n6586 ) | ( ~n6580 & n6587 ) | ( n6586 & n6587 ) ;
  assign n6589 = ( n6332 & n6578 ) | ( n6332 & n6588 ) | ( n6578 & n6588 ) ;
  assign n6590 = ( ~n6332 & n6578 ) | ( ~n6332 & n6588 ) | ( n6578 & n6588 ) ;
  assign n6591 = ( n6332 & ~n6589 ) | ( n6332 & n6590 ) | ( ~n6589 & n6590 ) ;
  assign n6592 = n840 & n3492 ;
  assign n6593 = x38 & n6592 ;
  assign n6594 = x80 & n3499 ;
  assign n6595 = x79 & n3496 ;
  assign n6596 = n6594 | n6595 ;
  assign n6597 = x78 & n3662 ;
  assign n6598 = n6596 | n6597 ;
  assign n6599 = ( ~x38 & n6592 ) | ( ~x38 & n6598 ) | ( n6592 & n6598 ) ;
  assign n6600 = x38 & ~n6598 ;
  assign n6601 = ( ~n6593 & n6599 ) | ( ~n6593 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6602 = ( n6335 & n6591 ) | ( n6335 & n6601 ) | ( n6591 & n6601 ) ;
  assign n6603 = ( ~n6335 & n6591 ) | ( ~n6335 & n6601 ) | ( n6591 & n6601 ) ;
  assign n6604 = ( n6335 & ~n6602 ) | ( n6335 & n6603 ) | ( ~n6602 & n6603 ) ;
  assign n6605 = n1093 & n2982 ;
  assign n6606 = x35 & n6605 ;
  assign n6607 = x83 & n2989 ;
  assign n6608 = x82 & n2986 ;
  assign n6609 = n6607 | n6608 ;
  assign n6610 = x81 & n3159 ;
  assign n6611 = n6609 | n6610 ;
  assign n6612 = ( ~x35 & n6605 ) | ( ~x35 & n6611 ) | ( n6605 & n6611 ) ;
  assign n6613 = x35 & ~n6611 ;
  assign n6614 = ( ~n6606 & n6612 ) | ( ~n6606 & n6613 ) | ( n6612 & n6613 ) ;
  assign n6615 = ( n6349 & ~n6604 ) | ( n6349 & n6614 ) | ( ~n6604 & n6614 ) ;
  assign n6616 = ( n6349 & n6604 ) | ( n6349 & n6614 ) | ( n6604 & n6614 ) ;
  assign n6617 = ( n6604 & n6615 ) | ( n6604 & ~n6616 ) | ( n6615 & ~n6616 ) ;
  assign n6618 = ( n6351 & n6522 ) | ( n6351 & n6617 ) | ( n6522 & n6617 ) ;
  assign n6619 = ( ~n6351 & n6522 ) | ( ~n6351 & n6617 ) | ( n6522 & n6617 ) ;
  assign n6620 = ( n6351 & ~n6618 ) | ( n6351 & n6619 ) | ( ~n6618 & n6619 ) ;
  assign n6621 = ( ~n6354 & n6512 ) | ( ~n6354 & n6620 ) | ( n6512 & n6620 ) ;
  assign n6622 = ( n6354 & n6512 ) | ( n6354 & n6620 ) | ( n6512 & n6620 ) ;
  assign n6623 = ( n6354 & n6621 ) | ( n6354 & ~n6622 ) | ( n6621 & ~n6622 ) ;
  assign n6624 = n1755 & n2083 ;
  assign n6625 = x26 & n6624 ;
  assign n6626 = x92 & n1762 ;
  assign n6627 = x91 & n1759 ;
  assign n6628 = n6626 | n6627 ;
  assign n6629 = x90 & n1895 ;
  assign n6630 = n6628 | n6629 ;
  assign n6631 = ( ~x26 & n6624 ) | ( ~x26 & n6630 ) | ( n6624 & n6630 ) ;
  assign n6632 = x26 & ~n6630 ;
  assign n6633 = ( ~n6625 & n6631 ) | ( ~n6625 & n6632 ) | ( n6631 & n6632 ) ;
  assign n6634 = ( n6367 & ~n6623 ) | ( n6367 & n6633 ) | ( ~n6623 & n6633 ) ;
  assign n6635 = ( n6367 & n6623 ) | ( n6367 & n6633 ) | ( n6623 & n6633 ) ;
  assign n6636 = ( n6623 & n6634 ) | ( n6623 & ~n6635 ) | ( n6634 & ~n6635 ) ;
  assign n6637 = ( n6380 & n6502 ) | ( n6380 & n6636 ) | ( n6502 & n6636 ) ;
  assign n6638 = ( ~n6380 & n6502 ) | ( ~n6380 & n6636 ) | ( n6502 & n6636 ) ;
  assign n6639 = ( n6380 & ~n6637 ) | ( n6380 & n6638 ) | ( ~n6637 & n6638 ) ;
  assign n6640 = n1146 & n2939 ;
  assign n6641 = x20 & n6640 ;
  assign n6642 = x98 & n1153 ;
  assign n6643 = x97 & n1150 ;
  assign n6644 = n6642 | n6643 ;
  assign n6645 = x96 & n1217 ;
  assign n6646 = n6644 | n6645 ;
  assign n6647 = ( ~x20 & n6640 ) | ( ~x20 & n6646 ) | ( n6640 & n6646 ) ;
  assign n6648 = x20 & ~n6646 ;
  assign n6649 = ( ~n6641 & n6647 ) | ( ~n6641 & n6648 ) | ( n6647 & n6648 ) ;
  assign n6650 = ( n6393 & ~n6639 ) | ( n6393 & n6649 ) | ( ~n6639 & n6649 ) ;
  assign n6651 = ( n6393 & n6639 ) | ( n6393 & n6649 ) | ( n6639 & n6649 ) ;
  assign n6652 = ( n6639 & n6650 ) | ( n6639 & ~n6651 ) | ( n6650 & ~n6651 ) ;
  assign n6653 = ( n6407 & n6492 ) | ( n6407 & n6652 ) | ( n6492 & n6652 ) ;
  assign n6654 = ( ~n6407 & n6492 ) | ( ~n6407 & n6652 ) | ( n6492 & n6652 ) ;
  assign n6655 = ( n6407 & ~n6653 ) | ( n6407 & n6654 ) | ( ~n6653 & n6654 ) ;
  assign n6656 = n649 & n3957 ;
  assign n6657 = x14 & n6656 ;
  assign n6658 = x104 & n656 ;
  assign n6659 = x103 & n653 ;
  assign n6660 = n6658 | n6659 ;
  assign n6661 = x102 & n744 ;
  assign n6662 = n6660 | n6661 ;
  assign n6663 = ( ~x14 & n6656 ) | ( ~x14 & n6662 ) | ( n6656 & n6662 ) ;
  assign n6664 = x14 & ~n6662 ;
  assign n6665 = ( ~n6657 & n6663 ) | ( ~n6657 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = ( n6409 & ~n6655 ) | ( n6409 & n6665 ) | ( ~n6655 & n6665 ) ;
  assign n6667 = ( n6409 & n6655 ) | ( n6409 & n6665 ) | ( n6655 & n6665 ) ;
  assign n6668 = ( n6655 & n6666 ) | ( n6655 & ~n6667 ) | ( n6666 & ~n6667 ) ;
  assign n6669 = n449 & n4523 ;
  assign n6670 = x11 & n6669 ;
  assign n6671 = x107 & n456 ;
  assign n6672 = x106 & n453 ;
  assign n6673 = n6671 | n6672 ;
  assign n6674 = x105 & n536 ;
  assign n6675 = n6673 | n6674 ;
  assign n6676 = ( ~x11 & n6669 ) | ( ~x11 & n6675 ) | ( n6669 & n6675 ) ;
  assign n6677 = x11 & ~n6675 ;
  assign n6678 = ( ~n6670 & n6676 ) | ( ~n6670 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6679 = ( n6426 & ~n6668 ) | ( n6426 & n6678 ) | ( ~n6668 & n6678 ) ;
  assign n6680 = ( n6426 & n6668 ) | ( n6426 & n6678 ) | ( n6668 & n6678 ) ;
  assign n6681 = ( n6668 & n6679 ) | ( n6668 & ~n6680 ) | ( n6679 & ~n6680 ) ;
  assign n6682 = ( n6428 & n6482 ) | ( n6428 & n6681 ) | ( n6482 & n6681 ) ;
  assign n6683 = ( ~n6428 & n6482 ) | ( ~n6428 & n6681 ) | ( n6482 & n6681 ) ;
  assign n6684 = ( n6428 & ~n6682 ) | ( n6428 & n6683 ) | ( ~n6682 & n6683 ) ;
  assign n6685 = n206 & n5774 ;
  assign n6686 = x5 & n6685 ;
  assign n6687 = x113 & n205 ;
  assign n6688 = x112 & n201 ;
  assign n6689 = n6687 | n6688 ;
  assign n6690 = x111 & n221 ;
  assign n6691 = n6689 | n6690 ;
  assign n6692 = ( ~x5 & n6685 ) | ( ~x5 & n6691 ) | ( n6685 & n6691 ) ;
  assign n6693 = x5 & ~n6691 ;
  assign n6694 = ( ~n6686 & n6692 ) | ( ~n6686 & n6693 ) | ( n6692 & n6693 ) ;
  assign n6695 = ( n6441 & ~n6684 ) | ( n6441 & n6694 ) | ( ~n6684 & n6694 ) ;
  assign n6696 = ( n6441 & n6684 ) | ( n6441 & n6694 ) | ( n6684 & n6694 ) ;
  assign n6697 = ( n6684 & n6695 ) | ( n6684 & ~n6696 ) | ( n6695 & ~n6696 ) ;
  assign n6698 = ( n6458 & n6472 ) | ( n6458 & n6697 ) | ( n6472 & n6697 ) ;
  assign n6699 = ( ~n6458 & n6472 ) | ( ~n6458 & n6697 ) | ( n6472 & n6697 ) ;
  assign n6700 = ( n6458 & ~n6698 ) | ( n6458 & n6699 ) | ( ~n6698 & n6699 ) ;
  assign n6701 = n301 & n5347 ;
  assign n6702 = x8 & n6701 ;
  assign n6703 = x111 & n309 ;
  assign n6704 = x110 & n306 ;
  assign n6705 = n6703 | n6704 ;
  assign n6706 = x109 & n359 ;
  assign n6707 = n6705 | n6706 ;
  assign n6708 = ( ~x8 & n6701 ) | ( ~x8 & n6707 ) | ( n6701 & n6707 ) ;
  assign n6709 = x8 & ~n6707 ;
  assign n6710 = ( ~n6702 & n6708 ) | ( ~n6702 & n6709 ) | ( n6708 & n6709 ) ;
  assign n6711 = n874 & n3764 ;
  assign n6712 = x17 & n6711 ;
  assign n6713 = x102 & n881 ;
  assign n6714 = x101 & n878 ;
  assign n6715 = n6713 | n6714 ;
  assign n6716 = x100 & n959 ;
  assign n6717 = n6715 | n6716 ;
  assign n6718 = ( ~x17 & n6711 ) | ( ~x17 & n6717 ) | ( n6711 & n6717 ) ;
  assign n6719 = x17 & ~n6717 ;
  assign n6720 = ( ~n6712 & n6718 ) | ( ~n6712 & n6719 ) | ( n6718 & n6719 ) ;
  assign n6721 = n1427 & n2772 ;
  assign n6722 = x23 & n6721 ;
  assign n6723 = x96 & n1434 ;
  assign n6724 = x95 & n1431 ;
  assign n6725 = n6723 | n6724 ;
  assign n6726 = x94 & n1531 ;
  assign n6727 = n6725 | n6726 ;
  assign n6728 = ( ~x23 & n6721 ) | ( ~x23 & n6727 ) | ( n6721 & n6727 ) ;
  assign n6729 = x23 & ~n6727 ;
  assign n6730 = ( ~n6722 & n6728 ) | ( ~n6722 & n6729 ) | ( n6728 & n6729 ) ;
  assign n6731 = n1838 & n2137 ;
  assign n6732 = x29 & n6731 ;
  assign n6733 = x90 & n2144 ;
  assign n6734 = x89 & n2141 ;
  assign n6735 = n6733 | n6734 ;
  assign n6736 = x88 & n2267 ;
  assign n6737 = n6735 | n6736 ;
  assign n6738 = ( ~x29 & n6731 ) | ( ~x29 & n6737 ) | ( n6731 & n6737 ) ;
  assign n6739 = x29 & ~n6737 ;
  assign n6740 = ( ~n6732 & n6738 ) | ( ~n6732 & n6739 ) | ( n6738 & n6739 ) ;
  assign n6741 = n1190 & n2982 ;
  assign n6742 = x35 & n6741 ;
  assign n6743 = x84 & n2989 ;
  assign n6744 = x83 & n2986 ;
  assign n6745 = n6743 | n6744 ;
  assign n6746 = x82 & n3159 ;
  assign n6747 = n6745 | n6746 ;
  assign n6748 = ( ~x35 & n6741 ) | ( ~x35 & n6747 ) | ( n6741 & n6747 ) ;
  assign n6749 = x35 & ~n6747 ;
  assign n6750 = ( ~n6742 & n6748 ) | ( ~n6742 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = n697 & n4020 ;
  assign n6752 = x41 & n6751 ;
  assign n6753 = x78 & n4027 ;
  assign n6754 = x77 & n4024 ;
  assign n6755 = n6753 | n6754 ;
  assign n6756 = x76 & n4223 ;
  assign n6757 = n6755 | n6756 ;
  assign n6758 = ( ~x41 & n6751 ) | ( ~x41 & n6757 ) | ( n6751 & n6757 ) ;
  assign n6759 = x41 & ~n6757 ;
  assign n6760 = ( ~n6752 & n6758 ) | ( ~n6752 & n6759 ) | ( n6758 & n6759 ) ;
  assign n6761 = n372 & n5223 ;
  assign n6762 = x47 & n6761 ;
  assign n6763 = x72 & n5230 ;
  assign n6764 = x71 & n5227 ;
  assign n6765 = n6763 | n6764 ;
  assign n6766 = x70 & n5434 ;
  assign n6767 = n6765 | n6766 ;
  assign n6768 = ( ~x47 & n6761 ) | ( ~x47 & n6767 ) | ( n6761 & n6767 ) ;
  assign n6769 = x47 & ~n6767 ;
  assign n6770 = ( ~n6762 & n6768 ) | ( ~n6762 & n6769 ) | ( n6768 & n6769 ) ;
  assign n6771 = n240 & n5858 ;
  assign n6772 = x50 & n6771 ;
  assign n6773 = x69 & n5865 ;
  assign n6774 = x68 & n5862 ;
  assign n6775 = n6773 | n6774 ;
  assign n6776 = x67 & n6092 ;
  assign n6777 = n6775 | n6776 ;
  assign n6778 = ( ~x50 & n6771 ) | ( ~x50 & n6777 ) | ( n6771 & n6777 ) ;
  assign n6779 = x50 & ~n6777 ;
  assign n6780 = ( ~n6772 & n6778 ) | ( ~n6772 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = x66 & n6553 ;
  assign n6782 = x65 & n6550 ;
  assign n6783 = n6781 | n6782 ;
  assign n6784 = n226 & n6546 ;
  assign n6785 = n6783 | n6784 ;
  assign n6786 = ~n6309 & n6545 ;
  assign n6787 = ~n6550 & n6786 ;
  assign n6788 = x64 & n6787 ;
  assign n6789 = n6785 | n6788 ;
  assign n6790 = ~x53 & n6789 ;
  assign n6791 = ( x53 & n6556 ) | ( x53 & n6789 ) | ( n6556 & n6789 ) ;
  assign n6792 = n6556 & n6789 ;
  assign n6793 = ( n6790 & n6791 ) | ( n6790 & ~n6792 ) | ( n6791 & ~n6792 ) ;
  assign n6794 = ( n6561 & ~n6780 ) | ( n6561 & n6793 ) | ( ~n6780 & n6793 ) ;
  assign n6795 = ( n6561 & n6780 ) | ( n6561 & n6793 ) | ( n6780 & n6793 ) ;
  assign n6796 = ( n6780 & n6794 ) | ( n6780 & ~n6795 ) | ( n6794 & ~n6795 ) ;
  assign n6797 = ( n6574 & n6770 ) | ( n6574 & n6796 ) | ( n6770 & n6796 ) ;
  assign n6798 = ( ~n6574 & n6770 ) | ( ~n6574 & n6796 ) | ( n6770 & n6796 ) ;
  assign n6799 = ( n6574 & ~n6797 ) | ( n6574 & n6798 ) | ( ~n6797 & n6798 ) ;
  assign n6800 = n508 & n4625 ;
  assign n6801 = x44 & n6800 ;
  assign n6802 = x75 & n4791 ;
  assign n6803 = x74 & n4621 ;
  assign n6804 = n6802 | n6803 ;
  assign n6805 = x73 & n4795 ;
  assign n6806 = n6804 | n6805 ;
  assign n6807 = ( ~x44 & n6800 ) | ( ~x44 & n6806 ) | ( n6800 & n6806 ) ;
  assign n6808 = x44 & ~n6806 ;
  assign n6809 = ( ~n6801 & n6807 ) | ( ~n6801 & n6808 ) | ( n6807 & n6808 ) ;
  assign n6810 = ( n6576 & ~n6799 ) | ( n6576 & n6809 ) | ( ~n6799 & n6809 ) ;
  assign n6811 = ( n6576 & n6799 ) | ( n6576 & n6809 ) | ( n6799 & n6809 ) ;
  assign n6812 = ( n6799 & n6810 ) | ( n6799 & ~n6811 ) | ( n6810 & ~n6811 ) ;
  assign n6813 = ( n6589 & n6760 ) | ( n6589 & n6812 ) | ( n6760 & n6812 ) ;
  assign n6814 = ( ~n6589 & n6760 ) | ( ~n6589 & n6812 ) | ( n6760 & n6812 ) ;
  assign n6815 = ( n6589 & ~n6813 ) | ( n6589 & n6814 ) | ( ~n6813 & n6814 ) ;
  assign n6816 = n990 & n3492 ;
  assign n6817 = x38 & n6816 ;
  assign n6818 = x81 & n3499 ;
  assign n6819 = x80 & n3496 ;
  assign n6820 = n6818 | n6819 ;
  assign n6821 = x79 & n3662 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = ( ~x38 & n6816 ) | ( ~x38 & n6822 ) | ( n6816 & n6822 ) ;
  assign n6824 = x38 & ~n6822 ;
  assign n6825 = ( ~n6817 & n6823 ) | ( ~n6817 & n6824 ) | ( n6823 & n6824 ) ;
  assign n6826 = ( n6602 & ~n6815 ) | ( n6602 & n6825 ) | ( ~n6815 & n6825 ) ;
  assign n6827 = ( n6602 & n6815 ) | ( n6602 & n6825 ) | ( n6815 & n6825 ) ;
  assign n6828 = ( n6815 & n6826 ) | ( n6815 & ~n6827 ) | ( n6826 & ~n6827 ) ;
  assign n6829 = ( n6616 & n6750 ) | ( n6616 & n6828 ) | ( n6750 & n6828 ) ;
  assign n6830 = ( ~n6616 & n6750 ) | ( ~n6616 & n6828 ) | ( n6750 & n6828 ) ;
  assign n6831 = ( n6616 & ~n6829 ) | ( n6616 & n6830 ) | ( ~n6829 & n6830 ) ;
  assign n6832 = n1494 & n2545 ;
  assign n6833 = x32 & n6832 ;
  assign n6834 = x87 & n2552 ;
  assign n6835 = x86 & n2549 ;
  assign n6836 = n6834 | n6835 ;
  assign n6837 = x85 & n2696 ;
  assign n6838 = n6836 | n6837 ;
  assign n6839 = ( ~x32 & n6832 ) | ( ~x32 & n6838 ) | ( n6832 & n6838 ) ;
  assign n6840 = x32 & ~n6838 ;
  assign n6841 = ( ~n6833 & n6839 ) | ( ~n6833 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6842 = ( n6618 & ~n6831 ) | ( n6618 & n6841 ) | ( ~n6831 & n6841 ) ;
  assign n6843 = ( n6618 & n6831 ) | ( n6618 & n6841 ) | ( n6831 & n6841 ) ;
  assign n6844 = ( n6831 & n6842 ) | ( n6831 & ~n6843 ) | ( n6842 & ~n6843 ) ;
  assign n6845 = ( n6622 & n6740 ) | ( n6622 & n6844 ) | ( n6740 & n6844 ) ;
  assign n6846 = ( ~n6622 & n6740 ) | ( ~n6622 & n6844 ) | ( n6740 & n6844 ) ;
  assign n6847 = ( n6622 & ~n6845 ) | ( n6622 & n6846 ) | ( ~n6845 & n6846 ) ;
  assign n6848 = n1755 & n2220 ;
  assign n6849 = x26 & n6848 ;
  assign n6850 = x93 & n1762 ;
  assign n6851 = x92 & n1759 ;
  assign n6852 = n6850 | n6851 ;
  assign n6853 = x91 & n1895 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = ( ~x26 & n6848 ) | ( ~x26 & n6854 ) | ( n6848 & n6854 ) ;
  assign n6856 = x26 & ~n6854 ;
  assign n6857 = ( ~n6849 & n6855 ) | ( ~n6849 & n6856 ) | ( n6855 & n6856 ) ;
  assign n6858 = ( n6635 & ~n6847 ) | ( n6635 & n6857 ) | ( ~n6847 & n6857 ) ;
  assign n6859 = ( n6635 & n6847 ) | ( n6635 & n6857 ) | ( n6847 & n6857 ) ;
  assign n6860 = ( n6847 & n6858 ) | ( n6847 & ~n6859 ) | ( n6858 & ~n6859 ) ;
  assign n6861 = ( n6637 & n6730 ) | ( n6637 & n6860 ) | ( n6730 & n6860 ) ;
  assign n6862 = ( ~n6637 & n6730 ) | ( ~n6637 & n6860 ) | ( n6730 & n6860 ) ;
  assign n6863 = ( n6637 & ~n6861 ) | ( n6637 & n6862 ) | ( ~n6861 & n6862 ) ;
  assign n6864 = n1146 & n3248 ;
  assign n6865 = x20 & n6864 ;
  assign n6866 = x99 & n1153 ;
  assign n6867 = x98 & n1150 ;
  assign n6868 = n6866 | n6867 ;
  assign n6869 = x97 & n1217 ;
  assign n6870 = n6868 | n6869 ;
  assign n6871 = ( ~x20 & n6864 ) | ( ~x20 & n6870 ) | ( n6864 & n6870 ) ;
  assign n6872 = x20 & ~n6870 ;
  assign n6873 = ( ~n6865 & n6871 ) | ( ~n6865 & n6872 ) | ( n6871 & n6872 ) ;
  assign n6874 = ( n6651 & ~n6863 ) | ( n6651 & n6873 ) | ( ~n6863 & n6873 ) ;
  assign n6875 = ( n6651 & n6863 ) | ( n6651 & n6873 ) | ( n6863 & n6873 ) ;
  assign n6876 = ( n6863 & n6874 ) | ( n6863 & ~n6875 ) | ( n6874 & ~n6875 ) ;
  assign n6877 = ( n6653 & n6720 ) | ( n6653 & n6876 ) | ( n6720 & n6876 ) ;
  assign n6878 = ( ~n6653 & n6720 ) | ( ~n6653 & n6876 ) | ( n6720 & n6876 ) ;
  assign n6879 = ( n6653 & ~n6877 ) | ( n6653 & n6878 ) | ( ~n6877 & n6878 ) ;
  assign n6880 = n649 & n4145 ;
  assign n6881 = x14 & n6880 ;
  assign n6882 = x105 & n656 ;
  assign n6883 = x104 & n653 ;
  assign n6884 = n6882 | n6883 ;
  assign n6885 = x103 & n744 ;
  assign n6886 = n6884 | n6885 ;
  assign n6887 = ( ~x14 & n6880 ) | ( ~x14 & n6886 ) | ( n6880 & n6886 ) ;
  assign n6888 = x14 & ~n6886 ;
  assign n6889 = ( ~n6881 & n6887 ) | ( ~n6881 & n6888 ) | ( n6887 & n6888 ) ;
  assign n6890 = ( n6667 & ~n6879 ) | ( n6667 & n6889 ) | ( ~n6879 & n6889 ) ;
  assign n6891 = ( n6667 & n6879 ) | ( n6667 & n6889 ) | ( n6879 & n6889 ) ;
  assign n6892 = ( n6879 & n6890 ) | ( n6879 & ~n6891 ) | ( n6890 & ~n6891 ) ;
  assign n6893 = n449 & n4914 ;
  assign n6894 = x11 & n6893 ;
  assign n6895 = x108 & n456 ;
  assign n6896 = x107 & n453 ;
  assign n6897 = n6895 | n6896 ;
  assign n6898 = x106 & n536 ;
  assign n6899 = n6897 | n6898 ;
  assign n6900 = ( ~x11 & n6893 ) | ( ~x11 & n6899 ) | ( n6893 & n6899 ) ;
  assign n6901 = x11 & ~n6899 ;
  assign n6902 = ( ~n6894 & n6900 ) | ( ~n6894 & n6901 ) | ( n6900 & n6901 ) ;
  assign n6903 = ( n6680 & ~n6892 ) | ( n6680 & n6902 ) | ( ~n6892 & n6902 ) ;
  assign n6904 = ( n6680 & n6892 ) | ( n6680 & n6902 ) | ( n6892 & n6902 ) ;
  assign n6905 = ( n6892 & n6903 ) | ( n6892 & ~n6904 ) | ( n6903 & ~n6904 ) ;
  assign n6906 = ( n6682 & n6710 ) | ( n6682 & n6905 ) | ( n6710 & n6905 ) ;
  assign n6907 = ( ~n6682 & n6710 ) | ( ~n6682 & n6905 ) | ( n6710 & n6905 ) ;
  assign n6908 = ( n6682 & ~n6906 ) | ( n6682 & n6907 ) | ( ~n6906 & n6907 ) ;
  assign n6909 = n206 & n6002 ;
  assign n6910 = x5 & n6909 ;
  assign n6911 = x114 & n205 ;
  assign n6912 = x113 & n201 ;
  assign n6913 = n6911 | n6912 ;
  assign n6914 = x112 & n221 ;
  assign n6915 = n6913 | n6914 ;
  assign n6916 = ( ~x5 & n6909 ) | ( ~x5 & n6915 ) | ( n6909 & n6915 ) ;
  assign n6917 = x5 & ~n6915 ;
  assign n6918 = ( ~n6910 & n6916 ) | ( ~n6910 & n6917 ) | ( n6916 & n6917 ) ;
  assign n6919 = ( n6696 & n6908 ) | ( n6696 & n6918 ) | ( n6908 & n6918 ) ;
  assign n6920 = ( ~n6696 & n6908 ) | ( ~n6696 & n6918 ) | ( n6908 & n6918 ) ;
  assign n6921 = ( n6696 & ~n6919 ) | ( n6696 & n6920 ) | ( ~n6919 & n6920 ) ;
  assign n6922 = ( ~x116 & x117 ) | ( ~x116 & n6461 ) | ( x117 & n6461 ) ;
  assign n6923 = ( x116 & x117 ) | ( x116 & n6461 ) | ( x117 & n6461 ) ;
  assign n6924 = ( x116 & n6922 ) | ( x116 & ~n6923 ) | ( n6922 & ~n6923 ) ;
  assign n6925 = x0 & n6924 ;
  assign n6926 = ( x1 & x2 ) | ( x1 & n6925 ) | ( x2 & n6925 ) ;
  assign n6927 = x116 & n172 ;
  assign n6928 = x117 | n6927 ;
  assign n6929 = ( n147 & n6927 ) | ( n147 & n6928 ) | ( n6927 & n6928 ) ;
  assign n6930 = ( ~x115 & n135 ) | ( ~x115 & n174 ) | ( n135 & n174 ) ;
  assign n6931 = n6929 | n6930 ;
  assign n6932 = n6926 | n6931 ;
  assign n6933 = n6926 & n6931 ;
  assign n6934 = n6932 & ~n6933 ;
  assign n6935 = ( n6698 & ~n6921 ) | ( n6698 & n6934 ) | ( ~n6921 & n6934 ) ;
  assign n6936 = ( n6698 & n6921 ) | ( n6698 & n6934 ) | ( n6921 & n6934 ) ;
  assign n6937 = ( n6921 & n6935 ) | ( n6921 & ~n6936 ) | ( n6935 & ~n6936 ) ;
  assign n6938 = ( ~x117 & x118 ) | ( ~x117 & n6923 ) | ( x118 & n6923 ) ;
  assign n6939 = ( x117 & x118 ) | ( x117 & n6923 ) | ( x118 & n6923 ) ;
  assign n6940 = ( x117 & n6938 ) | ( x117 & ~n6939 ) | ( n6938 & ~n6939 ) ;
  assign n6941 = x0 & n6940 ;
  assign n6942 = ( x1 & x2 ) | ( x1 & n6941 ) | ( x2 & n6941 ) ;
  assign n6943 = x117 & n172 ;
  assign n6944 = x118 | n6943 ;
  assign n6945 = ( n147 & n6943 ) | ( n147 & n6944 ) | ( n6943 & n6944 ) ;
  assign n6946 = ( ~x116 & n135 ) | ( ~x116 & n174 ) | ( n135 & n174 ) ;
  assign n6947 = n6945 | n6946 ;
  assign n6948 = n6942 | n6947 ;
  assign n6949 = n6942 & n6947 ;
  assign n6950 = n6948 & ~n6949 ;
  assign n6951 = n301 & n5558 ;
  assign n6952 = x8 & n6951 ;
  assign n6953 = x112 & n309 ;
  assign n6954 = x111 & n306 ;
  assign n6955 = n6953 | n6954 ;
  assign n6956 = x110 & n359 ;
  assign n6957 = n6955 | n6956 ;
  assign n6958 = ( ~x8 & n6951 ) | ( ~x8 & n6957 ) | ( n6951 & n6957 ) ;
  assign n6959 = x8 & ~n6957 ;
  assign n6960 = ( ~n6952 & n6958 ) | ( ~n6952 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = n449 & n4930 ;
  assign n6962 = x11 & n6961 ;
  assign n6963 = x109 & n456 ;
  assign n6964 = x108 & n453 ;
  assign n6965 = n6963 | n6964 ;
  assign n6966 = x107 & n536 ;
  assign n6967 = n6965 | n6966 ;
  assign n6968 = ( ~x11 & n6961 ) | ( ~x11 & n6967 ) | ( n6961 & n6967 ) ;
  assign n6969 = x11 & ~n6967 ;
  assign n6970 = ( ~n6962 & n6968 ) | ( ~n6962 & n6969 ) | ( n6968 & n6969 ) ;
  assign n6971 = n1146 & n3264 ;
  assign n6972 = x20 & n6971 ;
  assign n6973 = x100 & n1153 ;
  assign n6974 = x99 & n1150 ;
  assign n6975 = n6973 | n6974 ;
  assign n6976 = x98 & n1217 ;
  assign n6977 = n6975 | n6976 ;
  assign n6978 = ( ~x20 & n6971 ) | ( ~x20 & n6977 ) | ( n6971 & n6977 ) ;
  assign n6979 = x20 & ~n6977 ;
  assign n6980 = ( ~n6972 & n6978 ) | ( ~n6972 & n6979 ) | ( n6978 & n6979 ) ;
  assign n6981 = n1427 & n2788 ;
  assign n6982 = x23 & n6981 ;
  assign n6983 = x97 & n1434 ;
  assign n6984 = x96 & n1431 ;
  assign n6985 = n6983 | n6984 ;
  assign n6986 = x95 & n1531 ;
  assign n6987 = n6985 | n6986 ;
  assign n6988 = ( ~x23 & n6981 ) | ( ~x23 & n6987 ) | ( n6981 & n6987 ) ;
  assign n6989 = x23 & ~n6987 ;
  assign n6990 = ( ~n6982 & n6988 ) | ( ~n6982 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6991 = n1959 & n2137 ;
  assign n6992 = x29 & n6991 ;
  assign n6993 = x91 & n2144 ;
  assign n6994 = x90 & n2141 ;
  assign n6995 = n6993 | n6994 ;
  assign n6996 = x89 & n2267 ;
  assign n6997 = n6995 | n6996 ;
  assign n6998 = ( ~x29 & n6991 ) | ( ~x29 & n6997 ) | ( n6991 & n6997 ) ;
  assign n6999 = x29 & ~n6997 ;
  assign n7000 = ( ~n6992 & n6998 ) | ( ~n6992 & n6999 ) | ( n6998 & n6999 ) ;
  assign n7001 = n1602 & n2545 ;
  assign n7002 = x32 & n7001 ;
  assign n7003 = x88 & n2552 ;
  assign n7004 = x87 & n2549 ;
  assign n7005 = n7003 | n7004 ;
  assign n7006 = x86 & n2696 ;
  assign n7007 = n7005 | n7006 ;
  assign n7008 = ( ~x32 & n7001 ) | ( ~x32 & n7007 ) | ( n7001 & n7007 ) ;
  assign n7009 = x32 & ~n7007 ;
  assign n7010 = ( ~n7002 & n7008 ) | ( ~n7002 & n7009 ) | ( n7008 & n7009 ) ;
  assign n7011 = n565 & n4625 ;
  assign n7012 = x44 & n7011 ;
  assign n7013 = x76 & n4791 ;
  assign n7014 = x75 & n4621 ;
  assign n7015 = n7013 | n7014 ;
  assign n7016 = x74 & n4795 ;
  assign n7017 = n7015 | n7016 ;
  assign n7018 = ( ~x44 & n7011 ) | ( ~x44 & n7017 ) | ( n7011 & n7017 ) ;
  assign n7019 = x44 & ~n7017 ;
  assign n7020 = ( ~n7012 & n7018 ) | ( ~n7012 & n7019 ) | ( n7018 & n7019 ) ;
  assign n7021 = x67 & n6553 ;
  assign n7022 = x66 & n6550 ;
  assign n7023 = n7021 | n7022 ;
  assign n7024 = x65 & n6787 ;
  assign n7025 = n7023 | n7024 ;
  assign n7026 = n169 & n6546 ;
  assign n7027 = n7025 | n7026 ;
  assign n7028 = x53 | n7027 ;
  assign n7029 = n6556 | n6789 ;
  assign n7030 = n7027 & n7029 ;
  assign n7031 = ( x53 & n7027 ) | ( x53 & n7029 ) | ( n7027 & n7029 ) ;
  assign n7032 = ( n7028 & n7030 ) | ( n7028 & ~n7031 ) | ( n7030 & ~n7031 ) ;
  assign n7033 = x53 & ~x54 ;
  assign n7034 = ( x53 & x54 ) | ( x53 & x64 ) | ( x54 & x64 ) ;
  assign n7035 = ( n7032 & n7033 ) | ( n7032 & n7034 ) | ( n7033 & n7034 ) ;
  assign n7036 = ( ~n7032 & n7033 ) | ( ~n7032 & n7034 ) | ( n7033 & n7034 ) ;
  assign n7037 = ( n7032 & ~n7035 ) | ( n7032 & n7036 ) | ( ~n7035 & n7036 ) ;
  assign n7038 = n276 & n5858 ;
  assign n7039 = x50 & n7038 ;
  assign n7040 = x70 & n5865 ;
  assign n7041 = x69 & n5862 ;
  assign n7042 = n7040 | n7041 ;
  assign n7043 = x68 & n6092 ;
  assign n7044 = n7042 | n7043 ;
  assign n7045 = ( ~x50 & n7038 ) | ( ~x50 & n7044 ) | ( n7038 & n7044 ) ;
  assign n7046 = x50 & ~n7044 ;
  assign n7047 = ( ~n7039 & n7045 ) | ( ~n7039 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = ( n6795 & n7037 ) | ( n6795 & n7047 ) | ( n7037 & n7047 ) ;
  assign n7049 = ( ~n6795 & n7037 ) | ( ~n6795 & n7047 ) | ( n7037 & n7047 ) ;
  assign n7050 = ( n6795 & ~n7048 ) | ( n6795 & n7049 ) | ( ~n7048 & n7049 ) ;
  assign n7051 = n388 & n5223 ;
  assign n7052 = x47 & n7051 ;
  assign n7053 = x73 & n5230 ;
  assign n7054 = x72 & n5227 ;
  assign n7055 = n7053 | n7054 ;
  assign n7056 = x71 & n5434 ;
  assign n7057 = n7055 | n7056 ;
  assign n7058 = ( ~x47 & n7051 ) | ( ~x47 & n7057 ) | ( n7051 & n7057 ) ;
  assign n7059 = x47 & ~n7057 ;
  assign n7060 = ( ~n7052 & n7058 ) | ( ~n7052 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7061 = ( n6797 & ~n7050 ) | ( n6797 & n7060 ) | ( ~n7050 & n7060 ) ;
  assign n7062 = ( n6797 & n7050 ) | ( n6797 & n7060 ) | ( n7050 & n7060 ) ;
  assign n7063 = ( n7050 & n7061 ) | ( n7050 & ~n7062 ) | ( n7061 & ~n7062 ) ;
  assign n7064 = ( n6811 & n7020 ) | ( n6811 & n7063 ) | ( n7020 & n7063 ) ;
  assign n7065 = ( ~n6811 & n7020 ) | ( ~n6811 & n7063 ) | ( n7020 & n7063 ) ;
  assign n7066 = ( n6811 & ~n7064 ) | ( n6811 & n7065 ) | ( ~n7064 & n7065 ) ;
  assign n7067 = n823 & n4020 ;
  assign n7068 = x41 & n7067 ;
  assign n7069 = x79 & n4027 ;
  assign n7070 = x78 & n4024 ;
  assign n7071 = n7069 | n7070 ;
  assign n7072 = x77 & n4223 ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = ( ~x41 & n7067 ) | ( ~x41 & n7073 ) | ( n7067 & n7073 ) ;
  assign n7075 = x41 & ~n7073 ;
  assign n7076 = ( ~n7068 & n7074 ) | ( ~n7068 & n7075 ) | ( n7074 & n7075 ) ;
  assign n7077 = ( n6813 & n7066 ) | ( n6813 & n7076 ) | ( n7066 & n7076 ) ;
  assign n7078 = ( ~n6813 & n7066 ) | ( ~n6813 & n7076 ) | ( n7066 & n7076 ) ;
  assign n7079 = ( n6813 & ~n7077 ) | ( n6813 & n7078 ) | ( ~n7077 & n7078 ) ;
  assign n7080 = n1006 & n3492 ;
  assign n7081 = x38 & n7080 ;
  assign n7082 = x82 & n3499 ;
  assign n7083 = x81 & n3496 ;
  assign n7084 = n7082 | n7083 ;
  assign n7085 = x80 & n3662 ;
  assign n7086 = n7084 | n7085 ;
  assign n7087 = ( ~x38 & n7080 ) | ( ~x38 & n7086 ) | ( n7080 & n7086 ) ;
  assign n7088 = x38 & ~n7086 ;
  assign n7089 = ( ~n7081 & n7087 ) | ( ~n7081 & n7088 ) | ( n7087 & n7088 ) ;
  assign n7090 = ( ~n6827 & n7079 ) | ( ~n6827 & n7089 ) | ( n7079 & n7089 ) ;
  assign n7091 = ( n6827 & n7079 ) | ( n6827 & n7089 ) | ( n7079 & n7089 ) ;
  assign n7092 = ( n6827 & n7090 ) | ( n6827 & ~n7091 ) | ( n7090 & ~n7091 ) ;
  assign n7093 = n1368 & n2982 ;
  assign n7094 = x35 & n7093 ;
  assign n7095 = x85 & n2989 ;
  assign n7096 = x84 & n2986 ;
  assign n7097 = n7095 | n7096 ;
  assign n7098 = x83 & n3159 ;
  assign n7099 = n7097 | n7098 ;
  assign n7100 = ( ~x35 & n7093 ) | ( ~x35 & n7099 ) | ( n7093 & n7099 ) ;
  assign n7101 = x35 & ~n7099 ;
  assign n7102 = ( ~n7094 & n7100 ) | ( ~n7094 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7103 = ( n6829 & ~n7092 ) | ( n6829 & n7102 ) | ( ~n7092 & n7102 ) ;
  assign n7104 = ( n6829 & n7092 ) | ( n6829 & n7102 ) | ( n7092 & n7102 ) ;
  assign n7105 = ( n7092 & n7103 ) | ( n7092 & ~n7104 ) | ( n7103 & ~n7104 ) ;
  assign n7106 = ( n6843 & n7010 ) | ( n6843 & n7105 ) | ( n7010 & n7105 ) ;
  assign n7107 = ( ~n6843 & n7010 ) | ( ~n6843 & n7105 ) | ( n7010 & n7105 ) ;
  assign n7108 = ( n6843 & ~n7106 ) | ( n6843 & n7107 ) | ( ~n7106 & n7107 ) ;
  assign n7109 = ( ~n6845 & n7000 ) | ( ~n6845 & n7108 ) | ( n7000 & n7108 ) ;
  assign n7110 = ( n6845 & n7000 ) | ( n6845 & n7108 ) | ( n7000 & n7108 ) ;
  assign n7111 = ( n6845 & n7109 ) | ( n6845 & ~n7110 ) | ( n7109 & ~n7110 ) ;
  assign n7112 = n1755 & n2476 ;
  assign n7113 = x26 & n7112 ;
  assign n7114 = x94 & n1762 ;
  assign n7115 = x93 & n1759 ;
  assign n7116 = n7114 | n7115 ;
  assign n7117 = x92 & n1895 ;
  assign n7118 = n7116 | n7117 ;
  assign n7119 = ( ~x26 & n7112 ) | ( ~x26 & n7118 ) | ( n7112 & n7118 ) ;
  assign n7120 = x26 & ~n7118 ;
  assign n7121 = ( ~n7113 & n7119 ) | ( ~n7113 & n7120 ) | ( n7119 & n7120 ) ;
  assign n7122 = ( n6859 & ~n7111 ) | ( n6859 & n7121 ) | ( ~n7111 & n7121 ) ;
  assign n7123 = ( n6859 & n7111 ) | ( n6859 & n7121 ) | ( n7111 & n7121 ) ;
  assign n7124 = ( n7111 & n7122 ) | ( n7111 & ~n7123 ) | ( n7122 & ~n7123 ) ;
  assign n7125 = ( n6861 & n6990 ) | ( n6861 & n7124 ) | ( n6990 & n7124 ) ;
  assign n7126 = ( ~n6861 & n6990 ) | ( ~n6861 & n7124 ) | ( n6990 & n7124 ) ;
  assign n7127 = ( n6861 & ~n7125 ) | ( n6861 & n7126 ) | ( ~n7125 & n7126 ) ;
  assign n7128 = ( n6875 & n6980 ) | ( n6875 & n7127 ) | ( n6980 & n7127 ) ;
  assign n7129 = ( ~n6875 & n6980 ) | ( ~n6875 & n7127 ) | ( n6980 & n7127 ) ;
  assign n7130 = ( n6875 & ~n7128 ) | ( n6875 & n7129 ) | ( ~n7128 & n7129 ) ;
  assign n7131 = n874 & n3941 ;
  assign n7132 = x17 & n7131 ;
  assign n7133 = x103 & n881 ;
  assign n7134 = x102 & n878 ;
  assign n7135 = n7133 | n7134 ;
  assign n7136 = x101 & n959 ;
  assign n7137 = n7135 | n7136 ;
  assign n7138 = ( ~x17 & n7131 ) | ( ~x17 & n7137 ) | ( n7131 & n7137 ) ;
  assign n7139 = x17 & ~n7137 ;
  assign n7140 = ( ~n7132 & n7138 ) | ( ~n7132 & n7139 ) | ( n7138 & n7139 ) ;
  assign n7141 = ( n6877 & n7130 ) | ( n6877 & n7140 ) | ( n7130 & n7140 ) ;
  assign n7142 = ( ~n6877 & n7130 ) | ( ~n6877 & n7140 ) | ( n7130 & n7140 ) ;
  assign n7143 = ( n6877 & ~n7141 ) | ( n6877 & n7142 ) | ( ~n7141 & n7142 ) ;
  assign n7144 = n649 & n4331 ;
  assign n7145 = x14 & n7144 ;
  assign n7146 = x106 & n656 ;
  assign n7147 = x105 & n653 ;
  assign n7148 = n7146 | n7147 ;
  assign n7149 = x104 & n744 ;
  assign n7150 = n7148 | n7149 ;
  assign n7151 = ( ~x14 & n7144 ) | ( ~x14 & n7150 ) | ( n7144 & n7150 ) ;
  assign n7152 = x14 & ~n7150 ;
  assign n7153 = ( ~n7145 & n7151 ) | ( ~n7145 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7154 = ( ~n6891 & n7143 ) | ( ~n6891 & n7153 ) | ( n7143 & n7153 ) ;
  assign n7155 = ( n6891 & n7143 ) | ( n6891 & n7153 ) | ( n7143 & n7153 ) ;
  assign n7156 = ( n6891 & n7154 ) | ( n6891 & ~n7155 ) | ( n7154 & ~n7155 ) ;
  assign n7157 = ( n6904 & ~n6970 ) | ( n6904 & n7156 ) | ( ~n6970 & n7156 ) ;
  assign n7158 = ( n6904 & n6970 ) | ( n6904 & n7156 ) | ( n6970 & n7156 ) ;
  assign n7159 = ( n6970 & n7157 ) | ( n6970 & ~n7158 ) | ( n7157 & ~n7158 ) ;
  assign n7160 = ( n6906 & n6960 ) | ( n6906 & n7159 ) | ( n6960 & n7159 ) ;
  assign n7161 = ( ~n6906 & n6960 ) | ( ~n6906 & n7159 ) | ( n6960 & n7159 ) ;
  assign n7162 = ( n6906 & ~n7160 ) | ( n6906 & n7161 ) | ( ~n7160 & n7161 ) ;
  assign n7163 = n206 & n6446 ;
  assign n7164 = x5 & n7163 ;
  assign n7165 = x115 & n205 ;
  assign n7166 = x114 & n201 ;
  assign n7167 = n7165 | n7166 ;
  assign n7168 = x113 & n221 ;
  assign n7169 = n7167 | n7168 ;
  assign n7170 = ( ~x5 & n7163 ) | ( ~x5 & n7169 ) | ( n7163 & n7169 ) ;
  assign n7171 = x5 & ~n7169 ;
  assign n7172 = ( ~n7164 & n7170 ) | ( ~n7164 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7173 = ( n6919 & ~n7162 ) | ( n6919 & n7172 ) | ( ~n7162 & n7172 ) ;
  assign n7174 = ( n6919 & n7162 ) | ( n6919 & n7172 ) | ( n7162 & n7172 ) ;
  assign n7175 = ( n7162 & n7173 ) | ( n7162 & ~n7174 ) | ( n7173 & ~n7174 ) ;
  assign n7176 = ( n6936 & n6950 ) | ( n6936 & n7175 ) | ( n6950 & n7175 ) ;
  assign n7177 = ( ~n6936 & n6950 ) | ( ~n6936 & n7175 ) | ( n6950 & n7175 ) ;
  assign n7178 = ( n6936 & ~n7176 ) | ( n6936 & n7177 ) | ( ~n7176 & n7177 ) ;
  assign n7179 = ( ~x118 & x119 ) | ( ~x118 & n6939 ) | ( x119 & n6939 ) ;
  assign n7180 = ( x118 & x119 ) | ( x118 & n6939 ) | ( x119 & n6939 ) ;
  assign n7181 = ( x118 & n7179 ) | ( x118 & ~n7180 ) | ( n7179 & ~n7180 ) ;
  assign n7182 = x0 & n7181 ;
  assign n7183 = ( x1 & x2 ) | ( x1 & n7182 ) | ( x2 & n7182 ) ;
  assign n7184 = x118 & n172 ;
  assign n7185 = x119 | n7184 ;
  assign n7186 = ( n147 & n7184 ) | ( n147 & n7185 ) | ( n7184 & n7185 ) ;
  assign n7187 = ( ~x117 & n135 ) | ( ~x117 & n174 ) | ( n135 & n174 ) ;
  assign n7188 = n7186 | n7187 ;
  assign n7189 = n7183 | n7188 ;
  assign n7190 = n7183 & n7188 ;
  assign n7191 = n7189 & ~n7190 ;
  assign n7192 = n649 & n4523 ;
  assign n7193 = x14 & n7192 ;
  assign n7194 = x107 & n656 ;
  assign n7195 = x106 & n653 ;
  assign n7196 = n7194 | n7195 ;
  assign n7197 = x105 & n744 ;
  assign n7198 = n7196 | n7197 ;
  assign n7199 = ( ~x14 & n7192 ) | ( ~x14 & n7198 ) | ( n7192 & n7198 ) ;
  assign n7200 = x14 & ~n7198 ;
  assign n7201 = ( ~n7193 & n7199 ) | ( ~n7193 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7202 = n1146 & n3591 ;
  assign n7203 = x20 & n7202 ;
  assign n7204 = x101 & n1153 ;
  assign n7205 = x100 & n1150 ;
  assign n7206 = n7204 | n7205 ;
  assign n7207 = x99 & n1217 ;
  assign n7208 = n7206 | n7207 ;
  assign n7209 = ( ~x20 & n7202 ) | ( ~x20 & n7208 ) | ( n7202 & n7208 ) ;
  assign n7210 = x20 & ~n7208 ;
  assign n7211 = ( ~n7203 & n7209 ) | ( ~n7203 & n7210 ) | ( n7209 & n7210 ) ;
  assign n7212 = n1427 & n2939 ;
  assign n7213 = x23 & n7212 ;
  assign n7214 = x98 & n1434 ;
  assign n7215 = x97 & n1431 ;
  assign n7216 = n7214 | n7215 ;
  assign n7217 = x96 & n1531 ;
  assign n7218 = n7216 | n7217 ;
  assign n7219 = ( ~x23 & n7212 ) | ( ~x23 & n7218 ) | ( n7212 & n7218 ) ;
  assign n7220 = x23 & ~n7218 ;
  assign n7221 = ( ~n7213 & n7219 ) | ( ~n7213 & n7220 ) | ( n7219 & n7220 ) ;
  assign n7222 = n2083 & n2137 ;
  assign n7223 = x29 & n7222 ;
  assign n7224 = x92 & n2144 ;
  assign n7225 = x91 & n2141 ;
  assign n7226 = n7224 | n7225 ;
  assign n7227 = x90 & n2267 ;
  assign n7228 = n7226 | n7227 ;
  assign n7229 = ( ~x29 & n7222 ) | ( ~x29 & n7228 ) | ( n7222 & n7228 ) ;
  assign n7230 = x29 & ~n7228 ;
  assign n7231 = ( ~n7223 & n7229 ) | ( ~n7223 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7232 = n1822 & n2545 ;
  assign n7233 = x32 & n7232 ;
  assign n7234 = x89 & n2552 ;
  assign n7235 = x88 & n2549 ;
  assign n7236 = n7234 | n7235 ;
  assign n7237 = x87 & n2696 ;
  assign n7238 = n7236 | n7237 ;
  assign n7239 = ( ~x32 & n7232 ) | ( ~x32 & n7238 ) | ( n7232 & n7238 ) ;
  assign n7240 = x32 & ~n7238 ;
  assign n7241 = ( ~n7233 & n7239 ) | ( ~n7233 & n7240 ) | ( n7239 & n7240 ) ;
  assign n7242 = n1093 & n3492 ;
  assign n7243 = x38 & n7242 ;
  assign n7244 = x83 & n3499 ;
  assign n7245 = x82 & n3496 ;
  assign n7246 = n7244 | n7245 ;
  assign n7247 = x81 & n3662 ;
  assign n7248 = n7246 | n7247 ;
  assign n7249 = ( ~x38 & n7242 ) | ( ~x38 & n7248 ) | ( n7242 & n7248 ) ;
  assign n7250 = x38 & ~n7248 ;
  assign n7251 = ( ~n7243 & n7249 ) | ( ~n7243 & n7250 ) | ( n7249 & n7250 ) ;
  assign n7252 = n626 & n4625 ;
  assign n7253 = x44 & n7252 ;
  assign n7254 = x77 & n4791 ;
  assign n7255 = x76 & n4621 ;
  assign n7256 = n7254 | n7255 ;
  assign n7257 = x75 & n4795 ;
  assign n7258 = n7256 | n7257 ;
  assign n7259 = ( ~x44 & n7252 ) | ( ~x44 & n7258 ) | ( n7252 & n7258 ) ;
  assign n7260 = x44 & ~n7258 ;
  assign n7261 = ( ~n7253 & n7259 ) | ( ~n7253 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = x53 & x54 ;
  assign n7263 = ( x54 & n7033 ) | ( x54 & ~n7262 ) | ( n7033 & ~n7262 ) ;
  assign n7264 = x64 & n7263 ;
  assign n7265 = ~x53 & n7264 ;
  assign n7266 = n7027 & ~n7265 ;
  assign n7267 = x53 & x64 ;
  assign n7268 = ( x54 & ~n7266 ) | ( x54 & n7267 ) | ( ~n7266 & n7267 ) ;
  assign n7269 = ~x54 & n7268 ;
  assign n7270 = ( n7032 & ~n7266 ) | ( n7032 & n7269 ) | ( ~n7266 & n7269 ) ;
  assign n7271 = ~x53 & x55 ;
  assign n7272 = x54 & x55 ;
  assign n7273 = ( n7262 & n7271 ) | ( n7262 & ~n7272 ) | ( n7271 & ~n7272 ) ;
  assign n7274 = x55 & x56 ;
  assign n7275 = x55 | x56 ;
  assign n7276 = ~n7274 & n7275 ;
  assign n7277 = n7263 & n7276 ;
  assign n7278 = x65 & ~n7273 ;
  assign n7279 = ( n7273 & n7277 ) | ( n7273 & ~n7278 ) | ( n7277 & ~n7278 ) ;
  assign n7280 = x64 & n7279 ;
  assign n7281 = ( x65 & n138 ) | ( x65 & ~n7276 ) | ( n138 & ~n7276 ) ;
  assign n7282 = n7263 & n7281 ;
  assign n7283 = n7280 | n7282 ;
  assign n7284 = x56 | n7283 ;
  assign n7285 = ~n7264 & n7283 ;
  assign n7286 = ( x56 & ~n7264 ) | ( x56 & n7283 ) | ( ~n7264 & n7283 ) ;
  assign n7287 = ( n7284 & n7285 ) | ( n7284 & ~n7286 ) | ( n7285 & ~n7286 ) ;
  assign n7288 = n193 & n6546 ;
  assign n7289 = x53 & n7288 ;
  assign n7290 = x68 & n6553 ;
  assign n7291 = x67 & n6550 ;
  assign n7292 = n7290 | n7291 ;
  assign n7293 = x66 & n6787 ;
  assign n7294 = n7292 | n7293 ;
  assign n7295 = ( ~x53 & n7288 ) | ( ~x53 & n7294 ) | ( n7288 & n7294 ) ;
  assign n7296 = x53 & ~n7294 ;
  assign n7297 = ( ~n7289 & n7295 ) | ( ~n7289 & n7296 ) | ( n7295 & n7296 ) ;
  assign n7298 = ( n7270 & n7287 ) | ( n7270 & n7297 ) | ( n7287 & n7297 ) ;
  assign n7299 = ( ~n7270 & n7287 ) | ( ~n7270 & n7297 ) | ( n7287 & n7297 ) ;
  assign n7300 = ( n7270 & ~n7298 ) | ( n7270 & n7299 ) | ( ~n7298 & n7299 ) ;
  assign n7301 = n322 & n5858 ;
  assign n7302 = x50 & n7301 ;
  assign n7303 = x71 & n5865 ;
  assign n7304 = x70 & n5862 ;
  assign n7305 = n7303 | n7304 ;
  assign n7306 = x69 & n6092 ;
  assign n7307 = n7305 | n7306 ;
  assign n7308 = ( ~x50 & n7301 ) | ( ~x50 & n7307 ) | ( n7301 & n7307 ) ;
  assign n7309 = x50 & ~n7307 ;
  assign n7310 = ( ~n7302 & n7308 ) | ( ~n7302 & n7309 ) | ( n7308 & n7309 ) ;
  assign n7311 = ( n7048 & n7300 ) | ( n7048 & n7310 ) | ( n7300 & n7310 ) ;
  assign n7312 = ( ~n7048 & n7300 ) | ( ~n7048 & n7310 ) | ( n7300 & n7310 ) ;
  assign n7313 = ( n7048 & ~n7311 ) | ( n7048 & n7312 ) | ( ~n7311 & n7312 ) ;
  assign n7314 = n436 & n5223 ;
  assign n7315 = x47 & n7314 ;
  assign n7316 = x74 & n5230 ;
  assign n7317 = x73 & n5227 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = x72 & n5434 ;
  assign n7320 = n7318 | n7319 ;
  assign n7321 = ( ~x47 & n7314 ) | ( ~x47 & n7320 ) | ( n7314 & n7320 ) ;
  assign n7322 = x47 & ~n7320 ;
  assign n7323 = ( ~n7315 & n7321 ) | ( ~n7315 & n7322 ) | ( n7321 & n7322 ) ;
  assign n7324 = ( n7062 & ~n7313 ) | ( n7062 & n7323 ) | ( ~n7313 & n7323 ) ;
  assign n7325 = ( n7062 & n7313 ) | ( n7062 & n7323 ) | ( n7313 & n7323 ) ;
  assign n7326 = ( n7313 & n7324 ) | ( n7313 & ~n7325 ) | ( n7324 & ~n7325 ) ;
  assign n7327 = ( n7064 & n7261 ) | ( n7064 & n7326 ) | ( n7261 & n7326 ) ;
  assign n7328 = ( ~n7064 & n7261 ) | ( ~n7064 & n7326 ) | ( n7261 & n7326 ) ;
  assign n7329 = ( n7064 & ~n7327 ) | ( n7064 & n7328 ) | ( ~n7327 & n7328 ) ;
  assign n7330 = n840 & n4020 ;
  assign n7331 = x41 & n7330 ;
  assign n7332 = x80 & n4027 ;
  assign n7333 = x79 & n4024 ;
  assign n7334 = n7332 | n7333 ;
  assign n7335 = x78 & n4223 ;
  assign n7336 = n7334 | n7335 ;
  assign n7337 = ( ~x41 & n7330 ) | ( ~x41 & n7336 ) | ( n7330 & n7336 ) ;
  assign n7338 = x41 & ~n7336 ;
  assign n7339 = ( ~n7331 & n7337 ) | ( ~n7331 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7340 = ( n7077 & ~n7329 ) | ( n7077 & n7339 ) | ( ~n7329 & n7339 ) ;
  assign n7341 = ( n7077 & n7329 ) | ( n7077 & n7339 ) | ( n7329 & n7339 ) ;
  assign n7342 = ( n7329 & n7340 ) | ( n7329 & ~n7341 ) | ( n7340 & ~n7341 ) ;
  assign n7343 = ( ~n7091 & n7251 ) | ( ~n7091 & n7342 ) | ( n7251 & n7342 ) ;
  assign n7344 = ( n7091 & n7251 ) | ( n7091 & n7342 ) | ( n7251 & n7342 ) ;
  assign n7345 = ( n7091 & n7343 ) | ( n7091 & ~n7344 ) | ( n7343 & ~n7344 ) ;
  assign n7346 = n1384 & n2982 ;
  assign n7347 = x35 & n7346 ;
  assign n7348 = x86 & n2989 ;
  assign n7349 = x85 & n2986 ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = x84 & n3159 ;
  assign n7352 = n7350 | n7351 ;
  assign n7353 = ( ~x35 & n7346 ) | ( ~x35 & n7352 ) | ( n7346 & n7352 ) ;
  assign n7354 = x35 & ~n7352 ;
  assign n7355 = ( ~n7347 & n7353 ) | ( ~n7347 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7356 = ( n7104 & ~n7345 ) | ( n7104 & n7355 ) | ( ~n7345 & n7355 ) ;
  assign n7357 = ( n7104 & n7345 ) | ( n7104 & n7355 ) | ( n7345 & n7355 ) ;
  assign n7358 = ( n7345 & n7356 ) | ( n7345 & ~n7357 ) | ( n7356 & ~n7357 ) ;
  assign n7359 = ( n7106 & n7241 ) | ( n7106 & n7358 ) | ( n7241 & n7358 ) ;
  assign n7360 = ( ~n7106 & n7241 ) | ( ~n7106 & n7358 ) | ( n7241 & n7358 ) ;
  assign n7361 = ( n7106 & ~n7359 ) | ( n7106 & n7360 ) | ( ~n7359 & n7360 ) ;
  assign n7362 = ( n7110 & n7231 ) | ( n7110 & n7361 ) | ( n7231 & n7361 ) ;
  assign n7363 = ( ~n7110 & n7231 ) | ( ~n7110 & n7361 ) | ( n7231 & n7361 ) ;
  assign n7364 = ( n7110 & ~n7362 ) | ( n7110 & n7363 ) | ( ~n7362 & n7363 ) ;
  assign n7365 = n1755 & n2492 ;
  assign n7366 = x26 & n7365 ;
  assign n7367 = x95 & n1762 ;
  assign n7368 = x94 & n1759 ;
  assign n7369 = n7367 | n7368 ;
  assign n7370 = x93 & n1895 ;
  assign n7371 = n7369 | n7370 ;
  assign n7372 = ( ~x26 & n7365 ) | ( ~x26 & n7371 ) | ( n7365 & n7371 ) ;
  assign n7373 = x26 & ~n7371 ;
  assign n7374 = ( ~n7366 & n7372 ) | ( ~n7366 & n7373 ) | ( n7372 & n7373 ) ;
  assign n7375 = ( n7123 & ~n7364 ) | ( n7123 & n7374 ) | ( ~n7364 & n7374 ) ;
  assign n7376 = ( n7123 & n7364 ) | ( n7123 & n7374 ) | ( n7364 & n7374 ) ;
  assign n7377 = ( n7364 & n7375 ) | ( n7364 & ~n7376 ) | ( n7375 & ~n7376 ) ;
  assign n7378 = ( n7125 & n7221 ) | ( n7125 & n7377 ) | ( n7221 & n7377 ) ;
  assign n7379 = ( ~n7125 & n7221 ) | ( ~n7125 & n7377 ) | ( n7221 & n7377 ) ;
  assign n7380 = ( n7125 & ~n7378 ) | ( n7125 & n7379 ) | ( ~n7378 & n7379 ) ;
  assign n7381 = ( n7128 & n7211 ) | ( n7128 & n7380 ) | ( n7211 & n7380 ) ;
  assign n7382 = ( ~n7128 & n7211 ) | ( ~n7128 & n7380 ) | ( n7211 & n7380 ) ;
  assign n7383 = ( n7128 & ~n7381 ) | ( n7128 & n7382 ) | ( ~n7381 & n7382 ) ;
  assign n7384 = n874 & n3957 ;
  assign n7385 = x17 & n7384 ;
  assign n7386 = x104 & n881 ;
  assign n7387 = x103 & n878 ;
  assign n7388 = n7386 | n7387 ;
  assign n7389 = x102 & n959 ;
  assign n7390 = n7388 | n7389 ;
  assign n7391 = ( ~x17 & n7384 ) | ( ~x17 & n7390 ) | ( n7384 & n7390 ) ;
  assign n7392 = x17 & ~n7390 ;
  assign n7393 = ( ~n7385 & n7391 ) | ( ~n7385 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7394 = ( n7141 & ~n7383 ) | ( n7141 & n7393 ) | ( ~n7383 & n7393 ) ;
  assign n7395 = ( n7141 & n7383 ) | ( n7141 & n7393 ) | ( n7383 & n7393 ) ;
  assign n7396 = ( n7383 & n7394 ) | ( n7383 & ~n7395 ) | ( n7394 & ~n7395 ) ;
  assign n7397 = ( n7155 & n7201 ) | ( n7155 & n7396 ) | ( n7201 & n7396 ) ;
  assign n7398 = ( ~n7155 & n7201 ) | ( ~n7155 & n7396 ) | ( n7201 & n7396 ) ;
  assign n7399 = ( n7155 & ~n7397 ) | ( n7155 & n7398 ) | ( ~n7397 & n7398 ) ;
  assign n7400 = n449 & n5331 ;
  assign n7401 = x11 & n7400 ;
  assign n7402 = x110 & n456 ;
  assign n7403 = x109 & n453 ;
  assign n7404 = n7402 | n7403 ;
  assign n7405 = x108 & n536 ;
  assign n7406 = n7404 | n7405 ;
  assign n7407 = ( ~x11 & n7400 ) | ( ~x11 & n7406 ) | ( n7400 & n7406 ) ;
  assign n7408 = x11 & ~n7406 ;
  assign n7409 = ( ~n7401 & n7407 ) | ( ~n7401 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = ( n7158 & n7399 ) | ( n7158 & n7409 ) | ( n7399 & n7409 ) ;
  assign n7411 = ( ~n7158 & n7399 ) | ( ~n7158 & n7409 ) | ( n7399 & n7409 ) ;
  assign n7412 = ( n7158 & ~n7410 ) | ( n7158 & n7411 ) | ( ~n7410 & n7411 ) ;
  assign n7413 = n301 & n5774 ;
  assign n7414 = x8 & n7413 ;
  assign n7415 = x113 & n309 ;
  assign n7416 = x112 & n306 ;
  assign n7417 = n7415 | n7416 ;
  assign n7418 = x111 & n359 ;
  assign n7419 = n7417 | n7418 ;
  assign n7420 = ( ~x8 & n7413 ) | ( ~x8 & n7419 ) | ( n7413 & n7419 ) ;
  assign n7421 = x8 & ~n7419 ;
  assign n7422 = ( ~n7414 & n7420 ) | ( ~n7414 & n7421 ) | ( n7420 & n7421 ) ;
  assign n7423 = ( n7160 & ~n7412 ) | ( n7160 & n7422 ) | ( ~n7412 & n7422 ) ;
  assign n7424 = ( n7160 & n7412 ) | ( n7160 & n7422 ) | ( n7412 & n7422 ) ;
  assign n7425 = ( n7412 & n7423 ) | ( n7412 & ~n7424 ) | ( n7423 & ~n7424 ) ;
  assign n7426 = n206 & n6462 ;
  assign n7427 = x5 & n7426 ;
  assign n7428 = x116 & n205 ;
  assign n7429 = x115 & n201 ;
  assign n7430 = n7428 | n7429 ;
  assign n7431 = x114 & n221 ;
  assign n7432 = n7430 | n7431 ;
  assign n7433 = ( ~x5 & n7426 ) | ( ~x5 & n7432 ) | ( n7426 & n7432 ) ;
  assign n7434 = x5 & ~n7432 ;
  assign n7435 = ( ~n7427 & n7433 ) | ( ~n7427 & n7434 ) | ( n7433 & n7434 ) ;
  assign n7436 = ( n7174 & ~n7425 ) | ( n7174 & n7435 ) | ( ~n7425 & n7435 ) ;
  assign n7437 = ( n7174 & n7425 ) | ( n7174 & n7435 ) | ( n7425 & n7435 ) ;
  assign n7438 = ( n7425 & n7436 ) | ( n7425 & ~n7437 ) | ( n7436 & ~n7437 ) ;
  assign n7439 = ( n7176 & n7191 ) | ( n7176 & n7438 ) | ( n7191 & n7438 ) ;
  assign n7440 = ( ~n7176 & n7191 ) | ( ~n7176 & n7438 ) | ( n7191 & n7438 ) ;
  assign n7441 = ( n7176 & ~n7439 ) | ( n7176 & n7440 ) | ( ~n7439 & n7440 ) ;
  assign n7442 = ( ~x119 & x120 ) | ( ~x119 & n7180 ) | ( x120 & n7180 ) ;
  assign n7443 = ( x119 & x120 ) | ( x119 & n7180 ) | ( x120 & n7180 ) ;
  assign n7444 = ( x119 & n7442 ) | ( x119 & ~n7443 ) | ( n7442 & ~n7443 ) ;
  assign n7445 = x0 & n7444 ;
  assign n7446 = ( x1 & x2 ) | ( x1 & n7445 ) | ( x2 & n7445 ) ;
  assign n7447 = x119 & n172 ;
  assign n7448 = x120 | n7447 ;
  assign n7449 = ( n147 & n7447 ) | ( n147 & n7448 ) | ( n7447 & n7448 ) ;
  assign n7450 = ( ~x118 & n135 ) | ( ~x118 & n174 ) | ( n135 & n174 ) ;
  assign n7451 = n7449 | n7450 ;
  assign n7452 = n7446 | n7451 ;
  assign n7453 = n7446 & n7451 ;
  assign n7454 = n7452 & ~n7453 ;
  assign n7455 = n206 & n6924 ;
  assign n7456 = x5 & n7455 ;
  assign n7457 = x117 & n205 ;
  assign n7458 = x116 & n201 ;
  assign n7459 = n7457 | n7458 ;
  assign n7460 = x115 & n221 ;
  assign n7461 = n7459 | n7460 ;
  assign n7462 = ( ~x5 & n7455 ) | ( ~x5 & n7461 ) | ( n7455 & n7461 ) ;
  assign n7463 = x5 & ~n7461 ;
  assign n7464 = ( ~n7456 & n7462 ) | ( ~n7456 & n7463 ) | ( n7462 & n7463 ) ;
  assign n7465 = n301 & n6002 ;
  assign n7466 = x8 & n7465 ;
  assign n7467 = x114 & n309 ;
  assign n7468 = x113 & n306 ;
  assign n7469 = n7467 | n7468 ;
  assign n7470 = x112 & n359 ;
  assign n7471 = n7469 | n7470 ;
  assign n7472 = ( ~x8 & n7465 ) | ( ~x8 & n7471 ) | ( n7465 & n7471 ) ;
  assign n7473 = x8 & ~n7471 ;
  assign n7474 = ( ~n7466 & n7472 ) | ( ~n7466 & n7473 ) | ( n7472 & n7473 ) ;
  assign n7475 = n874 & n4145 ;
  assign n7476 = x17 & n7475 ;
  assign n7477 = x105 & n881 ;
  assign n7478 = x104 & n878 ;
  assign n7479 = n7477 | n7478 ;
  assign n7480 = x103 & n959 ;
  assign n7481 = n7479 | n7480 ;
  assign n7482 = ( ~x17 & n7475 ) | ( ~x17 & n7481 ) | ( n7475 & n7481 ) ;
  assign n7483 = x17 & ~n7481 ;
  assign n7484 = ( ~n7476 & n7482 ) | ( ~n7476 & n7483 ) | ( n7482 & n7483 ) ;
  assign n7485 = n2137 & n2220 ;
  assign n7486 = x29 & n7485 ;
  assign n7487 = x93 & n2144 ;
  assign n7488 = x92 & n2141 ;
  assign n7489 = n7487 | n7488 ;
  assign n7490 = x91 & n2267 ;
  assign n7491 = n7489 | n7490 ;
  assign n7492 = ( ~x29 & n7485 ) | ( ~x29 & n7491 ) | ( n7485 & n7491 ) ;
  assign n7493 = x29 & ~n7491 ;
  assign n7494 = ( ~n7486 & n7492 ) | ( ~n7486 & n7493 ) | ( n7492 & n7493 ) ;
  assign n7495 = n1838 & n2545 ;
  assign n7496 = x32 & n7495 ;
  assign n7497 = x90 & n2552 ;
  assign n7498 = x89 & n2549 ;
  assign n7499 = n7497 | n7498 ;
  assign n7500 = x88 & n2696 ;
  assign n7501 = n7499 | n7500 ;
  assign n7502 = ( ~x32 & n7495 ) | ( ~x32 & n7501 ) | ( n7495 & n7501 ) ;
  assign n7503 = x32 & ~n7501 ;
  assign n7504 = ( ~n7496 & n7502 ) | ( ~n7496 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7505 = n1190 & n3492 ;
  assign n7506 = x38 & n7505 ;
  assign n7507 = x84 & n3499 ;
  assign n7508 = x83 & n3496 ;
  assign n7509 = n7507 | n7508 ;
  assign n7510 = x82 & n3662 ;
  assign n7511 = n7509 | n7510 ;
  assign n7512 = ( ~x38 & n7505 ) | ( ~x38 & n7511 ) | ( n7505 & n7511 ) ;
  assign n7513 = x38 & ~n7511 ;
  assign n7514 = ( ~n7506 & n7512 ) | ( ~n7506 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7515 = n508 & n5223 ;
  assign n7516 = x47 & n7515 ;
  assign n7517 = x75 & n5230 ;
  assign n7518 = x74 & n5227 ;
  assign n7519 = n7517 | n7518 ;
  assign n7520 = x73 & n5434 ;
  assign n7521 = n7519 | n7520 ;
  assign n7522 = ( ~x47 & n7515 ) | ( ~x47 & n7521 ) | ( n7515 & n7521 ) ;
  assign n7523 = x47 & ~n7521 ;
  assign n7524 = ( ~n7516 & n7522 ) | ( ~n7516 & n7523 ) | ( n7522 & n7523 ) ;
  assign n7525 = n372 & n5858 ;
  assign n7526 = x50 & n7525 ;
  assign n7527 = x72 & n5865 ;
  assign n7528 = x71 & n5862 ;
  assign n7529 = n7527 | n7528 ;
  assign n7530 = x70 & n6092 ;
  assign n7531 = n7529 | n7530 ;
  assign n7532 = ( ~x50 & n7525 ) | ( ~x50 & n7531 ) | ( n7525 & n7531 ) ;
  assign n7533 = x50 & ~n7531 ;
  assign n7534 = ( ~n7526 & n7532 ) | ( ~n7526 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = n240 & n6546 ;
  assign n7536 = x53 & n7535 ;
  assign n7537 = x69 & n6553 ;
  assign n7538 = x68 & n6550 ;
  assign n7539 = n7537 | n7538 ;
  assign n7540 = x67 & n6787 ;
  assign n7541 = n7539 | n7540 ;
  assign n7542 = ( ~x53 & n7535 ) | ( ~x53 & n7541 ) | ( n7535 & n7541 ) ;
  assign n7543 = x53 & ~n7541 ;
  assign n7544 = ( ~n7536 & n7542 ) | ( ~n7536 & n7543 ) | ( n7542 & n7543 ) ;
  assign n7545 = ( n7263 & n7274 ) | ( n7263 & ~n7275 ) | ( n7274 & ~n7275 ) ;
  assign n7546 = x66 & n7545 ;
  assign n7547 = x65 & n7273 ;
  assign n7548 = n7546 | n7547 ;
  assign n7549 = n226 & n7277 ;
  assign n7550 = n7548 | n7549 ;
  assign n7551 = ~n7263 & n7276 ;
  assign n7552 = ~n7273 & n7551 ;
  assign n7553 = x64 & n7552 ;
  assign n7554 = n7550 | n7553 ;
  assign n7555 = x56 & n7264 ;
  assign n7556 = ( x56 & n7283 ) | ( x56 & n7555 ) | ( n7283 & n7555 ) ;
  assign n7557 = ~n7554 & n7556 ;
  assign n7558 = n7554 & ~n7556 ;
  assign n7559 = n7557 | n7558 ;
  assign n7560 = ( n7298 & ~n7544 ) | ( n7298 & n7559 ) | ( ~n7544 & n7559 ) ;
  assign n7561 = ( n7298 & n7544 ) | ( n7298 & n7559 ) | ( n7544 & n7559 ) ;
  assign n7562 = ( n7544 & n7560 ) | ( n7544 & ~n7561 ) | ( n7560 & ~n7561 ) ;
  assign n7563 = ( n7311 & n7534 ) | ( n7311 & n7562 ) | ( n7534 & n7562 ) ;
  assign n7564 = ( ~n7311 & n7534 ) | ( ~n7311 & n7562 ) | ( n7534 & n7562 ) ;
  assign n7565 = ( n7311 & ~n7563 ) | ( n7311 & n7564 ) | ( ~n7563 & n7564 ) ;
  assign n7566 = ( n7325 & n7524 ) | ( n7325 & n7565 ) | ( n7524 & n7565 ) ;
  assign n7567 = ( ~n7325 & n7524 ) | ( ~n7325 & n7565 ) | ( n7524 & n7565 ) ;
  assign n7568 = ( n7325 & ~n7566 ) | ( n7325 & n7567 ) | ( ~n7566 & n7567 ) ;
  assign n7569 = n697 & n4625 ;
  assign n7570 = x44 & n7569 ;
  assign n7571 = x78 & n4791 ;
  assign n7572 = x77 & n4621 ;
  assign n7573 = n7571 | n7572 ;
  assign n7574 = x76 & n4795 ;
  assign n7575 = n7573 | n7574 ;
  assign n7576 = ( ~x44 & n7569 ) | ( ~x44 & n7575 ) | ( n7569 & n7575 ) ;
  assign n7577 = x44 & ~n7575 ;
  assign n7578 = ( ~n7570 & n7576 ) | ( ~n7570 & n7577 ) | ( n7576 & n7577 ) ;
  assign n7579 = ( n7327 & n7568 ) | ( n7327 & n7578 ) | ( n7568 & n7578 ) ;
  assign n7580 = ( ~n7327 & n7568 ) | ( ~n7327 & n7578 ) | ( n7568 & n7578 ) ;
  assign n7581 = ( n7327 & ~n7579 ) | ( n7327 & n7580 ) | ( ~n7579 & n7580 ) ;
  assign n7582 = n990 & n4020 ;
  assign n7583 = x41 & n7582 ;
  assign n7584 = x81 & n4027 ;
  assign n7585 = x80 & n4024 ;
  assign n7586 = n7584 | n7585 ;
  assign n7587 = x79 & n4223 ;
  assign n7588 = n7586 | n7587 ;
  assign n7589 = ( ~x41 & n7582 ) | ( ~x41 & n7588 ) | ( n7582 & n7588 ) ;
  assign n7590 = x41 & ~n7588 ;
  assign n7591 = ( ~n7583 & n7589 ) | ( ~n7583 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7592 = ( n7341 & ~n7581 ) | ( n7341 & n7591 ) | ( ~n7581 & n7591 ) ;
  assign n7593 = ( n7341 & n7581 ) | ( n7341 & n7591 ) | ( n7581 & n7591 ) ;
  assign n7594 = ( n7581 & n7592 ) | ( n7581 & ~n7593 ) | ( n7592 & ~n7593 ) ;
  assign n7595 = ( n7344 & n7514 ) | ( n7344 & n7594 ) | ( n7514 & n7594 ) ;
  assign n7596 = ( ~n7344 & n7514 ) | ( ~n7344 & n7594 ) | ( n7514 & n7594 ) ;
  assign n7597 = ( n7344 & ~n7595 ) | ( n7344 & n7596 ) | ( ~n7595 & n7596 ) ;
  assign n7598 = n1494 & n2982 ;
  assign n7599 = x35 & n7598 ;
  assign n7600 = x87 & n2989 ;
  assign n7601 = x86 & n2986 ;
  assign n7602 = n7600 | n7601 ;
  assign n7603 = x85 & n3159 ;
  assign n7604 = n7602 | n7603 ;
  assign n7605 = ( ~x35 & n7598 ) | ( ~x35 & n7604 ) | ( n7598 & n7604 ) ;
  assign n7606 = x35 & ~n7604 ;
  assign n7607 = ( ~n7599 & n7605 ) | ( ~n7599 & n7606 ) | ( n7605 & n7606 ) ;
  assign n7608 = ( n7357 & ~n7597 ) | ( n7357 & n7607 ) | ( ~n7597 & n7607 ) ;
  assign n7609 = ( n7357 & n7597 ) | ( n7357 & n7607 ) | ( n7597 & n7607 ) ;
  assign n7610 = ( n7597 & n7608 ) | ( n7597 & ~n7609 ) | ( n7608 & ~n7609 ) ;
  assign n7611 = ( n7359 & n7504 ) | ( n7359 & n7610 ) | ( n7504 & n7610 ) ;
  assign n7612 = ( ~n7359 & n7504 ) | ( ~n7359 & n7610 ) | ( n7504 & n7610 ) ;
  assign n7613 = ( n7359 & ~n7611 ) | ( n7359 & n7612 ) | ( ~n7611 & n7612 ) ;
  assign n7614 = ( n7362 & n7494 ) | ( n7362 & n7613 ) | ( n7494 & n7613 ) ;
  assign n7615 = ( ~n7362 & n7494 ) | ( ~n7362 & n7613 ) | ( n7494 & n7613 ) ;
  assign n7616 = ( n7362 & ~n7614 ) | ( n7362 & n7615 ) | ( ~n7614 & n7615 ) ;
  assign n7617 = n1755 & n2772 ;
  assign n7618 = x26 & n7617 ;
  assign n7619 = x96 & n1762 ;
  assign n7620 = x95 & n1759 ;
  assign n7621 = n7619 | n7620 ;
  assign n7622 = x94 & n1895 ;
  assign n7623 = n7621 | n7622 ;
  assign n7624 = ( ~x26 & n7617 ) | ( ~x26 & n7623 ) | ( n7617 & n7623 ) ;
  assign n7625 = x26 & ~n7623 ;
  assign n7626 = ( ~n7618 & n7624 ) | ( ~n7618 & n7625 ) | ( n7624 & n7625 ) ;
  assign n7627 = ( n7376 & n7616 ) | ( n7376 & n7626 ) | ( n7616 & n7626 ) ;
  assign n7628 = ( ~n7376 & n7616 ) | ( ~n7376 & n7626 ) | ( n7616 & n7626 ) ;
  assign n7629 = ( n7376 & ~n7627 ) | ( n7376 & n7628 ) | ( ~n7627 & n7628 ) ;
  assign n7630 = n1427 & n3248 ;
  assign n7631 = x23 & n7630 ;
  assign n7632 = x99 & n1434 ;
  assign n7633 = x98 & n1431 ;
  assign n7634 = n7632 | n7633 ;
  assign n7635 = x97 & n1531 ;
  assign n7636 = n7634 | n7635 ;
  assign n7637 = ( ~x23 & n7630 ) | ( ~x23 & n7636 ) | ( n7630 & n7636 ) ;
  assign n7638 = x23 & ~n7636 ;
  assign n7639 = ( ~n7631 & n7637 ) | ( ~n7631 & n7638 ) | ( n7637 & n7638 ) ;
  assign n7640 = ( n7378 & n7629 ) | ( n7378 & n7639 ) | ( n7629 & n7639 ) ;
  assign n7641 = ( ~n7378 & n7629 ) | ( ~n7378 & n7639 ) | ( n7629 & n7639 ) ;
  assign n7642 = ( n7378 & ~n7640 ) | ( n7378 & n7641 ) | ( ~n7640 & n7641 ) ;
  assign n7643 = n1146 & n3764 ;
  assign n7644 = x20 & n7643 ;
  assign n7645 = x102 & n1153 ;
  assign n7646 = x101 & n1150 ;
  assign n7647 = n7645 | n7646 ;
  assign n7648 = x100 & n1217 ;
  assign n7649 = n7647 | n7648 ;
  assign n7650 = ( ~x20 & n7643 ) | ( ~x20 & n7649 ) | ( n7643 & n7649 ) ;
  assign n7651 = x20 & ~n7649 ;
  assign n7652 = ( ~n7644 & n7650 ) | ( ~n7644 & n7651 ) | ( n7650 & n7651 ) ;
  assign n7653 = ( n7381 & ~n7642 ) | ( n7381 & n7652 ) | ( ~n7642 & n7652 ) ;
  assign n7654 = ( n7381 & n7642 ) | ( n7381 & n7652 ) | ( n7642 & n7652 ) ;
  assign n7655 = ( n7642 & n7653 ) | ( n7642 & ~n7654 ) | ( n7653 & ~n7654 ) ;
  assign n7656 = ( n7395 & n7484 ) | ( n7395 & n7655 ) | ( n7484 & n7655 ) ;
  assign n7657 = ( ~n7395 & n7484 ) | ( ~n7395 & n7655 ) | ( n7484 & n7655 ) ;
  assign n7658 = ( n7395 & ~n7656 ) | ( n7395 & n7657 ) | ( ~n7656 & n7657 ) ;
  assign n7659 = n649 & n4914 ;
  assign n7660 = x14 & n7659 ;
  assign n7661 = x108 & n656 ;
  assign n7662 = x107 & n653 ;
  assign n7663 = n7661 | n7662 ;
  assign n7664 = x106 & n744 ;
  assign n7665 = n7663 | n7664 ;
  assign n7666 = ( ~x14 & n7659 ) | ( ~x14 & n7665 ) | ( n7659 & n7665 ) ;
  assign n7667 = x14 & ~n7665 ;
  assign n7668 = ( ~n7660 & n7666 ) | ( ~n7660 & n7667 ) | ( n7666 & n7667 ) ;
  assign n7669 = ( n7397 & ~n7658 ) | ( n7397 & n7668 ) | ( ~n7658 & n7668 ) ;
  assign n7670 = ( n7397 & n7658 ) | ( n7397 & n7668 ) | ( n7658 & n7668 ) ;
  assign n7671 = ( n7658 & n7669 ) | ( n7658 & ~n7670 ) | ( n7669 & ~n7670 ) ;
  assign n7672 = n449 & n5347 ;
  assign n7673 = x11 & n7672 ;
  assign n7674 = x111 & n456 ;
  assign n7675 = x110 & n453 ;
  assign n7676 = n7674 | n7675 ;
  assign n7677 = x109 & n536 ;
  assign n7678 = n7676 | n7677 ;
  assign n7679 = ( ~x11 & n7672 ) | ( ~x11 & n7678 ) | ( n7672 & n7678 ) ;
  assign n7680 = x11 & ~n7678 ;
  assign n7681 = ( ~n7673 & n7679 ) | ( ~n7673 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7682 = ( n7410 & ~n7671 ) | ( n7410 & n7681 ) | ( ~n7671 & n7681 ) ;
  assign n7683 = ( n7410 & n7671 ) | ( n7410 & n7681 ) | ( n7671 & n7681 ) ;
  assign n7684 = ( n7671 & n7682 ) | ( n7671 & ~n7683 ) | ( n7682 & ~n7683 ) ;
  assign n7685 = ( n7424 & n7474 ) | ( n7424 & n7684 ) | ( n7474 & n7684 ) ;
  assign n7686 = ( ~n7424 & n7474 ) | ( ~n7424 & n7684 ) | ( n7474 & n7684 ) ;
  assign n7687 = ( n7424 & ~n7685 ) | ( n7424 & n7686 ) | ( ~n7685 & n7686 ) ;
  assign n7688 = ( n7437 & ~n7464 ) | ( n7437 & n7687 ) | ( ~n7464 & n7687 ) ;
  assign n7689 = ( n7437 & n7464 ) | ( n7437 & n7687 ) | ( n7464 & n7687 ) ;
  assign n7690 = ( n7464 & n7688 ) | ( n7464 & ~n7689 ) | ( n7688 & ~n7689 ) ;
  assign n7691 = ( n7439 & n7454 ) | ( n7439 & n7690 ) | ( n7454 & n7690 ) ;
  assign n7692 = ( ~n7439 & n7454 ) | ( ~n7439 & n7690 ) | ( n7454 & n7690 ) ;
  assign n7693 = ( n7439 & ~n7691 ) | ( n7439 & n7692 ) | ( ~n7691 & n7692 ) ;
  assign n7694 = ( ~x120 & x121 ) | ( ~x120 & n7443 ) | ( x121 & n7443 ) ;
  assign n7695 = ( x120 & x121 ) | ( x120 & n7443 ) | ( x121 & n7443 ) ;
  assign n7696 = ( x120 & n7694 ) | ( x120 & ~n7695 ) | ( n7694 & ~n7695 ) ;
  assign n7697 = x0 & n7696 ;
  assign n7698 = ( x1 & x2 ) | ( x1 & n7697 ) | ( x2 & n7697 ) ;
  assign n7699 = x120 & n172 ;
  assign n7700 = x121 | n7699 ;
  assign n7701 = ( n147 & n7699 ) | ( n147 & n7700 ) | ( n7699 & n7700 ) ;
  assign n7702 = ( ~x119 & n135 ) | ( ~x119 & n174 ) | ( n135 & n174 ) ;
  assign n7703 = n7701 | n7702 ;
  assign n7704 = n7698 | n7703 ;
  assign n7705 = n7698 & n7703 ;
  assign n7706 = n7704 & ~n7705 ;
  assign n7707 = n206 & n6940 ;
  assign n7708 = x5 & n7707 ;
  assign n7709 = x118 & n205 ;
  assign n7710 = x117 & n201 ;
  assign n7711 = n7709 | n7710 ;
  assign n7712 = x116 & n221 ;
  assign n7713 = n7711 | n7712 ;
  assign n7714 = ( ~x5 & n7707 ) | ( ~x5 & n7713 ) | ( n7707 & n7713 ) ;
  assign n7715 = x5 & ~n7713 ;
  assign n7716 = ( ~n7708 & n7714 ) | ( ~n7708 & n7715 ) | ( n7714 & n7715 ) ;
  assign n7717 = n301 & n6446 ;
  assign n7718 = x8 & n7717 ;
  assign n7719 = x115 & n309 ;
  assign n7720 = x114 & n306 ;
  assign n7721 = n7719 | n7720 ;
  assign n7722 = x113 & n359 ;
  assign n7723 = n7721 | n7722 ;
  assign n7724 = ( ~x8 & n7717 ) | ( ~x8 & n7723 ) | ( n7717 & n7723 ) ;
  assign n7725 = x8 & ~n7723 ;
  assign n7726 = ( ~n7718 & n7724 ) | ( ~n7718 & n7725 ) | ( n7724 & n7725 ) ;
  assign n7727 = n449 & n5558 ;
  assign n7728 = x11 & n7727 ;
  assign n7729 = x112 & n456 ;
  assign n7730 = x111 & n453 ;
  assign n7731 = n7729 | n7730 ;
  assign n7732 = x110 & n536 ;
  assign n7733 = n7731 | n7732 ;
  assign n7734 = ( ~x11 & n7727 ) | ( ~x11 & n7733 ) | ( n7727 & n7733 ) ;
  assign n7735 = x11 & ~n7733 ;
  assign n7736 = ( ~n7728 & n7734 ) | ( ~n7728 & n7735 ) | ( n7734 & n7735 ) ;
  assign n7737 = n649 & n4930 ;
  assign n7738 = x14 & n7737 ;
  assign n7739 = x109 & n656 ;
  assign n7740 = x108 & n653 ;
  assign n7741 = n7739 | n7740 ;
  assign n7742 = x107 & n744 ;
  assign n7743 = n7741 | n7742 ;
  assign n7744 = ( ~x14 & n7737 ) | ( ~x14 & n7743 ) | ( n7737 & n7743 ) ;
  assign n7745 = x14 & ~n7743 ;
  assign n7746 = ( ~n7738 & n7744 ) | ( ~n7738 & n7745 ) | ( n7744 & n7745 ) ;
  assign n7747 = n874 & n4331 ;
  assign n7748 = x17 & n7747 ;
  assign n7749 = x106 & n881 ;
  assign n7750 = x105 & n878 ;
  assign n7751 = n7749 | n7750 ;
  assign n7752 = x104 & n959 ;
  assign n7753 = n7751 | n7752 ;
  assign n7754 = ( ~x17 & n7747 ) | ( ~x17 & n7753 ) | ( n7747 & n7753 ) ;
  assign n7755 = x17 & ~n7753 ;
  assign n7756 = ( ~n7748 & n7754 ) | ( ~n7748 & n7755 ) | ( n7754 & n7755 ) ;
  assign n7757 = n1427 & n3264 ;
  assign n7758 = x23 & n7757 ;
  assign n7759 = x100 & n1434 ;
  assign n7760 = x99 & n1431 ;
  assign n7761 = n7759 | n7760 ;
  assign n7762 = x98 & n1531 ;
  assign n7763 = n7761 | n7762 ;
  assign n7764 = ( ~x23 & n7757 ) | ( ~x23 & n7763 ) | ( n7757 & n7763 ) ;
  assign n7765 = x23 & ~n7763 ;
  assign n7766 = ( ~n7758 & n7764 ) | ( ~n7758 & n7765 ) | ( n7764 & n7765 ) ;
  assign n7767 = n2137 & n2476 ;
  assign n7768 = x29 & n7767 ;
  assign n7769 = x94 & n2144 ;
  assign n7770 = x93 & n2141 ;
  assign n7771 = n7769 | n7770 ;
  assign n7772 = x92 & n2267 ;
  assign n7773 = n7771 | n7772 ;
  assign n7774 = ( ~x29 & n7767 ) | ( ~x29 & n7773 ) | ( n7767 & n7773 ) ;
  assign n7775 = x29 & ~n7773 ;
  assign n7776 = ( ~n7768 & n7774 ) | ( ~n7768 & n7775 ) | ( n7774 & n7775 ) ;
  assign n7777 = n1602 & n2982 ;
  assign n7778 = x35 & n7777 ;
  assign n7779 = x88 & n2989 ;
  assign n7780 = x87 & n2986 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = x86 & n3159 ;
  assign n7783 = n7781 | n7782 ;
  assign n7784 = ( ~x35 & n7777 ) | ( ~x35 & n7783 ) | ( n7777 & n7783 ) ;
  assign n7785 = x35 & ~n7783 ;
  assign n7786 = ( ~n7778 & n7784 ) | ( ~n7778 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7787 = n1006 & n4020 ;
  assign n7788 = x41 & n7787 ;
  assign n7789 = x82 & n4027 ;
  assign n7790 = x81 & n4024 ;
  assign n7791 = n7789 | n7790 ;
  assign n7792 = x80 & n4223 ;
  assign n7793 = n7791 | n7792 ;
  assign n7794 = ( ~x41 & n7787 ) | ( ~x41 & n7793 ) | ( n7787 & n7793 ) ;
  assign n7795 = x41 & ~n7793 ;
  assign n7796 = ( ~n7788 & n7794 ) | ( ~n7788 & n7795 ) | ( n7794 & n7795 ) ;
  assign n7797 = n565 & n5223 ;
  assign n7798 = x47 & n7797 ;
  assign n7799 = x76 & n5230 ;
  assign n7800 = x75 & n5227 ;
  assign n7801 = n7799 | n7800 ;
  assign n7802 = x74 & n5434 ;
  assign n7803 = n7801 | n7802 ;
  assign n7804 = ( ~x47 & n7797 ) | ( ~x47 & n7803 ) | ( n7797 & n7803 ) ;
  assign n7805 = x47 & ~n7803 ;
  assign n7806 = ( ~n7798 & n7804 ) | ( ~n7798 & n7805 ) | ( n7804 & n7805 ) ;
  assign n7807 = x56 & ~n7556 ;
  assign n7808 = ~n7554 & n7807 ;
  assign n7809 = x66 & n7273 ;
  assign n7810 = x56 & n7809 ;
  assign n7811 = x67 & n7545 ;
  assign n7812 = x65 & n7552 ;
  assign n7813 = n7811 | n7812 ;
  assign n7814 = n169 & n7277 ;
  assign n7815 = n7813 | n7814 ;
  assign n7816 = ( ~x56 & n7809 ) | ( ~x56 & n7815 ) | ( n7809 & n7815 ) ;
  assign n7817 = x56 & ~n7815 ;
  assign n7818 = ( ~n7810 & n7816 ) | ( ~n7810 & n7817 ) | ( n7816 & n7817 ) ;
  assign n7819 = x56 & x57 ;
  assign n7820 = x56 | x57 ;
  assign n7821 = ~n7819 & n7820 ;
  assign n7822 = x64 & n7821 ;
  assign n7823 = ( ~n7808 & n7818 ) | ( ~n7808 & n7822 ) | ( n7818 & n7822 ) ;
  assign n7824 = ( n7808 & n7818 ) | ( n7808 & n7822 ) | ( n7818 & n7822 ) ;
  assign n7825 = ( n7808 & n7823 ) | ( n7808 & ~n7824 ) | ( n7823 & ~n7824 ) ;
  assign n7826 = n276 & n6546 ;
  assign n7827 = x53 & n7826 ;
  assign n7828 = x70 & n6553 ;
  assign n7829 = x69 & n6550 ;
  assign n7830 = n7828 | n7829 ;
  assign n7831 = x68 & n6787 ;
  assign n7832 = n7830 | n7831 ;
  assign n7833 = ( ~x53 & n7826 ) | ( ~x53 & n7832 ) | ( n7826 & n7832 ) ;
  assign n7834 = x53 & ~n7832 ;
  assign n7835 = ( ~n7827 & n7833 ) | ( ~n7827 & n7834 ) | ( n7833 & n7834 ) ;
  assign n7836 = ( n7561 & n7825 ) | ( n7561 & n7835 ) | ( n7825 & n7835 ) ;
  assign n7837 = ( ~n7561 & n7825 ) | ( ~n7561 & n7835 ) | ( n7825 & n7835 ) ;
  assign n7838 = ( n7561 & ~n7836 ) | ( n7561 & n7837 ) | ( ~n7836 & n7837 ) ;
  assign n7839 = n388 & n5858 ;
  assign n7840 = x50 & n7839 ;
  assign n7841 = x73 & n5865 ;
  assign n7842 = x72 & n5862 ;
  assign n7843 = n7841 | n7842 ;
  assign n7844 = x71 & n6092 ;
  assign n7845 = n7843 | n7844 ;
  assign n7846 = ( ~x50 & n7839 ) | ( ~x50 & n7845 ) | ( n7839 & n7845 ) ;
  assign n7847 = x50 & ~n7845 ;
  assign n7848 = ( ~n7840 & n7846 ) | ( ~n7840 & n7847 ) | ( n7846 & n7847 ) ;
  assign n7849 = ( n7563 & ~n7838 ) | ( n7563 & n7848 ) | ( ~n7838 & n7848 ) ;
  assign n7850 = ( n7563 & n7838 ) | ( n7563 & n7848 ) | ( n7838 & n7848 ) ;
  assign n7851 = ( n7838 & n7849 ) | ( n7838 & ~n7850 ) | ( n7849 & ~n7850 ) ;
  assign n7852 = ( n7566 & n7806 ) | ( n7566 & n7851 ) | ( n7806 & n7851 ) ;
  assign n7853 = ( ~n7566 & n7806 ) | ( ~n7566 & n7851 ) | ( n7806 & n7851 ) ;
  assign n7854 = ( n7566 & ~n7852 ) | ( n7566 & n7853 ) | ( ~n7852 & n7853 ) ;
  assign n7855 = n823 & n4625 ;
  assign n7856 = x44 & n7855 ;
  assign n7857 = x79 & n4791 ;
  assign n7858 = x78 & n4621 ;
  assign n7859 = n7857 | n7858 ;
  assign n7860 = x77 & n4795 ;
  assign n7861 = n7859 | n7860 ;
  assign n7862 = ( ~x44 & n7855 ) | ( ~x44 & n7861 ) | ( n7855 & n7861 ) ;
  assign n7863 = x44 & ~n7861 ;
  assign n7864 = ( ~n7856 & n7862 ) | ( ~n7856 & n7863 ) | ( n7862 & n7863 ) ;
  assign n7865 = ( n7579 & ~n7854 ) | ( n7579 & n7864 ) | ( ~n7854 & n7864 ) ;
  assign n7866 = ( n7579 & n7854 ) | ( n7579 & n7864 ) | ( n7854 & n7864 ) ;
  assign n7867 = ( n7854 & n7865 ) | ( n7854 & ~n7866 ) | ( n7865 & ~n7866 ) ;
  assign n7868 = ( n7593 & n7796 ) | ( n7593 & n7867 ) | ( n7796 & n7867 ) ;
  assign n7869 = ( ~n7593 & n7796 ) | ( ~n7593 & n7867 ) | ( n7796 & n7867 ) ;
  assign n7870 = ( n7593 & ~n7868 ) | ( n7593 & n7869 ) | ( ~n7868 & n7869 ) ;
  assign n7871 = n1368 & n3492 ;
  assign n7872 = x38 & n7871 ;
  assign n7873 = x85 & n3499 ;
  assign n7874 = x84 & n3496 ;
  assign n7875 = n7873 | n7874 ;
  assign n7876 = x83 & n3662 ;
  assign n7877 = n7875 | n7876 ;
  assign n7878 = ( ~x38 & n7871 ) | ( ~x38 & n7877 ) | ( n7871 & n7877 ) ;
  assign n7879 = x38 & ~n7877 ;
  assign n7880 = ( ~n7872 & n7878 ) | ( ~n7872 & n7879 ) | ( n7878 & n7879 ) ;
  assign n7881 = ( n7595 & ~n7870 ) | ( n7595 & n7880 ) | ( ~n7870 & n7880 ) ;
  assign n7882 = ( n7595 & n7870 ) | ( n7595 & n7880 ) | ( n7870 & n7880 ) ;
  assign n7883 = ( n7870 & n7881 ) | ( n7870 & ~n7882 ) | ( n7881 & ~n7882 ) ;
  assign n7884 = ( ~n7609 & n7786 ) | ( ~n7609 & n7883 ) | ( n7786 & n7883 ) ;
  assign n7885 = ( n7609 & n7786 ) | ( n7609 & n7883 ) | ( n7786 & n7883 ) ;
  assign n7886 = ( n7609 & n7884 ) | ( n7609 & ~n7885 ) | ( n7884 & ~n7885 ) ;
  assign n7887 = n1959 & n2545 ;
  assign n7888 = x32 & n7887 ;
  assign n7889 = x91 & n2552 ;
  assign n7890 = x90 & n2549 ;
  assign n7891 = n7889 | n7890 ;
  assign n7892 = x89 & n2696 ;
  assign n7893 = n7891 | n7892 ;
  assign n7894 = ( ~x32 & n7887 ) | ( ~x32 & n7893 ) | ( n7887 & n7893 ) ;
  assign n7895 = x32 & ~n7893 ;
  assign n7896 = ( ~n7888 & n7894 ) | ( ~n7888 & n7895 ) | ( n7894 & n7895 ) ;
  assign n7897 = ( n7611 & ~n7886 ) | ( n7611 & n7896 ) | ( ~n7886 & n7896 ) ;
  assign n7898 = ( n7611 & n7886 ) | ( n7611 & n7896 ) | ( n7886 & n7896 ) ;
  assign n7899 = ( n7886 & n7897 ) | ( n7886 & ~n7898 ) | ( n7897 & ~n7898 ) ;
  assign n7900 = ( n7614 & n7776 ) | ( n7614 & n7899 ) | ( n7776 & n7899 ) ;
  assign n7901 = ( ~n7614 & n7776 ) | ( ~n7614 & n7899 ) | ( n7776 & n7899 ) ;
  assign n7902 = ( n7614 & ~n7900 ) | ( n7614 & n7901 ) | ( ~n7900 & n7901 ) ;
  assign n7903 = n1755 & n2788 ;
  assign n7904 = x26 & n7903 ;
  assign n7905 = x97 & n1762 ;
  assign n7906 = x96 & n1759 ;
  assign n7907 = n7905 | n7906 ;
  assign n7908 = x95 & n1895 ;
  assign n7909 = n7907 | n7908 ;
  assign n7910 = ( ~x26 & n7903 ) | ( ~x26 & n7909 ) | ( n7903 & n7909 ) ;
  assign n7911 = x26 & ~n7909 ;
  assign n7912 = ( ~n7904 & n7910 ) | ( ~n7904 & n7911 ) | ( n7910 & n7911 ) ;
  assign n7913 = ( n7627 & ~n7902 ) | ( n7627 & n7912 ) | ( ~n7902 & n7912 ) ;
  assign n7914 = ( n7627 & n7902 ) | ( n7627 & n7912 ) | ( n7902 & n7912 ) ;
  assign n7915 = ( n7902 & n7913 ) | ( n7902 & ~n7914 ) | ( n7913 & ~n7914 ) ;
  assign n7916 = ( n7640 & n7766 ) | ( n7640 & n7915 ) | ( n7766 & n7915 ) ;
  assign n7917 = ( ~n7640 & n7766 ) | ( ~n7640 & n7915 ) | ( n7766 & n7915 ) ;
  assign n7918 = ( n7640 & ~n7916 ) | ( n7640 & n7917 ) | ( ~n7916 & n7917 ) ;
  assign n7919 = n1146 & n3941 ;
  assign n7920 = x20 & n7919 ;
  assign n7921 = x103 & n1153 ;
  assign n7922 = x102 & n1150 ;
  assign n7923 = n7921 | n7922 ;
  assign n7924 = x101 & n1217 ;
  assign n7925 = n7923 | n7924 ;
  assign n7926 = ( ~x20 & n7919 ) | ( ~x20 & n7925 ) | ( n7919 & n7925 ) ;
  assign n7927 = x20 & ~n7925 ;
  assign n7928 = ( ~n7920 & n7926 ) | ( ~n7920 & n7927 ) | ( n7926 & n7927 ) ;
  assign n7929 = ( n7654 & ~n7918 ) | ( n7654 & n7928 ) | ( ~n7918 & n7928 ) ;
  assign n7930 = ( n7654 & n7918 ) | ( n7654 & n7928 ) | ( n7918 & n7928 ) ;
  assign n7931 = ( n7918 & n7929 ) | ( n7918 & ~n7930 ) | ( n7929 & ~n7930 ) ;
  assign n7932 = ( n7656 & n7756 ) | ( n7656 & n7931 ) | ( n7756 & n7931 ) ;
  assign n7933 = ( ~n7656 & n7756 ) | ( ~n7656 & n7931 ) | ( n7756 & n7931 ) ;
  assign n7934 = ( n7656 & ~n7932 ) | ( n7656 & n7933 ) | ( ~n7932 & n7933 ) ;
  assign n7935 = ( ~n7670 & n7746 ) | ( ~n7670 & n7934 ) | ( n7746 & n7934 ) ;
  assign n7936 = ( n7670 & n7746 ) | ( n7670 & n7934 ) | ( n7746 & n7934 ) ;
  assign n7937 = ( n7670 & n7935 ) | ( n7670 & ~n7936 ) | ( n7935 & ~n7936 ) ;
  assign n7938 = ( n7683 & ~n7736 ) | ( n7683 & n7937 ) | ( ~n7736 & n7937 ) ;
  assign n7939 = ( n7683 & n7736 ) | ( n7683 & n7937 ) | ( n7736 & n7937 ) ;
  assign n7940 = ( n7736 & n7938 ) | ( n7736 & ~n7939 ) | ( n7938 & ~n7939 ) ;
  assign n7941 = ( n7685 & n7726 ) | ( n7685 & n7940 ) | ( n7726 & n7940 ) ;
  assign n7942 = ( ~n7685 & n7726 ) | ( ~n7685 & n7940 ) | ( n7726 & n7940 ) ;
  assign n7943 = ( n7685 & ~n7941 ) | ( n7685 & n7942 ) | ( ~n7941 & n7942 ) ;
  assign n7944 = ( n7689 & ~n7716 ) | ( n7689 & n7943 ) | ( ~n7716 & n7943 ) ;
  assign n7945 = ( n7689 & n7716 ) | ( n7689 & n7943 ) | ( n7716 & n7943 ) ;
  assign n7946 = ( n7716 & n7944 ) | ( n7716 & ~n7945 ) | ( n7944 & ~n7945 ) ;
  assign n7947 = ( n7691 & n7706 ) | ( n7691 & n7946 ) | ( n7706 & n7946 ) ;
  assign n7948 = ( ~n7691 & n7706 ) | ( ~n7691 & n7946 ) | ( n7706 & n7946 ) ;
  assign n7949 = ( n7691 & ~n7947 ) | ( n7691 & n7948 ) | ( ~n7947 & n7948 ) ;
  assign n7950 = n206 & n7181 ;
  assign n7951 = x5 & n7950 ;
  assign n7952 = x119 & n205 ;
  assign n7953 = x118 & n201 ;
  assign n7954 = n7952 | n7953 ;
  assign n7955 = x117 & n221 ;
  assign n7956 = n7954 | n7955 ;
  assign n7957 = ( ~x5 & n7950 ) | ( ~x5 & n7956 ) | ( n7950 & n7956 ) ;
  assign n7958 = x5 & ~n7956 ;
  assign n7959 = ( ~n7951 & n7957 ) | ( ~n7951 & n7958 ) | ( n7957 & n7958 ) ;
  assign n7960 = n301 & n6462 ;
  assign n7961 = x8 & n7960 ;
  assign n7962 = x116 & n309 ;
  assign n7963 = x115 & n306 ;
  assign n7964 = n7962 | n7963 ;
  assign n7965 = x114 & n359 ;
  assign n7966 = n7964 | n7965 ;
  assign n7967 = ( ~x8 & n7960 ) | ( ~x8 & n7966 ) | ( n7960 & n7966 ) ;
  assign n7968 = x8 & ~n7966 ;
  assign n7969 = ( ~n7961 & n7967 ) | ( ~n7961 & n7968 ) | ( n7967 & n7968 ) ;
  assign n7970 = n649 & n5331 ;
  assign n7971 = x14 & n7970 ;
  assign n7972 = x110 & n656 ;
  assign n7973 = x109 & n653 ;
  assign n7974 = n7972 | n7973 ;
  assign n7975 = x108 & n744 ;
  assign n7976 = n7974 | n7975 ;
  assign n7977 = ( ~x14 & n7970 ) | ( ~x14 & n7976 ) | ( n7970 & n7976 ) ;
  assign n7978 = x14 & ~n7976 ;
  assign n7979 = ( ~n7971 & n7977 ) | ( ~n7971 & n7978 ) | ( n7977 & n7978 ) ;
  assign n7980 = n1146 & n3957 ;
  assign n7981 = x20 & n7980 ;
  assign n7982 = x104 & n1153 ;
  assign n7983 = x103 & n1150 ;
  assign n7984 = n7982 | n7983 ;
  assign n7985 = x102 & n1217 ;
  assign n7986 = n7984 | n7985 ;
  assign n7987 = ( ~x20 & n7980 ) | ( ~x20 & n7986 ) | ( n7980 & n7986 ) ;
  assign n7988 = x20 & ~n7986 ;
  assign n7989 = ( ~n7981 & n7987 ) | ( ~n7981 & n7988 ) | ( n7987 & n7988 ) ;
  assign n7990 = n1755 & n2939 ;
  assign n7991 = x26 & n7990 ;
  assign n7992 = x98 & n1762 ;
  assign n7993 = x97 & n1759 ;
  assign n7994 = n7992 | n7993 ;
  assign n7995 = x96 & n1895 ;
  assign n7996 = n7994 | n7995 ;
  assign n7997 = ( ~x26 & n7990 ) | ( ~x26 & n7996 ) | ( n7990 & n7996 ) ;
  assign n7998 = x26 & ~n7996 ;
  assign n7999 = ( ~n7991 & n7997 ) | ( ~n7991 & n7998 ) | ( n7997 & n7998 ) ;
  assign n8000 = n2137 & n2492 ;
  assign n8001 = x29 & n8000 ;
  assign n8002 = x95 & n2144 ;
  assign n8003 = x94 & n2141 ;
  assign n8004 = n8002 | n8003 ;
  assign n8005 = x93 & n2267 ;
  assign n8006 = n8004 | n8005 ;
  assign n8007 = ( ~x29 & n8000 ) | ( ~x29 & n8006 ) | ( n8000 & n8006 ) ;
  assign n8008 = x29 & ~n8006 ;
  assign n8009 = ( ~n8001 & n8007 ) | ( ~n8001 & n8008 ) | ( n8007 & n8008 ) ;
  assign n8010 = n1822 & n2982 ;
  assign n8011 = x35 & n8010 ;
  assign n8012 = x89 & n2989 ;
  assign n8013 = x88 & n2986 ;
  assign n8014 = n8012 | n8013 ;
  assign n8015 = x87 & n3159 ;
  assign n8016 = n8014 | n8015 ;
  assign n8017 = ( ~x35 & n8010 ) | ( ~x35 & n8016 ) | ( n8010 & n8016 ) ;
  assign n8018 = x35 & ~n8016 ;
  assign n8019 = ( ~n8011 & n8017 ) | ( ~n8011 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8020 = n1093 & n4020 ;
  assign n8021 = x41 & n8020 ;
  assign n8022 = x83 & n4027 ;
  assign n8023 = x82 & n4024 ;
  assign n8024 = n8022 | n8023 ;
  assign n8025 = x81 & n4223 ;
  assign n8026 = n8024 | n8025 ;
  assign n8027 = ( ~x41 & n8020 ) | ( ~x41 & n8026 ) | ( n8020 & n8026 ) ;
  assign n8028 = x41 & ~n8026 ;
  assign n8029 = ( ~n8021 & n8027 ) | ( ~n8021 & n8028 ) | ( n8027 & n8028 ) ;
  assign n8030 = n840 & n4625 ;
  assign n8031 = x44 & n8030 ;
  assign n8032 = x80 & n4791 ;
  assign n8033 = x79 & n4621 ;
  assign n8034 = n8032 | n8033 ;
  assign n8035 = x78 & n4795 ;
  assign n8036 = n8034 | n8035 ;
  assign n8037 = ( ~x44 & n8030 ) | ( ~x44 & n8036 ) | ( n8030 & n8036 ) ;
  assign n8038 = x44 & ~n8036 ;
  assign n8039 = ( ~n8031 & n8037 ) | ( ~n8031 & n8038 ) | ( n8037 & n8038 ) ;
  assign n8040 = ~n8029 & n8039 ;
  assign n8041 = n8029 & ~n8039 ;
  assign n8042 = n8040 | n8041 ;
  assign n8043 = n626 & n5223 ;
  assign n8044 = x47 & n8043 ;
  assign n8045 = x77 & n5230 ;
  assign n8046 = x76 & n5227 ;
  assign n8047 = n8045 | n8046 ;
  assign n8048 = x75 & n5434 ;
  assign n8049 = n8047 | n8048 ;
  assign n8050 = ( ~x47 & n8043 ) | ( ~x47 & n8049 ) | ( n8043 & n8049 ) ;
  assign n8051 = x47 & ~n8049 ;
  assign n8052 = ( ~n8044 & n8050 ) | ( ~n8044 & n8051 ) | ( n8050 & n8051 ) ;
  assign n8053 = n7818 & n7824 ;
  assign n8054 = n193 & n7277 ;
  assign n8055 = x56 & n8054 ;
  assign n8056 = x68 & n7545 ;
  assign n8057 = x67 & n7273 ;
  assign n8058 = n8056 | n8057 ;
  assign n8059 = x66 & n7552 ;
  assign n8060 = n8058 | n8059 ;
  assign n8061 = ( ~x56 & n8054 ) | ( ~x56 & n8060 ) | ( n8054 & n8060 ) ;
  assign n8062 = x56 & ~n8060 ;
  assign n8063 = ( ~n8055 & n8061 ) | ( ~n8055 & n8062 ) | ( n8061 & n8062 ) ;
  assign n8064 = x58 & x59 ;
  assign n8065 = x58 | x59 ;
  assign n8066 = ~n8064 & n8065 ;
  assign n8067 = n7821 & n8066 ;
  assign n8068 = n302 & n8067 ;
  assign n8069 = ~x56 & x58 ;
  assign n8070 = x57 & x58 ;
  assign n8071 = ( n7819 & n8069 ) | ( n7819 & ~n8070 ) | ( n8069 & ~n8070 ) ;
  assign n8072 = x64 & n8071 ;
  assign n8073 = n8068 | n8072 ;
  assign n8074 = ( n7821 & n8064 ) | ( n7821 & ~n8065 ) | ( n8064 & ~n8065 ) ;
  assign n8075 = x65 & n8074 ;
  assign n8076 = n8073 | n8075 ;
  assign n8077 = n7822 | n8076 ;
  assign n8078 = ( x59 & n7822 ) | ( x59 & ~n8076 ) | ( n7822 & ~n8076 ) ;
  assign n8079 = x59 & ~n8076 ;
  assign n8080 = ( n8077 & ~n8078 ) | ( n8077 & n8079 ) | ( ~n8078 & n8079 ) ;
  assign n8081 = ( n8053 & n8063 ) | ( n8053 & n8080 ) | ( n8063 & n8080 ) ;
  assign n8082 = ( ~n8053 & n8063 ) | ( ~n8053 & n8080 ) | ( n8063 & n8080 ) ;
  assign n8083 = ( n8053 & ~n8081 ) | ( n8053 & n8082 ) | ( ~n8081 & n8082 ) ;
  assign n8084 = n322 & n6546 ;
  assign n8085 = x53 & n8084 ;
  assign n8086 = x71 & n6553 ;
  assign n8087 = x70 & n6550 ;
  assign n8088 = n8086 | n8087 ;
  assign n8089 = x69 & n6787 ;
  assign n8090 = n8088 | n8089 ;
  assign n8091 = ( ~x53 & n8084 ) | ( ~x53 & n8090 ) | ( n8084 & n8090 ) ;
  assign n8092 = x53 & ~n8090 ;
  assign n8093 = ( ~n8085 & n8091 ) | ( ~n8085 & n8092 ) | ( n8091 & n8092 ) ;
  assign n8094 = ( n7836 & n8083 ) | ( n7836 & n8093 ) | ( n8083 & n8093 ) ;
  assign n8095 = ( ~n7836 & n8083 ) | ( ~n7836 & n8093 ) | ( n8083 & n8093 ) ;
  assign n8096 = ( n7836 & ~n8094 ) | ( n7836 & n8095 ) | ( ~n8094 & n8095 ) ;
  assign n8097 = n436 & n5858 ;
  assign n8098 = x50 & n8097 ;
  assign n8099 = x74 & n5865 ;
  assign n8100 = x73 & n5862 ;
  assign n8101 = n8099 | n8100 ;
  assign n8102 = x72 & n6092 ;
  assign n8103 = n8101 | n8102 ;
  assign n8104 = ( ~x50 & n8097 ) | ( ~x50 & n8103 ) | ( n8097 & n8103 ) ;
  assign n8105 = x50 & ~n8103 ;
  assign n8106 = ( ~n8098 & n8104 ) | ( ~n8098 & n8105 ) | ( n8104 & n8105 ) ;
  assign n8107 = ( n7850 & ~n8096 ) | ( n7850 & n8106 ) | ( ~n8096 & n8106 ) ;
  assign n8108 = ( n7850 & n8096 ) | ( n7850 & n8106 ) | ( n8096 & n8106 ) ;
  assign n8109 = ( n8096 & n8107 ) | ( n8096 & ~n8108 ) | ( n8107 & ~n8108 ) ;
  assign n8110 = ( n7852 & n8052 ) | ( n7852 & n8109 ) | ( n8052 & n8109 ) ;
  assign n8111 = ( ~n7852 & n8052 ) | ( ~n7852 & n8109 ) | ( n8052 & n8109 ) ;
  assign n8112 = ( n7852 & ~n8110 ) | ( n7852 & n8111 ) | ( ~n8110 & n8111 ) ;
  assign n8113 = n7866 & ~n8112 ;
  assign n8114 = ~n7866 & n8112 ;
  assign n8115 = n8113 | n8114 ;
  assign n8116 = ( ~n7868 & n8042 ) | ( ~n7868 & n8115 ) | ( n8042 & n8115 ) ;
  assign n8117 = ( n7868 & n8042 ) | ( n7868 & ~n8115 ) | ( n8042 & ~n8115 ) ;
  assign n8118 = ( ~n8042 & n8116 ) | ( ~n8042 & n8117 ) | ( n8116 & n8117 ) ;
  assign n8119 = n1384 & n3492 ;
  assign n8120 = x38 & n8119 ;
  assign n8121 = x86 & n3499 ;
  assign n8122 = x85 & n3496 ;
  assign n8123 = n8121 | n8122 ;
  assign n8124 = x84 & n3662 ;
  assign n8125 = n8123 | n8124 ;
  assign n8126 = ( ~x38 & n8119 ) | ( ~x38 & n8125 ) | ( n8119 & n8125 ) ;
  assign n8127 = x38 & ~n8125 ;
  assign n8128 = ( ~n8120 & n8126 ) | ( ~n8120 & n8127 ) | ( n8126 & n8127 ) ;
  assign n8129 = ( n7882 & n8118 ) | ( n7882 & n8128 ) | ( n8118 & n8128 ) ;
  assign n8130 = ( ~n7882 & n8118 ) | ( ~n7882 & n8128 ) | ( n8118 & n8128 ) ;
  assign n8131 = ( n7882 & ~n8129 ) | ( n7882 & n8130 ) | ( ~n8129 & n8130 ) ;
  assign n8132 = ( ~n7885 & n8019 ) | ( ~n7885 & n8131 ) | ( n8019 & n8131 ) ;
  assign n8133 = ( n7885 & n8019 ) | ( n7885 & n8131 ) | ( n8019 & n8131 ) ;
  assign n8134 = ( n7885 & n8132 ) | ( n7885 & ~n8133 ) | ( n8132 & ~n8133 ) ;
  assign n8135 = n2083 & n2545 ;
  assign n8136 = x32 & n8135 ;
  assign n8137 = x92 & n2552 ;
  assign n8138 = x91 & n2549 ;
  assign n8139 = n8137 | n8138 ;
  assign n8140 = x90 & n2696 ;
  assign n8141 = n8139 | n8140 ;
  assign n8142 = ( ~x32 & n8135 ) | ( ~x32 & n8141 ) | ( n8135 & n8141 ) ;
  assign n8143 = x32 & ~n8141 ;
  assign n8144 = ( ~n8136 & n8142 ) | ( ~n8136 & n8143 ) | ( n8142 & n8143 ) ;
  assign n8145 = ( n7898 & ~n8134 ) | ( n7898 & n8144 ) | ( ~n8134 & n8144 ) ;
  assign n8146 = ( n7898 & n8134 ) | ( n7898 & n8144 ) | ( n8134 & n8144 ) ;
  assign n8147 = ( n8134 & n8145 ) | ( n8134 & ~n8146 ) | ( n8145 & ~n8146 ) ;
  assign n8148 = ( n7900 & n8009 ) | ( n7900 & n8147 ) | ( n8009 & n8147 ) ;
  assign n8149 = ( ~n7900 & n8009 ) | ( ~n7900 & n8147 ) | ( n8009 & n8147 ) ;
  assign n8150 = ( n7900 & ~n8148 ) | ( n7900 & n8149 ) | ( ~n8148 & n8149 ) ;
  assign n8151 = ( n7914 & n7999 ) | ( n7914 & n8150 ) | ( n7999 & n8150 ) ;
  assign n8152 = ( ~n7914 & n7999 ) | ( ~n7914 & n8150 ) | ( n7999 & n8150 ) ;
  assign n8153 = ( n7914 & ~n8151 ) | ( n7914 & n8152 ) | ( ~n8151 & n8152 ) ;
  assign n8154 = n1427 & n3591 ;
  assign n8155 = x23 & n8154 ;
  assign n8156 = x101 & n1434 ;
  assign n8157 = x100 & n1431 ;
  assign n8158 = n8156 | n8157 ;
  assign n8159 = x99 & n1531 ;
  assign n8160 = n8158 | n8159 ;
  assign n8161 = ( ~x23 & n8154 ) | ( ~x23 & n8160 ) | ( n8154 & n8160 ) ;
  assign n8162 = x23 & ~n8160 ;
  assign n8163 = ( ~n8155 & n8161 ) | ( ~n8155 & n8162 ) | ( n8161 & n8162 ) ;
  assign n8164 = ( n7916 & ~n8153 ) | ( n7916 & n8163 ) | ( ~n8153 & n8163 ) ;
  assign n8165 = ( n7916 & n8153 ) | ( n7916 & n8163 ) | ( n8153 & n8163 ) ;
  assign n8166 = ( n8153 & n8164 ) | ( n8153 & ~n8165 ) | ( n8164 & ~n8165 ) ;
  assign n8167 = ( n7930 & n7989 ) | ( n7930 & n8166 ) | ( n7989 & n8166 ) ;
  assign n8168 = ( ~n7930 & n7989 ) | ( ~n7930 & n8166 ) | ( n7989 & n8166 ) ;
  assign n8169 = ( n7930 & ~n8167 ) | ( n7930 & n8168 ) | ( ~n8167 & n8168 ) ;
  assign n8170 = n874 & n4523 ;
  assign n8171 = x17 & n8170 ;
  assign n8172 = x107 & n881 ;
  assign n8173 = x106 & n878 ;
  assign n8174 = n8172 | n8173 ;
  assign n8175 = x105 & n959 ;
  assign n8176 = n8174 | n8175 ;
  assign n8177 = ( ~x17 & n8170 ) | ( ~x17 & n8176 ) | ( n8170 & n8176 ) ;
  assign n8178 = x17 & ~n8176 ;
  assign n8179 = ( ~n8171 & n8177 ) | ( ~n8171 & n8178 ) | ( n8177 & n8178 ) ;
  assign n8180 = ( n7932 & ~n8169 ) | ( n7932 & n8179 ) | ( ~n8169 & n8179 ) ;
  assign n8181 = ( n7932 & n8169 ) | ( n7932 & n8179 ) | ( n8169 & n8179 ) ;
  assign n8182 = ( n8169 & n8180 ) | ( n8169 & ~n8181 ) | ( n8180 & ~n8181 ) ;
  assign n8183 = ( n7936 & n7979 ) | ( n7936 & n8182 ) | ( n7979 & n8182 ) ;
  assign n8184 = ( ~n7936 & n7979 ) | ( ~n7936 & n8182 ) | ( n7979 & n8182 ) ;
  assign n8185 = ( n7936 & ~n8183 ) | ( n7936 & n8184 ) | ( ~n8183 & n8184 ) ;
  assign n8186 = n449 & n5774 ;
  assign n8187 = x11 & n8186 ;
  assign n8188 = x113 & n456 ;
  assign n8189 = x112 & n453 ;
  assign n8190 = n8188 | n8189 ;
  assign n8191 = x111 & n536 ;
  assign n8192 = n8190 | n8191 ;
  assign n8193 = ( ~x11 & n8186 ) | ( ~x11 & n8192 ) | ( n8186 & n8192 ) ;
  assign n8194 = x11 & ~n8192 ;
  assign n8195 = ( ~n8187 & n8193 ) | ( ~n8187 & n8194 ) | ( n8193 & n8194 ) ;
  assign n8196 = ( n7939 & ~n8185 ) | ( n7939 & n8195 ) | ( ~n8185 & n8195 ) ;
  assign n8197 = ( n7939 & n8185 ) | ( n7939 & n8195 ) | ( n8185 & n8195 ) ;
  assign n8198 = ( n8185 & n8196 ) | ( n8185 & ~n8197 ) | ( n8196 & ~n8197 ) ;
  assign n8199 = ( n7941 & n7969 ) | ( n7941 & n8198 ) | ( n7969 & n8198 ) ;
  assign n8200 = ( ~n7941 & n7969 ) | ( ~n7941 & n8198 ) | ( n7969 & n8198 ) ;
  assign n8201 = ( n7941 & ~n8199 ) | ( n7941 & n8200 ) | ( ~n8199 & n8200 ) ;
  assign n8202 = ( n7945 & n7959 ) | ( n7945 & n8201 ) | ( n7959 & n8201 ) ;
  assign n8203 = ( ~n7945 & n7959 ) | ( ~n7945 & n8201 ) | ( n7959 & n8201 ) ;
  assign n8204 = ( n7945 & ~n8202 ) | ( n7945 & n8203 ) | ( ~n8202 & n8203 ) ;
  assign n8205 = ( ~x121 & x122 ) | ( ~x121 & n7695 ) | ( x122 & n7695 ) ;
  assign n8206 = ( x121 & x122 ) | ( x121 & n7695 ) | ( x122 & n7695 ) ;
  assign n8207 = ( x121 & n8205 ) | ( x121 & ~n8206 ) | ( n8205 & ~n8206 ) ;
  assign n8208 = x0 & n8207 ;
  assign n8209 = ( x1 & x2 ) | ( x1 & n8208 ) | ( x2 & n8208 ) ;
  assign n8210 = x121 & n172 ;
  assign n8211 = ( ~x120 & n135 ) | ( ~x120 & n174 ) | ( n135 & n174 ) ;
  assign n8212 = n8210 | n8211 ;
  assign n8213 = x122 & n147 ;
  assign n8214 = n8212 | n8213 ;
  assign n8215 = n8209 | n8214 ;
  assign n8216 = n8209 & n8214 ;
  assign n8217 = n8215 & ~n8216 ;
  assign n8218 = ( n7947 & n8204 ) | ( n7947 & n8217 ) | ( n8204 & n8217 ) ;
  assign n8219 = ( ~n7947 & n8204 ) | ( ~n7947 & n8217 ) | ( n8204 & n8217 ) ;
  assign n8220 = ( n7947 & ~n8218 ) | ( n7947 & n8219 ) | ( ~n8218 & n8219 ) ;
  assign n8221 = n301 & n6924 ;
  assign n8222 = x8 & n8221 ;
  assign n8223 = x117 & n309 ;
  assign n8224 = x116 & n306 ;
  assign n8225 = n8223 | n8224 ;
  assign n8226 = x115 & n359 ;
  assign n8227 = n8225 | n8226 ;
  assign n8228 = ( ~x8 & n8221 ) | ( ~x8 & n8227 ) | ( n8221 & n8227 ) ;
  assign n8229 = x8 & ~n8227 ;
  assign n8230 = ( ~n8222 & n8228 ) | ( ~n8222 & n8229 ) | ( n8228 & n8229 ) ;
  assign n8231 = n874 & n4914 ;
  assign n8232 = x17 & n8231 ;
  assign n8233 = x108 & n881 ;
  assign n8234 = x107 & n878 ;
  assign n8235 = n8233 | n8234 ;
  assign n8236 = x106 & n959 ;
  assign n8237 = n8235 | n8236 ;
  assign n8238 = ( ~x17 & n8231 ) | ( ~x17 & n8237 ) | ( n8231 & n8237 ) ;
  assign n8239 = x17 & ~n8237 ;
  assign n8240 = ( ~n8232 & n8238 ) | ( ~n8232 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8241 = n1427 & n3764 ;
  assign n8242 = x23 & n8241 ;
  assign n8243 = x102 & n1434 ;
  assign n8244 = x101 & n1431 ;
  assign n8245 = n8243 | n8244 ;
  assign n8246 = x100 & n1531 ;
  assign n8247 = n8245 | n8246 ;
  assign n8248 = ( ~x23 & n8241 ) | ( ~x23 & n8247 ) | ( n8241 & n8247 ) ;
  assign n8249 = x23 & ~n8247 ;
  assign n8250 = ( ~n8242 & n8248 ) | ( ~n8242 & n8249 ) | ( n8248 & n8249 ) ;
  assign n8251 = n2220 & n2545 ;
  assign n8252 = x32 & n8251 ;
  assign n8253 = x93 & n2552 ;
  assign n8254 = x92 & n2549 ;
  assign n8255 = n8253 | n8254 ;
  assign n8256 = x91 & n2696 ;
  assign n8257 = n8255 | n8256 ;
  assign n8258 = ( ~x32 & n8251 ) | ( ~x32 & n8257 ) | ( n8251 & n8257 ) ;
  assign n8259 = x32 & ~n8257 ;
  assign n8260 = ( ~n8252 & n8258 ) | ( ~n8252 & n8259 ) | ( n8258 & n8259 ) ;
  assign n8261 = ( n7866 & n8039 ) | ( n7866 & n8112 ) | ( n8039 & n8112 ) ;
  assign n8262 = n990 & n4625 ;
  assign n8263 = x44 & n8262 ;
  assign n8264 = x81 & n4791 ;
  assign n8265 = x80 & n4621 ;
  assign n8266 = n8264 | n8265 ;
  assign n8267 = x79 & n4795 ;
  assign n8268 = n8266 | n8267 ;
  assign n8269 = ( ~x44 & n8262 ) | ( ~x44 & n8268 ) | ( n8262 & n8268 ) ;
  assign n8270 = x44 & ~n8268 ;
  assign n8271 = ( ~n8263 & n8269 ) | ( ~n8263 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8272 = n508 & n5858 ;
  assign n8273 = x50 & n8272 ;
  assign n8274 = x75 & n5865 ;
  assign n8275 = x74 & n5862 ;
  assign n8276 = n8274 | n8275 ;
  assign n8277 = x73 & n6092 ;
  assign n8278 = n8276 | n8277 ;
  assign n8279 = ( ~x50 & n8272 ) | ( ~x50 & n8278 ) | ( n8272 & n8278 ) ;
  assign n8280 = x50 & ~n8278 ;
  assign n8281 = ( ~n8273 & n8279 ) | ( ~n8273 & n8280 ) | ( n8279 & n8280 ) ;
  assign n8282 = n240 & n7277 ;
  assign n8283 = x56 & n8282 ;
  assign n8284 = x69 & n7545 ;
  assign n8285 = x68 & n7273 ;
  assign n8286 = n8284 | n8285 ;
  assign n8287 = x67 & n7552 ;
  assign n8288 = n8286 | n8287 ;
  assign n8289 = ( ~x56 & n8282 ) | ( ~x56 & n8288 ) | ( n8282 & n8288 ) ;
  assign n8290 = x56 & ~n8288 ;
  assign n8291 = ( ~n8283 & n8289 ) | ( ~n8283 & n8290 ) | ( n8289 & n8290 ) ;
  assign n8292 = x66 & n8074 ;
  assign n8293 = x65 & n8071 ;
  assign n8294 = n8292 | n8293 ;
  assign n8295 = n226 & n8067 ;
  assign n8296 = n8294 | n8295 ;
  assign n8297 = ~n7821 & n8066 ;
  assign n8298 = ~n8071 & n8297 ;
  assign n8299 = x64 & n8298 ;
  assign n8300 = n8296 | n8299 ;
  assign n8301 = ~x59 & n8300 ;
  assign n8302 = ( x59 & n8077 ) | ( x59 & n8300 ) | ( n8077 & n8300 ) ;
  assign n8303 = n8077 & n8300 ;
  assign n8304 = ( n8301 & n8302 ) | ( n8301 & ~n8303 ) | ( n8302 & ~n8303 ) ;
  assign n8305 = ( n8081 & n8291 ) | ( n8081 & n8304 ) | ( n8291 & n8304 ) ;
  assign n8306 = ( ~n8081 & n8291 ) | ( ~n8081 & n8304 ) | ( n8291 & n8304 ) ;
  assign n8307 = ( n8081 & ~n8305 ) | ( n8081 & n8306 ) | ( ~n8305 & n8306 ) ;
  assign n8308 = n372 & n6546 ;
  assign n8309 = x53 & n8308 ;
  assign n8310 = x72 & n6553 ;
  assign n8311 = x71 & n6550 ;
  assign n8312 = n8310 | n8311 ;
  assign n8313 = x70 & n6787 ;
  assign n8314 = n8312 | n8313 ;
  assign n8315 = ( ~x53 & n8308 ) | ( ~x53 & n8314 ) | ( n8308 & n8314 ) ;
  assign n8316 = x53 & ~n8314 ;
  assign n8317 = ( ~n8309 & n8315 ) | ( ~n8309 & n8316 ) | ( n8315 & n8316 ) ;
  assign n8318 = ( n8094 & ~n8307 ) | ( n8094 & n8317 ) | ( ~n8307 & n8317 ) ;
  assign n8319 = ( n8094 & n8307 ) | ( n8094 & n8317 ) | ( n8307 & n8317 ) ;
  assign n8320 = ( n8307 & n8318 ) | ( n8307 & ~n8319 ) | ( n8318 & ~n8319 ) ;
  assign n8321 = ( n8108 & n8281 ) | ( n8108 & n8320 ) | ( n8281 & n8320 ) ;
  assign n8322 = ( ~n8108 & n8281 ) | ( ~n8108 & n8320 ) | ( n8281 & n8320 ) ;
  assign n8323 = ( n8108 & ~n8321 ) | ( n8108 & n8322 ) | ( ~n8321 & n8322 ) ;
  assign n8324 = n697 & n5223 ;
  assign n8325 = x47 & n8324 ;
  assign n8326 = x78 & n5230 ;
  assign n8327 = x77 & n5227 ;
  assign n8328 = n8326 | n8327 ;
  assign n8329 = x76 & n5434 ;
  assign n8330 = n8328 | n8329 ;
  assign n8331 = ( ~x47 & n8324 ) | ( ~x47 & n8330 ) | ( n8324 & n8330 ) ;
  assign n8332 = x47 & ~n8330 ;
  assign n8333 = ( ~n8325 & n8331 ) | ( ~n8325 & n8332 ) | ( n8331 & n8332 ) ;
  assign n8334 = ( n8110 & ~n8323 ) | ( n8110 & n8333 ) | ( ~n8323 & n8333 ) ;
  assign n8335 = ( n8110 & n8323 ) | ( n8110 & n8333 ) | ( n8323 & n8333 ) ;
  assign n8336 = ( n8323 & n8334 ) | ( n8323 & ~n8335 ) | ( n8334 & ~n8335 ) ;
  assign n8337 = ( n8261 & n8271 ) | ( n8261 & n8336 ) | ( n8271 & n8336 ) ;
  assign n8338 = ( ~n8261 & n8271 ) | ( ~n8261 & n8336 ) | ( n8271 & n8336 ) ;
  assign n8339 = ( n8261 & ~n8337 ) | ( n8261 & n8338 ) | ( ~n8337 & n8338 ) ;
  assign n8340 = ( n7866 & n8039 ) | ( n7866 & ~n8112 ) | ( n8039 & ~n8112 ) ;
  assign n8341 = ( n8112 & ~n8261 ) | ( n8112 & n8340 ) | ( ~n8261 & n8340 ) ;
  assign n8342 = ( n7868 & n8029 ) | ( n7868 & n8341 ) | ( n8029 & n8341 ) ;
  assign n8343 = n1190 & n4020 ;
  assign n8344 = x41 & n8343 ;
  assign n8345 = x84 & n4027 ;
  assign n8346 = x83 & n4024 ;
  assign n8347 = n8345 | n8346 ;
  assign n8348 = x82 & n4223 ;
  assign n8349 = n8347 | n8348 ;
  assign n8350 = ( ~x41 & n8343 ) | ( ~x41 & n8349 ) | ( n8343 & n8349 ) ;
  assign n8351 = x41 & ~n8349 ;
  assign n8352 = ( ~n8344 & n8350 ) | ( ~n8344 & n8351 ) | ( n8350 & n8351 ) ;
  assign n8353 = ( ~n8339 & n8342 ) | ( ~n8339 & n8352 ) | ( n8342 & n8352 ) ;
  assign n8354 = ( n8339 & n8342 ) | ( n8339 & n8352 ) | ( n8342 & n8352 ) ;
  assign n8355 = ( n8339 & n8353 ) | ( n8339 & ~n8354 ) | ( n8353 & ~n8354 ) ;
  assign n8356 = n1494 & n3492 ;
  assign n8357 = x38 & n8356 ;
  assign n8358 = x87 & n3499 ;
  assign n8359 = x86 & n3496 ;
  assign n8360 = n8358 | n8359 ;
  assign n8361 = x85 & n3662 ;
  assign n8362 = n8360 | n8361 ;
  assign n8363 = ( ~x38 & n8356 ) | ( ~x38 & n8362 ) | ( n8356 & n8362 ) ;
  assign n8364 = x38 & ~n8362 ;
  assign n8365 = ( ~n8357 & n8363 ) | ( ~n8357 & n8364 ) | ( n8363 & n8364 ) ;
  assign n8366 = ( n8129 & n8355 ) | ( n8129 & n8365 ) | ( n8355 & n8365 ) ;
  assign n8367 = ( n8129 & ~n8355 ) | ( n8129 & n8365 ) | ( ~n8355 & n8365 ) ;
  assign n8368 = ( n8355 & ~n8366 ) | ( n8355 & n8367 ) | ( ~n8366 & n8367 ) ;
  assign n8369 = n1838 & n2982 ;
  assign n8370 = x35 & n8369 ;
  assign n8371 = x90 & n2989 ;
  assign n8372 = x89 & n2986 ;
  assign n8373 = n8371 | n8372 ;
  assign n8374 = x88 & n3159 ;
  assign n8375 = n8373 | n8374 ;
  assign n8376 = ( ~x35 & n8369 ) | ( ~x35 & n8375 ) | ( n8369 & n8375 ) ;
  assign n8377 = x35 & ~n8375 ;
  assign n8378 = ( ~n8370 & n8376 ) | ( ~n8370 & n8377 ) | ( n8376 & n8377 ) ;
  assign n8379 = ( n8133 & n8368 ) | ( n8133 & n8378 ) | ( n8368 & n8378 ) ;
  assign n8380 = ( ~n8133 & n8368 ) | ( ~n8133 & n8378 ) | ( n8368 & n8378 ) ;
  assign n8381 = ( n8133 & ~n8379 ) | ( n8133 & n8380 ) | ( ~n8379 & n8380 ) ;
  assign n8382 = ( n8146 & n8260 ) | ( n8146 & n8381 ) | ( n8260 & n8381 ) ;
  assign n8383 = ( ~n8146 & n8260 ) | ( ~n8146 & n8381 ) | ( n8260 & n8381 ) ;
  assign n8384 = ( n8146 & ~n8382 ) | ( n8146 & n8383 ) | ( ~n8382 & n8383 ) ;
  assign n8385 = n2137 & n2772 ;
  assign n8386 = x29 & n8385 ;
  assign n8387 = x96 & n2144 ;
  assign n8388 = x95 & n2141 ;
  assign n8389 = n8387 | n8388 ;
  assign n8390 = x94 & n2267 ;
  assign n8391 = n8389 | n8390 ;
  assign n8392 = ( ~x29 & n8385 ) | ( ~x29 & n8391 ) | ( n8385 & n8391 ) ;
  assign n8393 = x29 & ~n8391 ;
  assign n8394 = ( ~n8386 & n8392 ) | ( ~n8386 & n8393 ) | ( n8392 & n8393 ) ;
  assign n8395 = ( ~n8148 & n8384 ) | ( ~n8148 & n8394 ) | ( n8384 & n8394 ) ;
  assign n8396 = ( n8148 & n8384 ) | ( n8148 & n8394 ) | ( n8384 & n8394 ) ;
  assign n8397 = ( n8148 & n8395 ) | ( n8148 & ~n8396 ) | ( n8395 & ~n8396 ) ;
  assign n8398 = x99 & n1762 ;
  assign n8399 = x97 & n1895 ;
  assign n8400 = n8398 | n8399 ;
  assign n8401 = n1755 | n8400 ;
  assign n8402 = ( n3248 & n8400 ) | ( n3248 & n8401 ) | ( n8400 & n8401 ) ;
  assign n8403 = x98 & n1759 ;
  assign n8404 = ( ~x26 & n8402 ) | ( ~x26 & n8403 ) | ( n8402 & n8403 ) ;
  assign n8405 = ( x26 & ~n8402 ) | ( x26 & n8403 ) | ( ~n8402 & n8403 ) ;
  assign n8406 = ~n8403 & n8405 ;
  assign n8407 = n8404 | n8406 ;
  assign n8408 = ( n8151 & ~n8397 ) | ( n8151 & n8407 ) | ( ~n8397 & n8407 ) ;
  assign n8409 = ( n8151 & n8397 ) | ( n8151 & n8407 ) | ( n8397 & n8407 ) ;
  assign n8410 = ( n8397 & n8408 ) | ( n8397 & ~n8409 ) | ( n8408 & ~n8409 ) ;
  assign n8411 = ( n8165 & n8250 ) | ( n8165 & n8410 ) | ( n8250 & n8410 ) ;
  assign n8412 = ( ~n8165 & n8250 ) | ( ~n8165 & n8410 ) | ( n8250 & n8410 ) ;
  assign n8413 = ( n8165 & ~n8411 ) | ( n8165 & n8412 ) | ( ~n8411 & n8412 ) ;
  assign n8414 = n1146 & n4145 ;
  assign n8415 = x20 & n8414 ;
  assign n8416 = x105 & n1153 ;
  assign n8417 = x104 & n1150 ;
  assign n8418 = n8416 | n8417 ;
  assign n8419 = x103 & n1217 ;
  assign n8420 = n8418 | n8419 ;
  assign n8421 = ( ~x20 & n8414 ) | ( ~x20 & n8420 ) | ( n8414 & n8420 ) ;
  assign n8422 = x20 & ~n8420 ;
  assign n8423 = ( ~n8415 & n8421 ) | ( ~n8415 & n8422 ) | ( n8421 & n8422 ) ;
  assign n8424 = ( n8167 & ~n8413 ) | ( n8167 & n8423 ) | ( ~n8413 & n8423 ) ;
  assign n8425 = ( n8167 & n8413 ) | ( n8167 & n8423 ) | ( n8413 & n8423 ) ;
  assign n8426 = ( n8413 & n8424 ) | ( n8413 & ~n8425 ) | ( n8424 & ~n8425 ) ;
  assign n8427 = ( n8181 & n8240 ) | ( n8181 & n8426 ) | ( n8240 & n8426 ) ;
  assign n8428 = ( ~n8181 & n8240 ) | ( ~n8181 & n8426 ) | ( n8240 & n8426 ) ;
  assign n8429 = ( n8181 & ~n8427 ) | ( n8181 & n8428 ) | ( ~n8427 & n8428 ) ;
  assign n8430 = n649 & n5347 ;
  assign n8431 = x14 & n8430 ;
  assign n8432 = x111 & n656 ;
  assign n8433 = x110 & n653 ;
  assign n8434 = n8432 | n8433 ;
  assign n8435 = x109 & n744 ;
  assign n8436 = n8434 | n8435 ;
  assign n8437 = ( ~x14 & n8430 ) | ( ~x14 & n8436 ) | ( n8430 & n8436 ) ;
  assign n8438 = x14 & ~n8436 ;
  assign n8439 = ( ~n8431 & n8437 ) | ( ~n8431 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8440 = ( n8183 & ~n8429 ) | ( n8183 & n8439 ) | ( ~n8429 & n8439 ) ;
  assign n8441 = ( n8183 & n8429 ) | ( n8183 & n8439 ) | ( n8429 & n8439 ) ;
  assign n8442 = ( n8429 & n8440 ) | ( n8429 & ~n8441 ) | ( n8440 & ~n8441 ) ;
  assign n8443 = n449 & n6002 ;
  assign n8444 = x11 & n8443 ;
  assign n8445 = x114 & n456 ;
  assign n8446 = x113 & n453 ;
  assign n8447 = n8445 | n8446 ;
  assign n8448 = x112 & n536 ;
  assign n8449 = n8447 | n8448 ;
  assign n8450 = ( ~x11 & n8443 ) | ( ~x11 & n8449 ) | ( n8443 & n8449 ) ;
  assign n8451 = x11 & ~n8449 ;
  assign n8452 = ( ~n8444 & n8450 ) | ( ~n8444 & n8451 ) | ( n8450 & n8451 ) ;
  assign n8453 = ( n8197 & ~n8442 ) | ( n8197 & n8452 ) | ( ~n8442 & n8452 ) ;
  assign n8454 = ( n8197 & n8442 ) | ( n8197 & n8452 ) | ( n8442 & n8452 ) ;
  assign n8455 = ( n8442 & n8453 ) | ( n8442 & ~n8454 ) | ( n8453 & ~n8454 ) ;
  assign n8456 = ( n8199 & n8230 ) | ( n8199 & n8455 ) | ( n8230 & n8455 ) ;
  assign n8457 = ( ~n8199 & n8230 ) | ( ~n8199 & n8455 ) | ( n8230 & n8455 ) ;
  assign n8458 = ( n8199 & ~n8456 ) | ( n8199 & n8457 ) | ( ~n8456 & n8457 ) ;
  assign n8459 = ( x122 & x123 ) | ( x122 & n8206 ) | ( x123 & n8206 ) ;
  assign n8460 = ( x122 & x123 ) | ( x122 & ~n8206 ) | ( x123 & ~n8206 ) ;
  assign n8461 = ( n8206 & ~n8459 ) | ( n8206 & n8460 ) | ( ~n8459 & n8460 ) ;
  assign n8462 = x0 & n8461 ;
  assign n8463 = ( x1 & x2 ) | ( x1 & n8462 ) | ( x2 & n8462 ) ;
  assign n8464 = x122 & n172 ;
  assign n8465 = ( ~x121 & n135 ) | ( ~x121 & n174 ) | ( n135 & n174 ) ;
  assign n8466 = n8464 | n8465 ;
  assign n8467 = x123 & n147 ;
  assign n8468 = n8466 | n8467 ;
  assign n8469 = n8463 | n8468 ;
  assign n8470 = n8463 & n8468 ;
  assign n8471 = n8469 & ~n8470 ;
  assign n8472 = n206 & n7444 ;
  assign n8473 = x5 & n8472 ;
  assign n8474 = x120 & n205 ;
  assign n8475 = x119 & n201 ;
  assign n8476 = n8474 | n8475 ;
  assign n8477 = x118 & n221 ;
  assign n8478 = n8476 | n8477 ;
  assign n8479 = ( ~x5 & n8472 ) | ( ~x5 & n8478 ) | ( n8472 & n8478 ) ;
  assign n8480 = x5 & ~n8478 ;
  assign n8481 = ( ~n8473 & n8479 ) | ( ~n8473 & n8480 ) | ( n8479 & n8480 ) ;
  assign n8482 = ( n8458 & n8471 ) | ( n8458 & n8481 ) | ( n8471 & n8481 ) ;
  assign n8483 = ( ~n8458 & n8471 ) | ( ~n8458 & n8481 ) | ( n8471 & n8481 ) ;
  assign n8484 = ( n8458 & ~n8482 ) | ( n8458 & n8483 ) | ( ~n8482 & n8483 ) ;
  assign n8485 = ( n8202 & n8218 ) | ( n8202 & n8484 ) | ( n8218 & n8484 ) ;
  assign n8486 = ( n8202 & ~n8218 ) | ( n8202 & n8484 ) | ( ~n8218 & n8484 ) ;
  assign n8487 = ( n8218 & ~n8485 ) | ( n8218 & n8486 ) | ( ~n8485 & n8486 ) ;
  assign n8488 = n301 & n6940 ;
  assign n8489 = x8 & n8488 ;
  assign n8490 = x118 & n309 ;
  assign n8491 = x117 & n306 ;
  assign n8492 = n8490 | n8491 ;
  assign n8493 = x116 & n359 ;
  assign n8494 = n8492 | n8493 ;
  assign n8495 = ( ~x8 & n8488 ) | ( ~x8 & n8494 ) | ( n8488 & n8494 ) ;
  assign n8496 = x8 & ~n8494 ;
  assign n8497 = ( ~n8489 & n8495 ) | ( ~n8489 & n8496 ) | ( n8495 & n8496 ) ;
  assign n8498 = n874 & n4930 ;
  assign n8499 = x17 & n8498 ;
  assign n8500 = x109 & n881 ;
  assign n8501 = x108 & n878 ;
  assign n8502 = n8500 | n8501 ;
  assign n8503 = x107 & n959 ;
  assign n8504 = n8502 | n8503 ;
  assign n8505 = ( ~x17 & n8498 ) | ( ~x17 & n8504 ) | ( n8498 & n8504 ) ;
  assign n8506 = x17 & ~n8504 ;
  assign n8507 = ( ~n8499 & n8505 ) | ( ~n8499 & n8506 ) | ( n8505 & n8506 ) ;
  assign n8508 = n1427 & n3941 ;
  assign n8509 = x23 & n8508 ;
  assign n8510 = x103 & n1434 ;
  assign n8511 = x102 & n1431 ;
  assign n8512 = n8510 | n8511 ;
  assign n8513 = x101 & n1531 ;
  assign n8514 = n8512 | n8513 ;
  assign n8515 = ( ~x23 & n8508 ) | ( ~x23 & n8514 ) | ( n8508 & n8514 ) ;
  assign n8516 = x23 & ~n8514 ;
  assign n8517 = ( ~n8509 & n8515 ) | ( ~n8509 & n8516 ) | ( n8515 & n8516 ) ;
  assign n8518 = n2137 & n2788 ;
  assign n8519 = x29 & n8518 ;
  assign n8520 = x97 & n2144 ;
  assign n8521 = x96 & n2141 ;
  assign n8522 = n8520 | n8521 ;
  assign n8523 = x95 & n2267 ;
  assign n8524 = n8522 | n8523 ;
  assign n8525 = ( ~x29 & n8518 ) | ( ~x29 & n8524 ) | ( n8518 & n8524 ) ;
  assign n8526 = x29 & ~n8524 ;
  assign n8527 = ( ~n8519 & n8525 ) | ( ~n8519 & n8526 ) | ( n8525 & n8526 ) ;
  assign n8528 = n1959 & n2982 ;
  assign n8529 = x35 & n8528 ;
  assign n8530 = x91 & n2989 ;
  assign n8531 = x90 & n2986 ;
  assign n8532 = n8530 | n8531 ;
  assign n8533 = x89 & n3159 ;
  assign n8534 = n8532 | n8533 ;
  assign n8535 = ( ~x35 & n8528 ) | ( ~x35 & n8534 ) | ( n8528 & n8534 ) ;
  assign n8536 = x35 & ~n8534 ;
  assign n8537 = ( ~n8529 & n8535 ) | ( ~n8529 & n8536 ) | ( n8535 & n8536 ) ;
  assign n8538 = n1368 & n4020 ;
  assign n8539 = x41 & n8538 ;
  assign n8540 = x85 & n4027 ;
  assign n8541 = x84 & n4024 ;
  assign n8542 = n8540 | n8541 ;
  assign n8543 = x83 & n4223 ;
  assign n8544 = n8542 | n8543 ;
  assign n8545 = ( ~x41 & n8538 ) | ( ~x41 & n8544 ) | ( n8538 & n8544 ) ;
  assign n8546 = x41 & ~n8544 ;
  assign n8547 = ( ~n8539 & n8545 ) | ( ~n8539 & n8546 ) | ( n8545 & n8546 ) ;
  assign n8548 = n823 & n5223 ;
  assign n8549 = x47 & n8548 ;
  assign n8550 = x79 & n5230 ;
  assign n8551 = x78 & n5227 ;
  assign n8552 = n8550 | n8551 ;
  assign n8553 = x77 & n5434 ;
  assign n8554 = n8552 | n8553 ;
  assign n8555 = ( ~x47 & n8548 ) | ( ~x47 & n8554 ) | ( n8548 & n8554 ) ;
  assign n8556 = x47 & ~n8554 ;
  assign n8557 = ( ~n8549 & n8555 ) | ( ~n8549 & n8556 ) | ( n8555 & n8556 ) ;
  assign n8558 = n388 & n6546 ;
  assign n8559 = x53 & n8558 ;
  assign n8560 = x73 & n6553 ;
  assign n8561 = x72 & n6550 ;
  assign n8562 = n8560 | n8561 ;
  assign n8563 = x71 & n6787 ;
  assign n8564 = n8562 | n8563 ;
  assign n8565 = ( ~x53 & n8558 ) | ( ~x53 & n8564 ) | ( n8558 & n8564 ) ;
  assign n8566 = x53 & ~n8564 ;
  assign n8567 = ( ~n8559 & n8565 ) | ( ~n8559 & n8566 ) | ( n8565 & n8566 ) ;
  assign n8568 = n276 & n7277 ;
  assign n8569 = x56 & n8568 ;
  assign n8570 = x70 & n7545 ;
  assign n8571 = x69 & n7273 ;
  assign n8572 = n8570 | n8571 ;
  assign n8573 = x68 & n7552 ;
  assign n8574 = n8572 | n8573 ;
  assign n8575 = ( ~x56 & n8568 ) | ( ~x56 & n8574 ) | ( n8568 & n8574 ) ;
  assign n8576 = x56 & ~n8574 ;
  assign n8577 = ( ~n8569 & n8575 ) | ( ~n8569 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = n8077 | n8300 ;
  assign n8579 = x59 & n8578 ;
  assign n8580 = x67 & n8074 ;
  assign n8581 = x66 & n8071 ;
  assign n8582 = n8580 | n8581 ;
  assign n8583 = x65 & n8298 ;
  assign n8584 = n8582 | n8583 ;
  assign n8585 = n169 & n8067 ;
  assign n8586 = n8584 | n8585 ;
  assign n8587 = x59 & x60 ;
  assign n8588 = x59 | x60 ;
  assign n8589 = ~n8587 & n8588 ;
  assign n8590 = x64 & n8589 ;
  assign n8591 = ( n8579 & ~n8586 ) | ( n8579 & n8590 ) | ( ~n8586 & n8590 ) ;
  assign n8592 = x59 & ~n8586 ;
  assign n8593 = ( ~n8579 & n8586 ) | ( ~n8579 & n8592 ) | ( n8586 & n8592 ) ;
  assign n8594 = ( n8590 & n8592 ) | ( n8590 & n8593 ) | ( n8592 & n8593 ) ;
  assign n8595 = ( n8591 & n8593 ) | ( n8591 & ~n8594 ) | ( n8593 & ~n8594 ) ;
  assign n8596 = ( n8305 & n8577 ) | ( n8305 & n8595 ) | ( n8577 & n8595 ) ;
  assign n8597 = ( ~n8305 & n8577 ) | ( ~n8305 & n8595 ) | ( n8577 & n8595 ) ;
  assign n8598 = ( n8305 & ~n8596 ) | ( n8305 & n8597 ) | ( ~n8596 & n8597 ) ;
  assign n8599 = ( n8319 & n8567 ) | ( n8319 & n8598 ) | ( n8567 & n8598 ) ;
  assign n8600 = ( ~n8319 & n8567 ) | ( ~n8319 & n8598 ) | ( n8567 & n8598 ) ;
  assign n8601 = ( n8319 & ~n8599 ) | ( n8319 & n8600 ) | ( ~n8599 & n8600 ) ;
  assign n8602 = n565 & n5858 ;
  assign n8603 = x50 & n8602 ;
  assign n8604 = x76 & n5865 ;
  assign n8605 = x75 & n5862 ;
  assign n8606 = n8604 | n8605 ;
  assign n8607 = x74 & n6092 ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = ( ~x50 & n8602 ) | ( ~x50 & n8608 ) | ( n8602 & n8608 ) ;
  assign n8610 = x50 & ~n8608 ;
  assign n8611 = ( ~n8603 & n8609 ) | ( ~n8603 & n8610 ) | ( n8609 & n8610 ) ;
  assign n8612 = ( n8321 & ~n8601 ) | ( n8321 & n8611 ) | ( ~n8601 & n8611 ) ;
  assign n8613 = ( n8321 & n8601 ) | ( n8321 & n8611 ) | ( n8601 & n8611 ) ;
  assign n8614 = ( n8601 & n8612 ) | ( n8601 & ~n8613 ) | ( n8612 & ~n8613 ) ;
  assign n8615 = ( n8335 & n8557 ) | ( n8335 & n8614 ) | ( n8557 & n8614 ) ;
  assign n8616 = ( ~n8335 & n8557 ) | ( ~n8335 & n8614 ) | ( n8557 & n8614 ) ;
  assign n8617 = ( n8335 & ~n8615 ) | ( n8335 & n8616 ) | ( ~n8615 & n8616 ) ;
  assign n8618 = n1006 & n4625 ;
  assign n8619 = x44 & n8618 ;
  assign n8620 = x82 & n4791 ;
  assign n8621 = x81 & n4621 ;
  assign n8622 = n8620 | n8621 ;
  assign n8623 = x80 & n4795 ;
  assign n8624 = n8622 | n8623 ;
  assign n8625 = ( ~x44 & n8618 ) | ( ~x44 & n8624 ) | ( n8618 & n8624 ) ;
  assign n8626 = x44 & ~n8624 ;
  assign n8627 = ( ~n8619 & n8625 ) | ( ~n8619 & n8626 ) | ( n8625 & n8626 ) ;
  assign n8628 = ( n8337 & ~n8617 ) | ( n8337 & n8627 ) | ( ~n8617 & n8627 ) ;
  assign n8629 = ( n8337 & n8617 ) | ( n8337 & n8627 ) | ( n8617 & n8627 ) ;
  assign n8630 = ( n8617 & n8628 ) | ( n8617 & ~n8629 ) | ( n8628 & ~n8629 ) ;
  assign n8631 = ( n8354 & n8547 ) | ( n8354 & n8630 ) | ( n8547 & n8630 ) ;
  assign n8632 = ( ~n8354 & n8547 ) | ( ~n8354 & n8630 ) | ( n8547 & n8630 ) ;
  assign n8633 = ( n8354 & ~n8631 ) | ( n8354 & n8632 ) | ( ~n8631 & n8632 ) ;
  assign n8634 = n1602 & n3492 ;
  assign n8635 = x38 & n8634 ;
  assign n8636 = x88 & n3499 ;
  assign n8637 = x87 & n3496 ;
  assign n8638 = n8636 | n8637 ;
  assign n8639 = x86 & n3662 ;
  assign n8640 = n8638 | n8639 ;
  assign n8641 = ( ~x38 & n8634 ) | ( ~x38 & n8640 ) | ( n8634 & n8640 ) ;
  assign n8642 = x38 & ~n8640 ;
  assign n8643 = ( ~n8635 & n8641 ) | ( ~n8635 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8644 = ( n8366 & ~n8633 ) | ( n8366 & n8643 ) | ( ~n8633 & n8643 ) ;
  assign n8645 = ( n8366 & n8633 ) | ( n8366 & n8643 ) | ( n8633 & n8643 ) ;
  assign n8646 = ( n8633 & n8644 ) | ( n8633 & ~n8645 ) | ( n8644 & ~n8645 ) ;
  assign n8647 = ( ~n8379 & n8537 ) | ( ~n8379 & n8646 ) | ( n8537 & n8646 ) ;
  assign n8648 = ( n8379 & n8537 ) | ( n8379 & n8646 ) | ( n8537 & n8646 ) ;
  assign n8649 = ( n8379 & n8647 ) | ( n8379 & ~n8648 ) | ( n8647 & ~n8648 ) ;
  assign n8650 = n2476 & n2545 ;
  assign n8651 = x32 & n8650 ;
  assign n8652 = x94 & n2552 ;
  assign n8653 = x93 & n2549 ;
  assign n8654 = n8652 | n8653 ;
  assign n8655 = x92 & n2696 ;
  assign n8656 = n8654 | n8655 ;
  assign n8657 = ( ~x32 & n8650 ) | ( ~x32 & n8656 ) | ( n8650 & n8656 ) ;
  assign n8658 = x32 & ~n8656 ;
  assign n8659 = ( ~n8651 & n8657 ) | ( ~n8651 & n8658 ) | ( n8657 & n8658 ) ;
  assign n8660 = ( n8382 & ~n8649 ) | ( n8382 & n8659 ) | ( ~n8649 & n8659 ) ;
  assign n8661 = ( n8382 & n8649 ) | ( n8382 & n8659 ) | ( n8649 & n8659 ) ;
  assign n8662 = ( n8649 & n8660 ) | ( n8649 & ~n8661 ) | ( n8660 & ~n8661 ) ;
  assign n8663 = ( n8396 & n8527 ) | ( n8396 & n8662 ) | ( n8527 & n8662 ) ;
  assign n8664 = ( ~n8396 & n8527 ) | ( ~n8396 & n8662 ) | ( n8527 & n8662 ) ;
  assign n8665 = ( n8396 & ~n8663 ) | ( n8396 & n8664 ) | ( ~n8663 & n8664 ) ;
  assign n8666 = n1755 & n3264 ;
  assign n8667 = x26 & n8666 ;
  assign n8668 = x100 & n1762 ;
  assign n8669 = x99 & n1759 ;
  assign n8670 = n8668 | n8669 ;
  assign n8671 = x98 & n1895 ;
  assign n8672 = n8670 | n8671 ;
  assign n8673 = ( ~x26 & n8666 ) | ( ~x26 & n8672 ) | ( n8666 & n8672 ) ;
  assign n8674 = x26 & ~n8672 ;
  assign n8675 = ( ~n8667 & n8673 ) | ( ~n8667 & n8674 ) | ( n8673 & n8674 ) ;
  assign n8676 = ( n8409 & ~n8665 ) | ( n8409 & n8675 ) | ( ~n8665 & n8675 ) ;
  assign n8677 = ( n8409 & n8665 ) | ( n8409 & n8675 ) | ( n8665 & n8675 ) ;
  assign n8678 = ( n8665 & n8676 ) | ( n8665 & ~n8677 ) | ( n8676 & ~n8677 ) ;
  assign n8679 = ( n8411 & n8517 ) | ( n8411 & n8678 ) | ( n8517 & n8678 ) ;
  assign n8680 = ( ~n8411 & n8517 ) | ( ~n8411 & n8678 ) | ( n8517 & n8678 ) ;
  assign n8681 = ( n8411 & ~n8679 ) | ( n8411 & n8680 ) | ( ~n8679 & n8680 ) ;
  assign n8682 = n1146 & n4331 ;
  assign n8683 = x20 & n8682 ;
  assign n8684 = x106 & n1153 ;
  assign n8685 = x105 & n1150 ;
  assign n8686 = n8684 | n8685 ;
  assign n8687 = x104 & n1217 ;
  assign n8688 = n8686 | n8687 ;
  assign n8689 = ( ~x20 & n8682 ) | ( ~x20 & n8688 ) | ( n8682 & n8688 ) ;
  assign n8690 = x20 & ~n8688 ;
  assign n8691 = ( ~n8683 & n8689 ) | ( ~n8683 & n8690 ) | ( n8689 & n8690 ) ;
  assign n8692 = ( n8425 & ~n8681 ) | ( n8425 & n8691 ) | ( ~n8681 & n8691 ) ;
  assign n8693 = ( n8425 & n8681 ) | ( n8425 & n8691 ) | ( n8681 & n8691 ) ;
  assign n8694 = ( n8681 & n8692 ) | ( n8681 & ~n8693 ) | ( n8692 & ~n8693 ) ;
  assign n8695 = ( n8427 & n8507 ) | ( n8427 & n8694 ) | ( n8507 & n8694 ) ;
  assign n8696 = ( ~n8427 & n8507 ) | ( ~n8427 & n8694 ) | ( n8507 & n8694 ) ;
  assign n8697 = ( n8427 & ~n8695 ) | ( n8427 & n8696 ) | ( ~n8695 & n8696 ) ;
  assign n8698 = n649 & n5558 ;
  assign n8699 = x14 & n8698 ;
  assign n8700 = x112 & n656 ;
  assign n8701 = x111 & n653 ;
  assign n8702 = n8700 | n8701 ;
  assign n8703 = x110 & n744 ;
  assign n8704 = n8702 | n8703 ;
  assign n8705 = ( ~x14 & n8698 ) | ( ~x14 & n8704 ) | ( n8698 & n8704 ) ;
  assign n8706 = x14 & ~n8704 ;
  assign n8707 = ( ~n8699 & n8705 ) | ( ~n8699 & n8706 ) | ( n8705 & n8706 ) ;
  assign n8708 = ( n8441 & ~n8697 ) | ( n8441 & n8707 ) | ( ~n8697 & n8707 ) ;
  assign n8709 = ( n8441 & n8697 ) | ( n8441 & n8707 ) | ( n8697 & n8707 ) ;
  assign n8710 = ( n8697 & n8708 ) | ( n8697 & ~n8709 ) | ( n8708 & ~n8709 ) ;
  assign n8711 = n449 & n6446 ;
  assign n8712 = x11 & n8711 ;
  assign n8713 = x115 & n456 ;
  assign n8714 = x114 & n453 ;
  assign n8715 = n8713 | n8714 ;
  assign n8716 = x113 & n536 ;
  assign n8717 = n8715 | n8716 ;
  assign n8718 = ( ~x11 & n8711 ) | ( ~x11 & n8717 ) | ( n8711 & n8717 ) ;
  assign n8719 = x11 & ~n8717 ;
  assign n8720 = ( ~n8712 & n8718 ) | ( ~n8712 & n8719 ) | ( n8718 & n8719 ) ;
  assign n8721 = ( n8454 & ~n8710 ) | ( n8454 & n8720 ) | ( ~n8710 & n8720 ) ;
  assign n8722 = ( n8454 & n8710 ) | ( n8454 & n8720 ) | ( n8710 & n8720 ) ;
  assign n8723 = ( n8710 & n8721 ) | ( n8710 & ~n8722 ) | ( n8721 & ~n8722 ) ;
  assign n8724 = ( n8456 & n8497 ) | ( n8456 & n8723 ) | ( n8497 & n8723 ) ;
  assign n8725 = ( ~n8456 & n8497 ) | ( ~n8456 & n8723 ) | ( n8497 & n8723 ) ;
  assign n8726 = ( n8456 & ~n8724 ) | ( n8456 & n8725 ) | ( ~n8724 & n8725 ) ;
  assign n8727 = ( x123 & x124 ) | ( x123 & n8459 ) | ( x124 & n8459 ) ;
  assign n8728 = ( x122 & x124 ) | ( x122 & ~n8460 ) | ( x124 & ~n8460 ) ;
  assign n8729 = ( x123 & ~n8727 ) | ( x123 & n8728 ) | ( ~n8727 & n8728 ) ;
  assign n8730 = x0 & n8729 ;
  assign n8731 = ( x1 & x2 ) | ( x1 & n8730 ) | ( x2 & n8730 ) ;
  assign n8732 = x123 & n172 ;
  assign n8733 = x124 | n8732 ;
  assign n8734 = ( n147 & n8732 ) | ( n147 & n8733 ) | ( n8732 & n8733 ) ;
  assign n8735 = ( ~x122 & n135 ) | ( ~x122 & n174 ) | ( n135 & n174 ) ;
  assign n8736 = n8734 | n8735 ;
  assign n8737 = n8731 | n8736 ;
  assign n8738 = n8731 & n8736 ;
  assign n8739 = n8737 & ~n8738 ;
  assign n8740 = n206 & n7696 ;
  assign n8741 = x5 & n8740 ;
  assign n8742 = x121 & n205 ;
  assign n8743 = x120 & n201 ;
  assign n8744 = n8742 | n8743 ;
  assign n8745 = x119 & n221 ;
  assign n8746 = n8744 | n8745 ;
  assign n8747 = ( ~x5 & n8740 ) | ( ~x5 & n8746 ) | ( n8740 & n8746 ) ;
  assign n8748 = x5 & ~n8746 ;
  assign n8749 = ( ~n8741 & n8747 ) | ( ~n8741 & n8748 ) | ( n8747 & n8748 ) ;
  assign n8750 = ( ~n8726 & n8739 ) | ( ~n8726 & n8749 ) | ( n8739 & n8749 ) ;
  assign n8751 = ( n8726 & n8739 ) | ( n8726 & n8749 ) | ( n8739 & n8749 ) ;
  assign n8752 = ( n8726 & n8750 ) | ( n8726 & ~n8751 ) | ( n8750 & ~n8751 ) ;
  assign n8753 = ( n8482 & ~n8485 ) | ( n8482 & n8752 ) | ( ~n8485 & n8752 ) ;
  assign n8754 = ( n8482 & n8485 ) | ( n8482 & n8752 ) | ( n8485 & n8752 ) ;
  assign n8755 = ( n8485 & n8753 ) | ( n8485 & ~n8754 ) | ( n8753 & ~n8754 ) ;
  assign n8756 = n301 & n7181 ;
  assign n8757 = x8 & n8756 ;
  assign n8758 = x119 & n309 ;
  assign n8759 = x118 & n306 ;
  assign n8760 = n8758 | n8759 ;
  assign n8761 = x117 & n359 ;
  assign n8762 = n8760 | n8761 ;
  assign n8763 = ( ~x8 & n8756 ) | ( ~x8 & n8762 ) | ( n8756 & n8762 ) ;
  assign n8764 = x8 & ~n8762 ;
  assign n8765 = ( ~n8757 & n8763 ) | ( ~n8757 & n8764 ) | ( n8763 & n8764 ) ;
  assign n8766 = n874 & n5331 ;
  assign n8767 = x17 & n8766 ;
  assign n8768 = x110 & n881 ;
  assign n8769 = x109 & n878 ;
  assign n8770 = n8768 | n8769 ;
  assign n8771 = x108 & n959 ;
  assign n8772 = n8770 | n8771 ;
  assign n8773 = ( ~x17 & n8766 ) | ( ~x17 & n8772 ) | ( n8766 & n8772 ) ;
  assign n8774 = x17 & ~n8772 ;
  assign n8775 = ( ~n8767 & n8773 ) | ( ~n8767 & n8774 ) | ( n8773 & n8774 ) ;
  assign n8776 = n1146 & n4523 ;
  assign n8777 = x20 & n8776 ;
  assign n8778 = x107 & n1153 ;
  assign n8779 = x106 & n1150 ;
  assign n8780 = n8778 | n8779 ;
  assign n8781 = x105 & n1217 ;
  assign n8782 = n8780 | n8781 ;
  assign n8783 = ( ~x20 & n8776 ) | ( ~x20 & n8782 ) | ( n8776 & n8782 ) ;
  assign n8784 = x20 & ~n8782 ;
  assign n8785 = ( ~n8777 & n8783 ) | ( ~n8777 & n8784 ) | ( n8783 & n8784 ) ;
  assign n8786 = n1755 & n3591 ;
  assign n8787 = x26 & n8786 ;
  assign n8788 = x101 & n1762 ;
  assign n8789 = x100 & n1759 ;
  assign n8790 = n8788 | n8789 ;
  assign n8791 = x99 & n1895 ;
  assign n8792 = n8790 | n8791 ;
  assign n8793 = ( ~x26 & n8786 ) | ( ~x26 & n8792 ) | ( n8786 & n8792 ) ;
  assign n8794 = x26 & ~n8792 ;
  assign n8795 = ( ~n8787 & n8793 ) | ( ~n8787 & n8794 ) | ( n8793 & n8794 ) ;
  assign n8796 = n2492 & n2545 ;
  assign n8797 = x32 & n8796 ;
  assign n8798 = x95 & n2552 ;
  assign n8799 = x94 & n2549 ;
  assign n8800 = n8798 | n8799 ;
  assign n8801 = x93 & n2696 ;
  assign n8802 = n8800 | n8801 ;
  assign n8803 = ( ~x32 & n8796 ) | ( ~x32 & n8802 ) | ( n8796 & n8802 ) ;
  assign n8804 = x32 & ~n8802 ;
  assign n8805 = ( ~n8797 & n8803 ) | ( ~n8797 & n8804 ) | ( n8803 & n8804 ) ;
  assign n8806 = n1384 & n4020 ;
  assign n8807 = x41 & n8806 ;
  assign n8808 = x86 & n4027 ;
  assign n8809 = x85 & n4024 ;
  assign n8810 = n8808 | n8809 ;
  assign n8811 = x84 & n4223 ;
  assign n8812 = n8810 | n8811 ;
  assign n8813 = ( ~x41 & n8806 ) | ( ~x41 & n8812 ) | ( n8806 & n8812 ) ;
  assign n8814 = x41 & ~n8812 ;
  assign n8815 = ( ~n8807 & n8813 ) | ( ~n8807 & n8814 ) | ( n8813 & n8814 ) ;
  assign n8816 = n1093 & n4625 ;
  assign n8817 = x44 & n8816 ;
  assign n8818 = x83 & n4791 ;
  assign n8819 = x82 & n4621 ;
  assign n8820 = n8818 | n8819 ;
  assign n8821 = x81 & n4795 ;
  assign n8822 = n8820 | n8821 ;
  assign n8823 = ( ~x44 & n8816 ) | ( ~x44 & n8822 ) | ( n8816 & n8822 ) ;
  assign n8824 = x44 & ~n8822 ;
  assign n8825 = ( ~n8817 & n8823 ) | ( ~n8817 & n8824 ) | ( n8823 & n8824 ) ;
  assign n8826 = n626 & n5858 ;
  assign n8827 = x50 & n8826 ;
  assign n8828 = x77 & n5865 ;
  assign n8829 = x76 & n5862 ;
  assign n8830 = n8828 | n8829 ;
  assign n8831 = x75 & n6092 ;
  assign n8832 = n8830 | n8831 ;
  assign n8833 = ( ~x50 & n8826 ) | ( ~x50 & n8832 ) | ( n8826 & n8832 ) ;
  assign n8834 = x50 & ~n8832 ;
  assign n8835 = ( ~n8827 & n8833 ) | ( ~n8827 & n8834 ) | ( n8833 & n8834 ) ;
  assign n8836 = n436 & n6546 ;
  assign n8837 = x53 & n8836 ;
  assign n8838 = x74 & n6553 ;
  assign n8839 = x73 & n6550 ;
  assign n8840 = n8838 | n8839 ;
  assign n8841 = x72 & n6787 ;
  assign n8842 = n8840 | n8841 ;
  assign n8843 = ( ~x53 & n8836 ) | ( ~x53 & n8842 ) | ( n8836 & n8842 ) ;
  assign n8844 = x53 & ~n8842 ;
  assign n8845 = ( ~n8837 & n8843 ) | ( ~n8837 & n8844 ) | ( n8843 & n8844 ) ;
  assign n8846 = n193 & n8067 ;
  assign n8847 = x59 & n8846 ;
  assign n8848 = x68 & n8074 ;
  assign n8849 = x67 & n8071 ;
  assign n8850 = n8848 | n8849 ;
  assign n8851 = x66 & n8298 ;
  assign n8852 = n8850 | n8851 ;
  assign n8853 = ( ~x59 & n8846 ) | ( ~x59 & n8852 ) | ( n8846 & n8852 ) ;
  assign n8854 = x59 & ~n8852 ;
  assign n8855 = ( ~n8847 & n8853 ) | ( ~n8847 & n8854 ) | ( n8853 & n8854 ) ;
  assign n8856 = x61 & x62 ;
  assign n8857 = x61 | x62 ;
  assign n8858 = ~n8856 & n8857 ;
  assign n8859 = n8589 & n8858 ;
  assign n8860 = n302 & n8859 ;
  assign n8861 = ~x59 & x61 ;
  assign n8862 = x60 & x61 ;
  assign n8863 = ( n8587 & n8861 ) | ( n8587 & ~n8862 ) | ( n8861 & ~n8862 ) ;
  assign n8864 = x64 & n8863 ;
  assign n8865 = n8860 | n8864 ;
  assign n8866 = ( n8589 & n8856 ) | ( n8589 & ~n8857 ) | ( n8856 & ~n8857 ) ;
  assign n8867 = x65 & n8866 ;
  assign n8868 = n8865 | n8867 ;
  assign n8869 = n8590 | n8868 ;
  assign n8870 = ( x62 & n8590 ) | ( x62 & ~n8868 ) | ( n8590 & ~n8868 ) ;
  assign n8871 = x62 & ~n8868 ;
  assign n8872 = ( n8869 & ~n8870 ) | ( n8869 & n8871 ) | ( ~n8870 & n8871 ) ;
  assign n8873 = ( ~n8594 & n8855 ) | ( ~n8594 & n8872 ) | ( n8855 & n8872 ) ;
  assign n8874 = ( n8594 & n8855 ) | ( n8594 & n8872 ) | ( n8855 & n8872 ) ;
  assign n8875 = ( n8594 & n8873 ) | ( n8594 & ~n8874 ) | ( n8873 & ~n8874 ) ;
  assign n8876 = n322 & n7277 ;
  assign n8877 = x56 & n8876 ;
  assign n8878 = x71 & n7545 ;
  assign n8879 = x70 & n7273 ;
  assign n8880 = n8878 | n8879 ;
  assign n8881 = x69 & n7552 ;
  assign n8882 = n8880 | n8881 ;
  assign n8883 = ( ~x56 & n8876 ) | ( ~x56 & n8882 ) | ( n8876 & n8882 ) ;
  assign n8884 = x56 & ~n8882 ;
  assign n8885 = ( ~n8877 & n8883 ) | ( ~n8877 & n8884 ) | ( n8883 & n8884 ) ;
  assign n8886 = ( n8596 & ~n8875 ) | ( n8596 & n8885 ) | ( ~n8875 & n8885 ) ;
  assign n8887 = ( n8596 & n8875 ) | ( n8596 & n8885 ) | ( n8875 & n8885 ) ;
  assign n8888 = ( n8875 & n8886 ) | ( n8875 & ~n8887 ) | ( n8886 & ~n8887 ) ;
  assign n8889 = ( n8599 & n8845 ) | ( n8599 & n8888 ) | ( n8845 & n8888 ) ;
  assign n8890 = ( ~n8599 & n8845 ) | ( ~n8599 & n8888 ) | ( n8845 & n8888 ) ;
  assign n8891 = ( n8599 & ~n8889 ) | ( n8599 & n8890 ) | ( ~n8889 & n8890 ) ;
  assign n8892 = ( n8613 & n8835 ) | ( n8613 & n8891 ) | ( n8835 & n8891 ) ;
  assign n8893 = ( ~n8613 & n8835 ) | ( ~n8613 & n8891 ) | ( n8835 & n8891 ) ;
  assign n8894 = ( n8613 & ~n8892 ) | ( n8613 & n8893 ) | ( ~n8892 & n8893 ) ;
  assign n8895 = n840 & n5223 ;
  assign n8896 = x47 & n8895 ;
  assign n8897 = x80 & n5230 ;
  assign n8898 = x79 & n5227 ;
  assign n8899 = n8897 | n8898 ;
  assign n8900 = x78 & n5434 ;
  assign n8901 = n8899 | n8900 ;
  assign n8902 = ( ~x47 & n8895 ) | ( ~x47 & n8901 ) | ( n8895 & n8901 ) ;
  assign n8903 = x47 & ~n8901 ;
  assign n8904 = ( ~n8896 & n8902 ) | ( ~n8896 & n8903 ) | ( n8902 & n8903 ) ;
  assign n8905 = ( n8615 & ~n8894 ) | ( n8615 & n8904 ) | ( ~n8894 & n8904 ) ;
  assign n8906 = ( n8615 & n8894 ) | ( n8615 & n8904 ) | ( n8894 & n8904 ) ;
  assign n8907 = ( n8894 & n8905 ) | ( n8894 & ~n8906 ) | ( n8905 & ~n8906 ) ;
  assign n8908 = ( n8629 & n8825 ) | ( n8629 & n8907 ) | ( n8825 & n8907 ) ;
  assign n8909 = ( ~n8629 & n8825 ) | ( ~n8629 & n8907 ) | ( n8825 & n8907 ) ;
  assign n8910 = ( n8629 & ~n8908 ) | ( n8629 & n8909 ) | ( ~n8908 & n8909 ) ;
  assign n8911 = ( n8631 & n8815 ) | ( n8631 & n8910 ) | ( n8815 & n8910 ) ;
  assign n8912 = ( ~n8631 & n8815 ) | ( ~n8631 & n8910 ) | ( n8815 & n8910 ) ;
  assign n8913 = ( n8631 & ~n8911 ) | ( n8631 & n8912 ) | ( ~n8911 & n8912 ) ;
  assign n8914 = n1822 & n3492 ;
  assign n8915 = x38 & n8914 ;
  assign n8916 = x89 & n3499 ;
  assign n8917 = x88 & n3496 ;
  assign n8918 = n8916 | n8917 ;
  assign n8919 = x87 & n3662 ;
  assign n8920 = n8918 | n8919 ;
  assign n8921 = ( ~x38 & n8914 ) | ( ~x38 & n8920 ) | ( n8914 & n8920 ) ;
  assign n8922 = x38 & ~n8920 ;
  assign n8923 = ( ~n8915 & n8921 ) | ( ~n8915 & n8922 ) | ( n8921 & n8922 ) ;
  assign n8924 = ( ~n8645 & n8913 ) | ( ~n8645 & n8923 ) | ( n8913 & n8923 ) ;
  assign n8925 = ( n8645 & n8913 ) | ( n8645 & n8923 ) | ( n8913 & n8923 ) ;
  assign n8926 = ( n8645 & n8924 ) | ( n8645 & ~n8925 ) | ( n8924 & ~n8925 ) ;
  assign n8927 = n2083 & n2982 ;
  assign n8928 = x35 & n8927 ;
  assign n8929 = x92 & n2989 ;
  assign n8930 = x91 & n2986 ;
  assign n8931 = n8929 | n8930 ;
  assign n8932 = x90 & n3159 ;
  assign n8933 = n8931 | n8932 ;
  assign n8934 = ( ~x35 & n8927 ) | ( ~x35 & n8933 ) | ( n8927 & n8933 ) ;
  assign n8935 = x35 & ~n8933 ;
  assign n8936 = ( ~n8928 & n8934 ) | ( ~n8928 & n8935 ) | ( n8934 & n8935 ) ;
  assign n8937 = ( n8648 & ~n8926 ) | ( n8648 & n8936 ) | ( ~n8926 & n8936 ) ;
  assign n8938 = ( n8648 & n8926 ) | ( n8648 & n8936 ) | ( n8926 & n8936 ) ;
  assign n8939 = ( n8926 & n8937 ) | ( n8926 & ~n8938 ) | ( n8937 & ~n8938 ) ;
  assign n8940 = ( n8661 & n8805 ) | ( n8661 & n8939 ) | ( n8805 & n8939 ) ;
  assign n8941 = ( ~n8661 & n8805 ) | ( ~n8661 & n8939 ) | ( n8805 & n8939 ) ;
  assign n8942 = ( n8661 & ~n8940 ) | ( n8661 & n8941 ) | ( ~n8940 & n8941 ) ;
  assign n8943 = n2137 & n2939 ;
  assign n8944 = x29 & n8943 ;
  assign n8945 = x98 & n2144 ;
  assign n8946 = x97 & n2141 ;
  assign n8947 = n8945 | n8946 ;
  assign n8948 = x96 & n2267 ;
  assign n8949 = n8947 | n8948 ;
  assign n8950 = ( ~x29 & n8943 ) | ( ~x29 & n8949 ) | ( n8943 & n8949 ) ;
  assign n8951 = x29 & ~n8949 ;
  assign n8952 = ( ~n8944 & n8950 ) | ( ~n8944 & n8951 ) | ( n8950 & n8951 ) ;
  assign n8953 = ( n8663 & ~n8942 ) | ( n8663 & n8952 ) | ( ~n8942 & n8952 ) ;
  assign n8954 = ( n8663 & n8942 ) | ( n8663 & n8952 ) | ( n8942 & n8952 ) ;
  assign n8955 = ( n8942 & n8953 ) | ( n8942 & ~n8954 ) | ( n8953 & ~n8954 ) ;
  assign n8956 = ( n8677 & n8795 ) | ( n8677 & n8955 ) | ( n8795 & n8955 ) ;
  assign n8957 = ( ~n8677 & n8795 ) | ( ~n8677 & n8955 ) | ( n8795 & n8955 ) ;
  assign n8958 = ( n8677 & ~n8956 ) | ( n8677 & n8957 ) | ( ~n8956 & n8957 ) ;
  assign n8959 = n1427 & n3957 ;
  assign n8960 = x23 & n8959 ;
  assign n8961 = x104 & n1434 ;
  assign n8962 = x103 & n1431 ;
  assign n8963 = n8961 | n8962 ;
  assign n8964 = x102 & n1531 ;
  assign n8965 = n8963 | n8964 ;
  assign n8966 = ( ~x23 & n8959 ) | ( ~x23 & n8965 ) | ( n8959 & n8965 ) ;
  assign n8967 = x23 & ~n8965 ;
  assign n8968 = ( ~n8960 & n8966 ) | ( ~n8960 & n8967 ) | ( n8966 & n8967 ) ;
  assign n8969 = ( n8679 & ~n8958 ) | ( n8679 & n8968 ) | ( ~n8958 & n8968 ) ;
  assign n8970 = ( n8679 & n8958 ) | ( n8679 & n8968 ) | ( n8958 & n8968 ) ;
  assign n8971 = ( n8958 & n8969 ) | ( n8958 & ~n8970 ) | ( n8969 & ~n8970 ) ;
  assign n8972 = ( n8693 & n8785 ) | ( n8693 & n8971 ) | ( n8785 & n8971 ) ;
  assign n8973 = ( ~n8693 & n8785 ) | ( ~n8693 & n8971 ) | ( n8785 & n8971 ) ;
  assign n8974 = ( n8693 & ~n8972 ) | ( n8693 & n8973 ) | ( ~n8972 & n8973 ) ;
  assign n8975 = ( n8695 & n8775 ) | ( n8695 & n8974 ) | ( n8775 & n8974 ) ;
  assign n8976 = ( ~n8695 & n8775 ) | ( ~n8695 & n8974 ) | ( n8775 & n8974 ) ;
  assign n8977 = ( n8695 & ~n8975 ) | ( n8695 & n8976 ) | ( ~n8975 & n8976 ) ;
  assign n8978 = n649 & n5774 ;
  assign n8979 = x14 & n8978 ;
  assign n8980 = x113 & n656 ;
  assign n8981 = x112 & n653 ;
  assign n8982 = n8980 | n8981 ;
  assign n8983 = x111 & n744 ;
  assign n8984 = n8982 | n8983 ;
  assign n8985 = ( ~x14 & n8978 ) | ( ~x14 & n8984 ) | ( n8978 & n8984 ) ;
  assign n8986 = x14 & ~n8984 ;
  assign n8987 = ( ~n8979 & n8985 ) | ( ~n8979 & n8986 ) | ( n8985 & n8986 ) ;
  assign n8988 = ( n8709 & ~n8977 ) | ( n8709 & n8987 ) | ( ~n8977 & n8987 ) ;
  assign n8989 = ( n8709 & n8977 ) | ( n8709 & n8987 ) | ( n8977 & n8987 ) ;
  assign n8990 = ( n8977 & n8988 ) | ( n8977 & ~n8989 ) | ( n8988 & ~n8989 ) ;
  assign n8991 = n449 & n6462 ;
  assign n8992 = x11 & n8991 ;
  assign n8993 = x116 & n456 ;
  assign n8994 = x115 & n453 ;
  assign n8995 = n8993 | n8994 ;
  assign n8996 = x114 & n536 ;
  assign n8997 = n8995 | n8996 ;
  assign n8998 = ( ~x11 & n8991 ) | ( ~x11 & n8997 ) | ( n8991 & n8997 ) ;
  assign n8999 = x11 & ~n8997 ;
  assign n9000 = ( ~n8992 & n8998 ) | ( ~n8992 & n8999 ) | ( n8998 & n8999 ) ;
  assign n9001 = ( n8722 & ~n8990 ) | ( n8722 & n9000 ) | ( ~n8990 & n9000 ) ;
  assign n9002 = ( n8722 & n8990 ) | ( n8722 & n9000 ) | ( n8990 & n9000 ) ;
  assign n9003 = ( n8990 & n9001 ) | ( n8990 & ~n9002 ) | ( n9001 & ~n9002 ) ;
  assign n9004 = ( n8724 & n8765 ) | ( n8724 & n9003 ) | ( n8765 & n9003 ) ;
  assign n9005 = ( ~n8724 & n8765 ) | ( ~n8724 & n9003 ) | ( n8765 & n9003 ) ;
  assign n9006 = ( n8724 & ~n9004 ) | ( n8724 & n9005 ) | ( ~n9004 & n9005 ) ;
  assign n9007 = ( ~x124 & x125 ) | ( ~x124 & n8727 ) | ( x125 & n8727 ) ;
  assign n9008 = ( x124 & x125 ) | ( x124 & n8727 ) | ( x125 & n8727 ) ;
  assign n9009 = ( x124 & n9007 ) | ( x124 & ~n9008 ) | ( n9007 & ~n9008 ) ;
  assign n9010 = x0 & n9009 ;
  assign n9011 = ( x1 & x2 ) | ( x1 & n9010 ) | ( x2 & n9010 ) ;
  assign n9012 = x124 & n172 ;
  assign n9013 = ( ~x123 & n135 ) | ( ~x123 & n174 ) | ( n135 & n174 ) ;
  assign n9014 = n9012 | n9013 ;
  assign n9015 = x125 & n147 ;
  assign n9016 = n9014 | n9015 ;
  assign n9017 = n9011 | n9016 ;
  assign n9018 = n9011 & n9016 ;
  assign n9019 = n9017 & ~n9018 ;
  assign n9020 = n206 & n8207 ;
  assign n9021 = x5 & n9020 ;
  assign n9022 = x122 & n205 ;
  assign n9023 = x121 & n201 ;
  assign n9024 = n9022 | n9023 ;
  assign n9025 = x120 & n221 ;
  assign n9026 = n9024 | n9025 ;
  assign n9027 = ( ~x5 & n9020 ) | ( ~x5 & n9026 ) | ( n9020 & n9026 ) ;
  assign n9028 = x5 & ~n9026 ;
  assign n9029 = ( ~n9021 & n9027 ) | ( ~n9021 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9030 = ( ~n9006 & n9019 ) | ( ~n9006 & n9029 ) | ( n9019 & n9029 ) ;
  assign n9031 = ( n9006 & n9019 ) | ( n9006 & n9029 ) | ( n9019 & n9029 ) ;
  assign n9032 = ( n9006 & n9030 ) | ( n9006 & ~n9031 ) | ( n9030 & ~n9031 ) ;
  assign n9033 = ( n8751 & n8754 ) | ( n8751 & n9032 ) | ( n8754 & n9032 ) ;
  assign n9034 = ( n8751 & ~n8754 ) | ( n8751 & n9032 ) | ( ~n8754 & n9032 ) ;
  assign n9035 = ( n8754 & ~n9033 ) | ( n8754 & n9034 ) | ( ~n9033 & n9034 ) ;
  assign n9036 = ( x125 & x126 ) | ( x125 & n9008 ) | ( x126 & n9008 ) ;
  assign n9037 = ( x125 & x126 ) | ( x125 & ~n9008 ) | ( x126 & ~n9008 ) ;
  assign n9038 = ( n9008 & ~n9036 ) | ( n9008 & n9037 ) | ( ~n9036 & n9037 ) ;
  assign n9039 = x0 & n9038 ;
  assign n9040 = ( x1 & x2 ) | ( x1 & n9039 ) | ( x2 & n9039 ) ;
  assign n9041 = x125 & n172 ;
  assign n9042 = ( ~x124 & n135 ) | ( ~x124 & n174 ) | ( n135 & n174 ) ;
  assign n9043 = n9041 | n9042 ;
  assign n9044 = x126 & n147 ;
  assign n9045 = n9043 | n9044 ;
  assign n9046 = n9040 | n9045 ;
  assign n9047 = n9040 & n9045 ;
  assign n9048 = n9046 & ~n9047 ;
  assign n9049 = n649 & n6002 ;
  assign n9050 = x14 & n9049 ;
  assign n9051 = x114 & n656 ;
  assign n9052 = x113 & n653 ;
  assign n9053 = n9051 | n9052 ;
  assign n9054 = x112 & n744 ;
  assign n9055 = n9053 | n9054 ;
  assign n9056 = ( ~x14 & n9049 ) | ( ~x14 & n9055 ) | ( n9049 & n9055 ) ;
  assign n9057 = x14 & ~n9055 ;
  assign n9058 = ( ~n9050 & n9056 ) | ( ~n9050 & n9057 ) | ( n9056 & n9057 ) ;
  assign n9059 = n1146 & n4914 ;
  assign n9060 = x20 & n9059 ;
  assign n9061 = x108 & n1153 ;
  assign n9062 = x107 & n1150 ;
  assign n9063 = n9061 | n9062 ;
  assign n9064 = x106 & n1217 ;
  assign n9065 = n9063 | n9064 ;
  assign n9066 = ( ~x20 & n9059 ) | ( ~x20 & n9065 ) | ( n9059 & n9065 ) ;
  assign n9067 = x20 & ~n9065 ;
  assign n9068 = ( ~n9060 & n9066 ) | ( ~n9060 & n9067 ) | ( n9066 & n9067 ) ;
  assign n9069 = n1755 & n3764 ;
  assign n9070 = x26 & n9069 ;
  assign n9071 = x102 & n1762 ;
  assign n9072 = x101 & n1759 ;
  assign n9073 = n9071 | n9072 ;
  assign n9074 = x100 & n1895 ;
  assign n9075 = n9073 | n9074 ;
  assign n9076 = ( ~x26 & n9069 ) | ( ~x26 & n9075 ) | ( n9069 & n9075 ) ;
  assign n9077 = x26 & ~n9075 ;
  assign n9078 = ( ~n9070 & n9076 ) | ( ~n9070 & n9077 ) | ( n9076 & n9077 ) ;
  assign n9079 = n2545 & n2772 ;
  assign n9080 = x32 & n9079 ;
  assign n9081 = x96 & n2552 ;
  assign n9082 = x95 & n2549 ;
  assign n9083 = n9081 | n9082 ;
  assign n9084 = x94 & n2696 ;
  assign n9085 = n9083 | n9084 ;
  assign n9086 = ( ~x32 & n9079 ) | ( ~x32 & n9085 ) | ( n9079 & n9085 ) ;
  assign n9087 = x32 & ~n9085 ;
  assign n9088 = ( ~n9080 & n9086 ) | ( ~n9080 & n9087 ) | ( n9086 & n9087 ) ;
  assign n9089 = n1838 & n3492 ;
  assign n9090 = x38 & n9089 ;
  assign n9091 = x90 & n3499 ;
  assign n9092 = x89 & n3496 ;
  assign n9093 = n9091 | n9092 ;
  assign n9094 = x88 & n3662 ;
  assign n9095 = n9093 | n9094 ;
  assign n9096 = ( ~x38 & n9089 ) | ( ~x38 & n9095 ) | ( n9089 & n9095 ) ;
  assign n9097 = x38 & ~n9095 ;
  assign n9098 = ( ~n9090 & n9096 ) | ( ~n9090 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9099 = n990 & n5223 ;
  assign n9100 = x47 & n9099 ;
  assign n9101 = x81 & n5230 ;
  assign n9102 = x80 & n5227 ;
  assign n9103 = n9101 | n9102 ;
  assign n9104 = x79 & n5434 ;
  assign n9105 = n9103 | n9104 ;
  assign n9106 = ( ~x47 & n9099 ) | ( ~x47 & n9105 ) | ( n9099 & n9105 ) ;
  assign n9107 = x47 & ~n9105 ;
  assign n9108 = ( ~n9100 & n9106 ) | ( ~n9100 & n9107 ) | ( n9106 & n9107 ) ;
  assign n9109 = n508 & n6546 ;
  assign n9110 = x53 & n9109 ;
  assign n9111 = x75 & n6553 ;
  assign n9112 = x74 & n6550 ;
  assign n9113 = n9111 | n9112 ;
  assign n9114 = x73 & n6787 ;
  assign n9115 = n9113 | n9114 ;
  assign n9116 = ( ~x53 & n9109 ) | ( ~x53 & n9115 ) | ( n9109 & n9115 ) ;
  assign n9117 = x53 & ~n9115 ;
  assign n9118 = ( ~n9110 & n9116 ) | ( ~n9110 & n9117 ) | ( n9116 & n9117 ) ;
  assign n9119 = x66 & n8866 ;
  assign n9120 = x65 & n8863 ;
  assign n9121 = n9119 | n9120 ;
  assign n9122 = n226 & n8859 ;
  assign n9123 = n9121 | n9122 ;
  assign n9124 = ~n8589 & n8858 ;
  assign n9125 = ~n8863 & n9124 ;
  assign n9126 = x64 & n9125 ;
  assign n9127 = n9123 | n9126 ;
  assign n9128 = ~x62 & n9127 ;
  assign n9129 = ( x62 & n8869 ) | ( x62 & n9127 ) | ( n8869 & n9127 ) ;
  assign n9130 = n8869 & n9127 ;
  assign n9131 = ( n9128 & n9129 ) | ( n9128 & ~n9130 ) | ( n9129 & ~n9130 ) ;
  assign n9132 = n240 & n8067 ;
  assign n9133 = x59 & n9132 ;
  assign n9134 = x69 & n8074 ;
  assign n9135 = x68 & n8071 ;
  assign n9136 = n9134 | n9135 ;
  assign n9137 = x67 & n8298 ;
  assign n9138 = n9136 | n9137 ;
  assign n9139 = ( ~x59 & n9132 ) | ( ~x59 & n9138 ) | ( n9132 & n9138 ) ;
  assign n9140 = x59 & ~n9138 ;
  assign n9141 = ( ~n9133 & n9139 ) | ( ~n9133 & n9140 ) | ( n9139 & n9140 ) ;
  assign n9142 = ( n8874 & n9131 ) | ( n8874 & n9141 ) | ( n9131 & n9141 ) ;
  assign n9143 = ( ~n8874 & n9131 ) | ( ~n8874 & n9141 ) | ( n9131 & n9141 ) ;
  assign n9144 = ( n8874 & ~n9142 ) | ( n8874 & n9143 ) | ( ~n9142 & n9143 ) ;
  assign n9145 = n372 & n7277 ;
  assign n9146 = x56 & n9145 ;
  assign n9147 = x72 & n7545 ;
  assign n9148 = x71 & n7273 ;
  assign n9149 = n9147 | n9148 ;
  assign n9150 = x70 & n7552 ;
  assign n9151 = n9149 | n9150 ;
  assign n9152 = ( ~x56 & n9145 ) | ( ~x56 & n9151 ) | ( n9145 & n9151 ) ;
  assign n9153 = x56 & ~n9151 ;
  assign n9154 = ( ~n9146 & n9152 ) | ( ~n9146 & n9153 ) | ( n9152 & n9153 ) ;
  assign n9155 = ( n8887 & ~n9144 ) | ( n8887 & n9154 ) | ( ~n9144 & n9154 ) ;
  assign n9156 = ( n8887 & n9144 ) | ( n8887 & n9154 ) | ( n9144 & n9154 ) ;
  assign n9157 = ( n9144 & n9155 ) | ( n9144 & ~n9156 ) | ( n9155 & ~n9156 ) ;
  assign n9158 = ( n8889 & n9118 ) | ( n8889 & n9157 ) | ( n9118 & n9157 ) ;
  assign n9159 = ( ~n8889 & n9118 ) | ( ~n8889 & n9157 ) | ( n9118 & n9157 ) ;
  assign n9160 = ( n8889 & ~n9158 ) | ( n8889 & n9159 ) | ( ~n9158 & n9159 ) ;
  assign n9161 = n697 & n5858 ;
  assign n9162 = x50 & n9161 ;
  assign n9163 = x78 & n5865 ;
  assign n9164 = x77 & n5862 ;
  assign n9165 = n9163 | n9164 ;
  assign n9166 = x76 & n6092 ;
  assign n9167 = n9165 | n9166 ;
  assign n9168 = ( ~x50 & n9161 ) | ( ~x50 & n9167 ) | ( n9161 & n9167 ) ;
  assign n9169 = x50 & ~n9167 ;
  assign n9170 = ( ~n9162 & n9168 ) | ( ~n9162 & n9169 ) | ( n9168 & n9169 ) ;
  assign n9171 = ( n8892 & ~n9160 ) | ( n8892 & n9170 ) | ( ~n9160 & n9170 ) ;
  assign n9172 = ( n8892 & n9160 ) | ( n8892 & n9170 ) | ( n9160 & n9170 ) ;
  assign n9173 = ( n9160 & n9171 ) | ( n9160 & ~n9172 ) | ( n9171 & ~n9172 ) ;
  assign n9174 = ( n8906 & n9108 ) | ( n8906 & n9173 ) | ( n9108 & n9173 ) ;
  assign n9175 = ( ~n8906 & n9108 ) | ( ~n8906 & n9173 ) | ( n9108 & n9173 ) ;
  assign n9176 = ( n8906 & ~n9174 ) | ( n8906 & n9175 ) | ( ~n9174 & n9175 ) ;
  assign n9177 = n1190 & n4625 ;
  assign n9178 = x44 & n9177 ;
  assign n9179 = x84 & n4791 ;
  assign n9180 = x83 & n4621 ;
  assign n9181 = n9179 | n9180 ;
  assign n9182 = x82 & n4795 ;
  assign n9183 = n9181 | n9182 ;
  assign n9184 = ( ~x44 & n9177 ) | ( ~x44 & n9183 ) | ( n9177 & n9183 ) ;
  assign n9185 = x44 & ~n9183 ;
  assign n9186 = ( ~n9178 & n9184 ) | ( ~n9178 & n9185 ) | ( n9184 & n9185 ) ;
  assign n9187 = ( n8908 & n9176 ) | ( n8908 & n9186 ) | ( n9176 & n9186 ) ;
  assign n9188 = ( ~n8908 & n9176 ) | ( ~n8908 & n9186 ) | ( n9176 & n9186 ) ;
  assign n9189 = ( n8908 & ~n9187 ) | ( n8908 & n9188 ) | ( ~n9187 & n9188 ) ;
  assign n9190 = n1494 & n4020 ;
  assign n9191 = x41 & n9190 ;
  assign n9192 = x87 & n4027 ;
  assign n9193 = x86 & n4024 ;
  assign n9194 = n9192 | n9193 ;
  assign n9195 = x85 & n4223 ;
  assign n9196 = n9194 | n9195 ;
  assign n9197 = ( ~x41 & n9190 ) | ( ~x41 & n9196 ) | ( n9190 & n9196 ) ;
  assign n9198 = x41 & ~n9196 ;
  assign n9199 = ( ~n9191 & n9197 ) | ( ~n9191 & n9198 ) | ( n9197 & n9198 ) ;
  assign n9200 = ( n8911 & ~n9189 ) | ( n8911 & n9199 ) | ( ~n9189 & n9199 ) ;
  assign n9201 = ( n8911 & n9189 ) | ( n8911 & n9199 ) | ( n9189 & n9199 ) ;
  assign n9202 = ( n9189 & n9200 ) | ( n9189 & ~n9201 ) | ( n9200 & ~n9201 ) ;
  assign n9203 = ( n8925 & n9098 ) | ( n8925 & n9202 ) | ( n9098 & n9202 ) ;
  assign n9204 = ( ~n8925 & n9098 ) | ( ~n8925 & n9202 ) | ( n9098 & n9202 ) ;
  assign n9205 = ( n8925 & ~n9203 ) | ( n8925 & n9204 ) | ( ~n9203 & n9204 ) ;
  assign n9206 = n2220 & n2982 ;
  assign n9207 = x35 & n9206 ;
  assign n9208 = x93 & n2989 ;
  assign n9209 = x92 & n2986 ;
  assign n9210 = n9208 | n9209 ;
  assign n9211 = x91 & n3159 ;
  assign n9212 = n9210 | n9211 ;
  assign n9213 = ( ~x35 & n9206 ) | ( ~x35 & n9212 ) | ( n9206 & n9212 ) ;
  assign n9214 = x35 & ~n9212 ;
  assign n9215 = ( ~n9207 & n9213 ) | ( ~n9207 & n9214 ) | ( n9213 & n9214 ) ;
  assign n9216 = ( n8938 & ~n9205 ) | ( n8938 & n9215 ) | ( ~n9205 & n9215 ) ;
  assign n9217 = ( n8938 & n9205 ) | ( n8938 & n9215 ) | ( n9205 & n9215 ) ;
  assign n9218 = ( n9205 & n9216 ) | ( n9205 & ~n9217 ) | ( n9216 & ~n9217 ) ;
  assign n9219 = ( n8940 & n9088 ) | ( n8940 & n9218 ) | ( n9088 & n9218 ) ;
  assign n9220 = ( ~n8940 & n9088 ) | ( ~n8940 & n9218 ) | ( n9088 & n9218 ) ;
  assign n9221 = ( n8940 & ~n9219 ) | ( n8940 & n9220 ) | ( ~n9219 & n9220 ) ;
  assign n9222 = n2137 & n3248 ;
  assign n9223 = x29 & n9222 ;
  assign n9224 = x99 & n2144 ;
  assign n9225 = x98 & n2141 ;
  assign n9226 = n9224 | n9225 ;
  assign n9227 = x97 & n2267 ;
  assign n9228 = n9226 | n9227 ;
  assign n9229 = ( ~x29 & n9222 ) | ( ~x29 & n9228 ) | ( n9222 & n9228 ) ;
  assign n9230 = x29 & ~n9228 ;
  assign n9231 = ( ~n9223 & n9229 ) | ( ~n9223 & n9230 ) | ( n9229 & n9230 ) ;
  assign n9232 = ( n8954 & ~n9221 ) | ( n8954 & n9231 ) | ( ~n9221 & n9231 ) ;
  assign n9233 = ( n8954 & n9221 ) | ( n8954 & n9231 ) | ( n9221 & n9231 ) ;
  assign n9234 = ( n9221 & n9232 ) | ( n9221 & ~n9233 ) | ( n9232 & ~n9233 ) ;
  assign n9235 = ( n8956 & n9078 ) | ( n8956 & n9234 ) | ( n9078 & n9234 ) ;
  assign n9236 = ( ~n8956 & n9078 ) | ( ~n8956 & n9234 ) | ( n9078 & n9234 ) ;
  assign n9237 = ( n8956 & ~n9235 ) | ( n8956 & n9236 ) | ( ~n9235 & n9236 ) ;
  assign n9238 = n1427 & n4145 ;
  assign n9239 = x23 & n9238 ;
  assign n9240 = x105 & n1434 ;
  assign n9241 = x104 & n1431 ;
  assign n9242 = n9240 | n9241 ;
  assign n9243 = x103 & n1531 ;
  assign n9244 = n9242 | n9243 ;
  assign n9245 = ( ~x23 & n9238 ) | ( ~x23 & n9244 ) | ( n9238 & n9244 ) ;
  assign n9246 = x23 & ~n9244 ;
  assign n9247 = ( ~n9239 & n9245 ) | ( ~n9239 & n9246 ) | ( n9245 & n9246 ) ;
  assign n9248 = ( n8970 & ~n9237 ) | ( n8970 & n9247 ) | ( ~n9237 & n9247 ) ;
  assign n9249 = ( n8970 & n9237 ) | ( n8970 & n9247 ) | ( n9237 & n9247 ) ;
  assign n9250 = ( n9237 & n9248 ) | ( n9237 & ~n9249 ) | ( n9248 & ~n9249 ) ;
  assign n9251 = ( n8972 & n9068 ) | ( n8972 & n9250 ) | ( n9068 & n9250 ) ;
  assign n9252 = ( ~n8972 & n9068 ) | ( ~n8972 & n9250 ) | ( n9068 & n9250 ) ;
  assign n9253 = ( n8972 & ~n9251 ) | ( n8972 & n9252 ) | ( ~n9251 & n9252 ) ;
  assign n9254 = n874 & n5347 ;
  assign n9255 = x17 & n9254 ;
  assign n9256 = x111 & n881 ;
  assign n9257 = x110 & n878 ;
  assign n9258 = n9256 | n9257 ;
  assign n9259 = x109 & n959 ;
  assign n9260 = n9258 | n9259 ;
  assign n9261 = ( ~x17 & n9254 ) | ( ~x17 & n9260 ) | ( n9254 & n9260 ) ;
  assign n9262 = x17 & ~n9260 ;
  assign n9263 = ( ~n9255 & n9261 ) | ( ~n9255 & n9262 ) | ( n9261 & n9262 ) ;
  assign n9264 = ( n8975 & ~n9253 ) | ( n8975 & n9263 ) | ( ~n9253 & n9263 ) ;
  assign n9265 = ( n8975 & n9253 ) | ( n8975 & n9263 ) | ( n9253 & n9263 ) ;
  assign n9266 = ( n9253 & n9264 ) | ( n9253 & ~n9265 ) | ( n9264 & ~n9265 ) ;
  assign n9267 = ( n8989 & n9058 ) | ( n8989 & n9266 ) | ( n9058 & n9266 ) ;
  assign n9268 = ( ~n8989 & n9058 ) | ( ~n8989 & n9266 ) | ( n9058 & n9266 ) ;
  assign n9269 = ( n8989 & ~n9267 ) | ( n8989 & n9268 ) | ( ~n9267 & n9268 ) ;
  assign n9270 = n449 & n6924 ;
  assign n9271 = x11 & n9270 ;
  assign n9272 = x117 & n456 ;
  assign n9273 = x116 & n453 ;
  assign n9274 = n9272 | n9273 ;
  assign n9275 = x115 & n536 ;
  assign n9276 = n9274 | n9275 ;
  assign n9277 = ( ~x11 & n9270 ) | ( ~x11 & n9276 ) | ( n9270 & n9276 ) ;
  assign n9278 = x11 & ~n9276 ;
  assign n9279 = ( ~n9271 & n9277 ) | ( ~n9271 & n9278 ) | ( n9277 & n9278 ) ;
  assign n9280 = ( n9002 & ~n9269 ) | ( n9002 & n9279 ) | ( ~n9269 & n9279 ) ;
  assign n9281 = ( n9002 & n9269 ) | ( n9002 & n9279 ) | ( n9269 & n9279 ) ;
  assign n9282 = ( n9269 & n9280 ) | ( n9269 & ~n9281 ) | ( n9280 & ~n9281 ) ;
  assign n9283 = n206 & n8461 ;
  assign n9284 = x5 & n9283 ;
  assign n9285 = x123 & n205 ;
  assign n9286 = x122 & n201 ;
  assign n9287 = n9285 | n9286 ;
  assign n9288 = x121 & n221 ;
  assign n9289 = n9287 | n9288 ;
  assign n9290 = ( ~x5 & n9283 ) | ( ~x5 & n9289 ) | ( n9283 & n9289 ) ;
  assign n9291 = x5 & ~n9289 ;
  assign n9292 = ( ~n9284 & n9290 ) | ( ~n9284 & n9291 ) | ( n9290 & n9291 ) ;
  assign n9293 = n301 & n7444 ;
  assign n9294 = x8 & n9293 ;
  assign n9295 = x120 & n309 ;
  assign n9296 = x119 & n306 ;
  assign n9297 = n9295 | n9296 ;
  assign n9298 = x118 & n359 ;
  assign n9299 = n9297 | n9298 ;
  assign n9300 = ( ~x8 & n9293 ) | ( ~x8 & n9299 ) | ( n9293 & n9299 ) ;
  assign n9301 = x8 & ~n9299 ;
  assign n9302 = ( ~n9294 & n9300 ) | ( ~n9294 & n9301 ) | ( n9300 & n9301 ) ;
  assign n9303 = ( n9282 & n9292 ) | ( n9282 & n9302 ) | ( n9292 & n9302 ) ;
  assign n9304 = ( ~n9282 & n9292 ) | ( ~n9282 & n9302 ) | ( n9292 & n9302 ) ;
  assign n9305 = ( n9282 & ~n9303 ) | ( n9282 & n9304 ) | ( ~n9303 & n9304 ) ;
  assign n9306 = ( n9004 & ~n9048 ) | ( n9004 & n9305 ) | ( ~n9048 & n9305 ) ;
  assign n9307 = ( n9004 & n9048 ) | ( n9004 & n9305 ) | ( n9048 & n9305 ) ;
  assign n9308 = ( n9048 & n9306 ) | ( n9048 & ~n9307 ) | ( n9306 & ~n9307 ) ;
  assign n9309 = ( n9031 & ~n9033 ) | ( n9031 & n9308 ) | ( ~n9033 & n9308 ) ;
  assign n9310 = ( n9031 & n9033 ) | ( n9031 & n9308 ) | ( n9033 & n9308 ) ;
  assign n9311 = ( n9033 & n9309 ) | ( n9033 & ~n9310 ) | ( n9309 & ~n9310 ) ;
  assign n9312 = n1146 & n4930 ;
  assign n9313 = x20 & n9312 ;
  assign n9314 = x109 & n1153 ;
  assign n9315 = x108 & n1150 ;
  assign n9316 = n9314 | n9315 ;
  assign n9317 = x107 & n1217 ;
  assign n9318 = n9316 | n9317 ;
  assign n9319 = ( ~x20 & n9312 ) | ( ~x20 & n9318 ) | ( n9312 & n9318 ) ;
  assign n9320 = x20 & ~n9318 ;
  assign n9321 = ( ~n9313 & n9319 ) | ( ~n9313 & n9320 ) | ( n9319 & n9320 ) ;
  assign n9322 = n1427 & n4331 ;
  assign n9323 = x23 & n9322 ;
  assign n9324 = x106 & n1434 ;
  assign n9325 = x105 & n1431 ;
  assign n9326 = n9324 | n9325 ;
  assign n9327 = x104 & n1531 ;
  assign n9328 = n9326 | n9327 ;
  assign n9329 = ( ~x23 & n9322 ) | ( ~x23 & n9328 ) | ( n9322 & n9328 ) ;
  assign n9330 = x23 & ~n9328 ;
  assign n9331 = ( ~n9323 & n9329 ) | ( ~n9323 & n9330 ) | ( n9329 & n9330 ) ;
  assign n9332 = ~n9321 & n9331 ;
  assign n9333 = n9321 & ~n9331 ;
  assign n9334 = n9332 | n9333 ;
  assign n9335 = n1755 & n3941 ;
  assign n9336 = x26 & n9335 ;
  assign n9337 = x103 & n1762 ;
  assign n9338 = x102 & n1759 ;
  assign n9339 = n9337 | n9338 ;
  assign n9340 = x101 & n1895 ;
  assign n9341 = n9339 | n9340 ;
  assign n9342 = ( ~x26 & n9335 ) | ( ~x26 & n9341 ) | ( n9335 & n9341 ) ;
  assign n9343 = x26 & ~n9341 ;
  assign n9344 = ( ~n9336 & n9342 ) | ( ~n9336 & n9343 ) | ( n9342 & n9343 ) ;
  assign n9345 = n2476 & n2982 ;
  assign n9346 = x35 & n9345 ;
  assign n9347 = x94 & n2989 ;
  assign n9348 = x93 & n2986 ;
  assign n9349 = n9347 | n9348 ;
  assign n9350 = x92 & n3159 ;
  assign n9351 = n9349 | n9350 ;
  assign n9352 = ( ~x35 & n9345 ) | ( ~x35 & n9351 ) | ( n9345 & n9351 ) ;
  assign n9353 = x35 & ~n9351 ;
  assign n9354 = ( ~n9346 & n9352 ) | ( ~n9346 & n9353 ) | ( n9352 & n9353 ) ;
  assign n9355 = n1602 & n4020 ;
  assign n9356 = x41 & n9355 ;
  assign n9357 = x88 & n4027 ;
  assign n9358 = x87 & n4024 ;
  assign n9359 = n9357 | n9358 ;
  assign n9360 = x86 & n4223 ;
  assign n9361 = n9359 | n9360 ;
  assign n9362 = ( ~x41 & n9355 ) | ( ~x41 & n9361 ) | ( n9355 & n9361 ) ;
  assign n9363 = x41 & ~n9361 ;
  assign n9364 = ( ~n9356 & n9362 ) | ( ~n9356 & n9363 ) | ( n9362 & n9363 ) ;
  assign n9365 = n1006 & n5223 ;
  assign n9366 = x47 & n9365 ;
  assign n9367 = x82 & n5230 ;
  assign n9368 = x81 & n5227 ;
  assign n9369 = n9367 | n9368 ;
  assign n9370 = x80 & n5434 ;
  assign n9371 = n9369 | n9370 ;
  assign n9372 = ( ~x47 & n9365 ) | ( ~x47 & n9371 ) | ( n9365 & n9371 ) ;
  assign n9373 = x47 & ~n9371 ;
  assign n9374 = ( ~n9366 & n9372 ) | ( ~n9366 & n9373 ) | ( n9372 & n9373 ) ;
  assign n9375 = n565 & n6546 ;
  assign n9376 = x53 & n9375 ;
  assign n9377 = x76 & n6553 ;
  assign n9378 = x75 & n6550 ;
  assign n9379 = n9377 | n9378 ;
  assign n9380 = x74 & n6787 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = ( ~x53 & n9375 ) | ( ~x53 & n9381 ) | ( n9375 & n9381 ) ;
  assign n9383 = x53 & ~n9381 ;
  assign n9384 = ( ~n9376 & n9382 ) | ( ~n9376 & n9383 ) | ( n9382 & n9383 ) ;
  assign n9385 = n8869 | n9127 ;
  assign n9386 = x62 & n9385 ;
  assign n9387 = x67 & n8866 ;
  assign n9388 = x66 & n8863 ;
  assign n9389 = n9387 | n9388 ;
  assign n9390 = x65 & n9125 ;
  assign n9391 = n9389 | n9390 ;
  assign n9392 = n169 & n8859 ;
  assign n9393 = n9391 | n9392 ;
  assign n9394 = x62 & ~x63 ;
  assign n9395 = ~x62 & x63 ;
  assign n9396 = ( x64 & n9394 ) | ( x64 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9397 = ( n9386 & n9393 ) | ( n9386 & ~n9396 ) | ( n9393 & ~n9396 ) ;
  assign n9398 = ( n9386 & ~n9393 ) | ( n9386 & n9396 ) | ( ~n9393 & n9396 ) ;
  assign n9399 = ( ~n9386 & n9397 ) | ( ~n9386 & n9398 ) | ( n9397 & n9398 ) ;
  assign n9400 = n276 & n8067 ;
  assign n9401 = x59 & n9400 ;
  assign n9402 = x70 & n8074 ;
  assign n9403 = x69 & n8071 ;
  assign n9404 = n9402 | n9403 ;
  assign n9405 = x68 & n8298 ;
  assign n9406 = n9404 | n9405 ;
  assign n9407 = ( ~x59 & n9400 ) | ( ~x59 & n9406 ) | ( n9400 & n9406 ) ;
  assign n9408 = x59 & ~n9406 ;
  assign n9409 = ( ~n9401 & n9407 ) | ( ~n9401 & n9408 ) | ( n9407 & n9408 ) ;
  assign n9410 = ( n9142 & n9399 ) | ( n9142 & n9409 ) | ( n9399 & n9409 ) ;
  assign n9411 = ( ~n9142 & n9399 ) | ( ~n9142 & n9409 ) | ( n9399 & n9409 ) ;
  assign n9412 = ( n9142 & ~n9410 ) | ( n9142 & n9411 ) | ( ~n9410 & n9411 ) ;
  assign n9413 = n388 & n7277 ;
  assign n9414 = x56 & n9413 ;
  assign n9415 = x73 & n7545 ;
  assign n9416 = x72 & n7273 ;
  assign n9417 = n9415 | n9416 ;
  assign n9418 = x71 & n7552 ;
  assign n9419 = n9417 | n9418 ;
  assign n9420 = ( ~x56 & n9413 ) | ( ~x56 & n9419 ) | ( n9413 & n9419 ) ;
  assign n9421 = x56 & ~n9419 ;
  assign n9422 = ( ~n9414 & n9420 ) | ( ~n9414 & n9421 ) | ( n9420 & n9421 ) ;
  assign n9423 = ( n9156 & ~n9412 ) | ( n9156 & n9422 ) | ( ~n9412 & n9422 ) ;
  assign n9424 = ( n9156 & n9412 ) | ( n9156 & n9422 ) | ( n9412 & n9422 ) ;
  assign n9425 = ( n9412 & n9423 ) | ( n9412 & ~n9424 ) | ( n9423 & ~n9424 ) ;
  assign n9426 = ( n9158 & n9384 ) | ( n9158 & n9425 ) | ( n9384 & n9425 ) ;
  assign n9427 = ( ~n9158 & n9384 ) | ( ~n9158 & n9425 ) | ( n9384 & n9425 ) ;
  assign n9428 = ( n9158 & ~n9426 ) | ( n9158 & n9427 ) | ( ~n9426 & n9427 ) ;
  assign n9429 = n823 & n5858 ;
  assign n9430 = x50 & n9429 ;
  assign n9431 = x79 & n5865 ;
  assign n9432 = x78 & n5862 ;
  assign n9433 = n9431 | n9432 ;
  assign n9434 = x77 & n6092 ;
  assign n9435 = n9433 | n9434 ;
  assign n9436 = ( ~x50 & n9429 ) | ( ~x50 & n9435 ) | ( n9429 & n9435 ) ;
  assign n9437 = x50 & ~n9435 ;
  assign n9438 = ( ~n9430 & n9436 ) | ( ~n9430 & n9437 ) | ( n9436 & n9437 ) ;
  assign n9439 = ( n9172 & ~n9428 ) | ( n9172 & n9438 ) | ( ~n9428 & n9438 ) ;
  assign n9440 = ( n9172 & n9428 ) | ( n9172 & n9438 ) | ( n9428 & n9438 ) ;
  assign n9441 = ( n9428 & n9439 ) | ( n9428 & ~n9440 ) | ( n9439 & ~n9440 ) ;
  assign n9442 = ( n9174 & n9374 ) | ( n9174 & n9441 ) | ( n9374 & n9441 ) ;
  assign n9443 = ( ~n9174 & n9374 ) | ( ~n9174 & n9441 ) | ( n9374 & n9441 ) ;
  assign n9444 = ( n9174 & ~n9442 ) | ( n9174 & n9443 ) | ( ~n9442 & n9443 ) ;
  assign n9445 = n1368 & n4625 ;
  assign n9446 = x44 & n9445 ;
  assign n9447 = x85 & n4791 ;
  assign n9448 = x84 & n4621 ;
  assign n9449 = n9447 | n9448 ;
  assign n9450 = x83 & n4795 ;
  assign n9451 = n9449 | n9450 ;
  assign n9452 = ( ~x44 & n9445 ) | ( ~x44 & n9451 ) | ( n9445 & n9451 ) ;
  assign n9453 = x44 & ~n9451 ;
  assign n9454 = ( ~n9446 & n9452 ) | ( ~n9446 & n9453 ) | ( n9452 & n9453 ) ;
  assign n9455 = ( n9187 & ~n9444 ) | ( n9187 & n9454 ) | ( ~n9444 & n9454 ) ;
  assign n9456 = ( n9187 & n9444 ) | ( n9187 & n9454 ) | ( n9444 & n9454 ) ;
  assign n9457 = ( n9444 & n9455 ) | ( n9444 & ~n9456 ) | ( n9455 & ~n9456 ) ;
  assign n9458 = ( n9201 & n9364 ) | ( n9201 & n9457 ) | ( n9364 & n9457 ) ;
  assign n9459 = ( ~n9201 & n9364 ) | ( ~n9201 & n9457 ) | ( n9364 & n9457 ) ;
  assign n9460 = ( n9201 & ~n9458 ) | ( n9201 & n9459 ) | ( ~n9458 & n9459 ) ;
  assign n9461 = n1959 & n3492 ;
  assign n9462 = x38 & n9461 ;
  assign n9463 = x91 & n3499 ;
  assign n9464 = x90 & n3496 ;
  assign n9465 = n9463 | n9464 ;
  assign n9466 = x89 & n3662 ;
  assign n9467 = n9465 | n9466 ;
  assign n9468 = ( ~x38 & n9461 ) | ( ~x38 & n9467 ) | ( n9461 & n9467 ) ;
  assign n9469 = x38 & ~n9467 ;
  assign n9470 = ( ~n9462 & n9468 ) | ( ~n9462 & n9469 ) | ( n9468 & n9469 ) ;
  assign n9471 = ( n9203 & n9460 ) | ( n9203 & n9470 ) | ( n9460 & n9470 ) ;
  assign n9472 = ( n9203 & ~n9460 ) | ( n9203 & n9470 ) | ( ~n9460 & n9470 ) ;
  assign n9473 = ( n9460 & ~n9471 ) | ( n9460 & n9472 ) | ( ~n9471 & n9472 ) ;
  assign n9474 = ( n9217 & n9354 ) | ( n9217 & n9473 ) | ( n9354 & n9473 ) ;
  assign n9475 = ( ~n9217 & n9354 ) | ( ~n9217 & n9473 ) | ( n9354 & n9473 ) ;
  assign n9476 = ( n9217 & ~n9474 ) | ( n9217 & n9475 ) | ( ~n9474 & n9475 ) ;
  assign n9477 = n2545 & n2788 ;
  assign n9478 = x32 & n9477 ;
  assign n9479 = x97 & n2552 ;
  assign n9480 = x96 & n2549 ;
  assign n9481 = n9479 | n9480 ;
  assign n9482 = x95 & n2696 ;
  assign n9483 = n9481 | n9482 ;
  assign n9484 = ( ~x32 & n9477 ) | ( ~x32 & n9483 ) | ( n9477 & n9483 ) ;
  assign n9485 = x32 & ~n9483 ;
  assign n9486 = ( ~n9478 & n9484 ) | ( ~n9478 & n9485 ) | ( n9484 & n9485 ) ;
  assign n9487 = ( n9219 & n9476 ) | ( n9219 & n9486 ) | ( n9476 & n9486 ) ;
  assign n9488 = ( ~n9219 & n9476 ) | ( ~n9219 & n9486 ) | ( n9476 & n9486 ) ;
  assign n9489 = ( n9219 & ~n9487 ) | ( n9219 & n9488 ) | ( ~n9487 & n9488 ) ;
  assign n9490 = n2137 & n3264 ;
  assign n9491 = x29 & n9490 ;
  assign n9492 = x100 & n2144 ;
  assign n9493 = x99 & n2141 ;
  assign n9494 = n9492 | n9493 ;
  assign n9495 = x98 & n2267 ;
  assign n9496 = n9494 | n9495 ;
  assign n9497 = ( ~x29 & n9490 ) | ( ~x29 & n9496 ) | ( n9490 & n9496 ) ;
  assign n9498 = x29 & ~n9496 ;
  assign n9499 = ( ~n9491 & n9497 ) | ( ~n9491 & n9498 ) | ( n9497 & n9498 ) ;
  assign n9500 = ( n9233 & ~n9489 ) | ( n9233 & n9499 ) | ( ~n9489 & n9499 ) ;
  assign n9501 = ( n9233 & n9489 ) | ( n9233 & n9499 ) | ( n9489 & n9499 ) ;
  assign n9502 = ( n9489 & n9500 ) | ( n9489 & ~n9501 ) | ( n9500 & ~n9501 ) ;
  assign n9503 = ( n9235 & n9344 ) | ( n9235 & n9502 ) | ( n9344 & n9502 ) ;
  assign n9504 = ( ~n9235 & n9344 ) | ( ~n9235 & n9502 ) | ( n9344 & n9502 ) ;
  assign n9505 = ( n9235 & ~n9503 ) | ( n9235 & n9504 ) | ( ~n9503 & n9504 ) ;
  assign n9506 = n9249 & ~n9505 ;
  assign n9507 = ~n9249 & n9505 ;
  assign n9508 = n9506 | n9507 ;
  assign n9509 = ( ~n9251 & n9334 ) | ( ~n9251 & n9508 ) | ( n9334 & n9508 ) ;
  assign n9510 = ( n9251 & n9334 ) | ( n9251 & ~n9508 ) | ( n9334 & ~n9508 ) ;
  assign n9511 = ( ~n9334 & n9509 ) | ( ~n9334 & n9510 ) | ( n9509 & n9510 ) ;
  assign n9512 = n874 & n5558 ;
  assign n9513 = x17 & n9512 ;
  assign n9514 = x112 & n881 ;
  assign n9515 = x111 & n878 ;
  assign n9516 = n9514 | n9515 ;
  assign n9517 = x110 & n959 ;
  assign n9518 = n9516 | n9517 ;
  assign n9519 = ( ~x17 & n9512 ) | ( ~x17 & n9518 ) | ( n9512 & n9518 ) ;
  assign n9520 = x17 & ~n9518 ;
  assign n9521 = ( ~n9513 & n9519 ) | ( ~n9513 & n9520 ) | ( n9519 & n9520 ) ;
  assign n9522 = ( n9265 & n9511 ) | ( n9265 & n9521 ) | ( n9511 & n9521 ) ;
  assign n9523 = ( ~n9265 & n9511 ) | ( ~n9265 & n9521 ) | ( n9511 & n9521 ) ;
  assign n9524 = ( n9265 & ~n9522 ) | ( n9265 & n9523 ) | ( ~n9522 & n9523 ) ;
  assign n9525 = n649 & n6446 ;
  assign n9526 = x14 & n9525 ;
  assign n9527 = x115 & n656 ;
  assign n9528 = x114 & n653 ;
  assign n9529 = n9527 | n9528 ;
  assign n9530 = x113 & n744 ;
  assign n9531 = n9529 | n9530 ;
  assign n9532 = ( ~x14 & n9525 ) | ( ~x14 & n9531 ) | ( n9525 & n9531 ) ;
  assign n9533 = x14 & ~n9531 ;
  assign n9534 = ( ~n9526 & n9532 ) | ( ~n9526 & n9533 ) | ( n9532 & n9533 ) ;
  assign n9535 = ( n9267 & ~n9524 ) | ( n9267 & n9534 ) | ( ~n9524 & n9534 ) ;
  assign n9536 = ( n9267 & n9524 ) | ( n9267 & n9534 ) | ( n9524 & n9534 ) ;
  assign n9537 = ( n9524 & n9535 ) | ( n9524 & ~n9536 ) | ( n9535 & ~n9536 ) ;
  assign n9538 = n449 & n6940 ;
  assign n9539 = x11 & n9538 ;
  assign n9540 = x118 & n456 ;
  assign n9541 = x117 & n453 ;
  assign n9542 = n9540 | n9541 ;
  assign n9543 = x116 & n536 ;
  assign n9544 = n9542 | n9543 ;
  assign n9545 = ( ~x11 & n9538 ) | ( ~x11 & n9544 ) | ( n9538 & n9544 ) ;
  assign n9546 = x11 & ~n9544 ;
  assign n9547 = ( ~n9539 & n9545 ) | ( ~n9539 & n9546 ) | ( n9545 & n9546 ) ;
  assign n9548 = ( n9281 & ~n9537 ) | ( n9281 & n9547 ) | ( ~n9537 & n9547 ) ;
  assign n9549 = ( n9281 & n9537 ) | ( n9281 & n9547 ) | ( n9537 & n9547 ) ;
  assign n9550 = ( n9537 & n9548 ) | ( n9537 & ~n9549 ) | ( n9548 & ~n9549 ) ;
  assign n9551 = n206 & n8729 ;
  assign n9552 = x5 & n9551 ;
  assign n9553 = x124 & n205 ;
  assign n9554 = x123 & n201 ;
  assign n9555 = n9553 | n9554 ;
  assign n9556 = x122 & n221 ;
  assign n9557 = n9555 | n9556 ;
  assign n9558 = ( ~x5 & n9551 ) | ( ~x5 & n9557 ) | ( n9551 & n9557 ) ;
  assign n9559 = x5 & ~n9557 ;
  assign n9560 = ( ~n9552 & n9558 ) | ( ~n9552 & n9559 ) | ( n9558 & n9559 ) ;
  assign n9561 = n301 & n7696 ;
  assign n9562 = x8 & n9561 ;
  assign n9563 = x121 & n309 ;
  assign n9564 = x120 & n306 ;
  assign n9565 = n9563 | n9564 ;
  assign n9566 = x119 & n359 ;
  assign n9567 = n9565 | n9566 ;
  assign n9568 = ( ~x8 & n9561 ) | ( ~x8 & n9567 ) | ( n9561 & n9567 ) ;
  assign n9569 = x8 & ~n9567 ;
  assign n9570 = ( ~n9562 & n9568 ) | ( ~n9562 & n9569 ) | ( n9568 & n9569 ) ;
  assign n9571 = ( n9550 & n9560 ) | ( n9550 & n9570 ) | ( n9560 & n9570 ) ;
  assign n9572 = ( ~n9550 & n9560 ) | ( ~n9550 & n9570 ) | ( n9560 & n9570 ) ;
  assign n9573 = ( n9550 & ~n9571 ) | ( n9550 & n9572 ) | ( ~n9571 & n9572 ) ;
  assign n9574 = ( ~x125 & x127 ) | ( ~x125 & n9037 ) | ( x127 & n9037 ) ;
  assign n9575 = ( x125 & x127 ) | ( x125 & n9037 ) | ( x127 & n9037 ) ;
  assign n9576 = ( x125 & n9574 ) | ( x125 & ~n9575 ) | ( n9574 & ~n9575 ) ;
  assign n9577 = x0 & n9576 ;
  assign n9578 = ( x1 & x2 ) | ( x1 & n9577 ) | ( x2 & n9577 ) ;
  assign n9579 = x126 & n172 ;
  assign n9580 = x127 | n9579 ;
  assign n9581 = ( n147 & n9579 ) | ( n147 & n9580 ) | ( n9579 & n9580 ) ;
  assign n9582 = ( ~x125 & n135 ) | ( ~x125 & n174 ) | ( n135 & n174 ) ;
  assign n9583 = n9581 | n9582 ;
  assign n9584 = n9578 | n9583 ;
  assign n9585 = n9578 & n9583 ;
  assign n9586 = n9584 & ~n9585 ;
  assign n9587 = ( n9303 & n9573 ) | ( n9303 & n9586 ) | ( n9573 & n9586 ) ;
  assign n9588 = ( n9303 & ~n9573 ) | ( n9303 & n9586 ) | ( ~n9573 & n9586 ) ;
  assign n9589 = ( n9573 & ~n9587 ) | ( n9573 & n9588 ) | ( ~n9587 & n9588 ) ;
  assign n9590 = ( n9307 & ~n9310 ) | ( n9307 & n9589 ) | ( ~n9310 & n9589 ) ;
  assign n9591 = ( n9307 & n9310 ) | ( n9307 & n9589 ) | ( n9310 & n9589 ) ;
  assign n9592 = ( n9310 & n9590 ) | ( n9310 & ~n9591 ) | ( n9590 & ~n9591 ) ;
  assign n9593 = n449 & n7181 ;
  assign n9594 = x11 & n9593 ;
  assign n9595 = x118 & n453 ;
  assign n9596 = x117 & n536 ;
  assign n9597 = n9595 | n9596 ;
  assign n9598 = x119 & n456 ;
  assign n9599 = n9597 | n9598 ;
  assign n9600 = ( ~x11 & n9593 ) | ( ~x11 & n9599 ) | ( n9593 & n9599 ) ;
  assign n9601 = x11 & ~n9599 ;
  assign n9602 = ( ~n9594 & n9600 ) | ( ~n9594 & n9601 ) | ( n9600 & n9601 ) ;
  assign n9603 = n874 & n5774 ;
  assign n9604 = x17 & n9603 ;
  assign n9605 = x113 & n881 ;
  assign n9606 = x112 & n878 ;
  assign n9607 = n9605 | n9606 ;
  assign n9608 = x111 & n959 ;
  assign n9609 = n9607 | n9608 ;
  assign n9610 = ( ~x17 & n9603 ) | ( ~x17 & n9609 ) | ( n9603 & n9609 ) ;
  assign n9611 = x17 & ~n9609 ;
  assign n9612 = ( ~n9604 & n9610 ) | ( ~n9604 & n9611 ) | ( n9610 & n9611 ) ;
  assign n9613 = ( n9249 & n9331 ) | ( n9249 & n9505 ) | ( n9331 & n9505 ) ;
  assign n9614 = n1427 & n4523 ;
  assign n9615 = x23 & n9614 ;
  assign n9616 = x107 & n1434 ;
  assign n9617 = x106 & n1431 ;
  assign n9618 = n9616 | n9617 ;
  assign n9619 = x105 & n1531 ;
  assign n9620 = n9618 | n9619 ;
  assign n9621 = ( ~x23 & n9614 ) | ( ~x23 & n9620 ) | ( n9614 & n9620 ) ;
  assign n9622 = x23 & ~n9620 ;
  assign n9623 = ( ~n9615 & n9621 ) | ( ~n9615 & n9622 ) | ( n9621 & n9622 ) ;
  assign n9624 = n2137 & n3591 ;
  assign n9625 = x29 & n9624 ;
  assign n9626 = x101 & n2144 ;
  assign n9627 = x100 & n2141 ;
  assign n9628 = n9626 | n9627 ;
  assign n9629 = x99 & n2267 ;
  assign n9630 = n9628 | n9629 ;
  assign n9631 = ( ~x29 & n9624 ) | ( ~x29 & n9630 ) | ( n9624 & n9630 ) ;
  assign n9632 = x29 & ~n9630 ;
  assign n9633 = ( ~n9625 & n9631 ) | ( ~n9625 & n9632 ) | ( n9631 & n9632 ) ;
  assign n9634 = n2492 & n2982 ;
  assign n9635 = x35 & n9634 ;
  assign n9636 = x95 & n2989 ;
  assign n9637 = x94 & n2986 ;
  assign n9638 = n9636 | n9637 ;
  assign n9639 = x93 & n3159 ;
  assign n9640 = n9638 | n9639 ;
  assign n9641 = ( ~x35 & n9634 ) | ( ~x35 & n9640 ) | ( n9634 & n9640 ) ;
  assign n9642 = x35 & ~n9640 ;
  assign n9643 = ( ~n9635 & n9641 ) | ( ~n9635 & n9642 ) | ( n9641 & n9642 ) ;
  assign n9644 = n1822 & n4020 ;
  assign n9645 = x41 & n9644 ;
  assign n9646 = x89 & n4027 ;
  assign n9647 = x88 & n4024 ;
  assign n9648 = n9646 | n9647 ;
  assign n9649 = x87 & n4223 ;
  assign n9650 = n9648 | n9649 ;
  assign n9651 = ( ~x41 & n9644 ) | ( ~x41 & n9650 ) | ( n9644 & n9650 ) ;
  assign n9652 = x41 & ~n9650 ;
  assign n9653 = ( ~n9645 & n9651 ) | ( ~n9645 & n9652 ) | ( n9651 & n9652 ) ;
  assign n9654 = n1093 & n5223 ;
  assign n9655 = x47 & n9654 ;
  assign n9656 = x83 & n5230 ;
  assign n9657 = x82 & n5227 ;
  assign n9658 = n9656 | n9657 ;
  assign n9659 = x81 & n5434 ;
  assign n9660 = n9658 | n9659 ;
  assign n9661 = ( ~x47 & n9654 ) | ( ~x47 & n9660 ) | ( n9654 & n9660 ) ;
  assign n9662 = x47 & ~n9660 ;
  assign n9663 = ( ~n9655 & n9661 ) | ( ~n9655 & n9662 ) | ( n9661 & n9662 ) ;
  assign n9664 = n626 & n6546 ;
  assign n9665 = x53 & n9664 ;
  assign n9666 = x77 & n6553 ;
  assign n9667 = x76 & n6550 ;
  assign n9668 = n9666 | n9667 ;
  assign n9669 = x75 & n6787 ;
  assign n9670 = n9668 | n9669 ;
  assign n9671 = ( ~x53 & n9664 ) | ( ~x53 & n9670 ) | ( n9664 & n9670 ) ;
  assign n9672 = x53 & ~n9670 ;
  assign n9673 = ( ~n9665 & n9671 ) | ( ~n9665 & n9672 ) | ( n9671 & n9672 ) ;
  assign n9674 = x62 & ~n9393 ;
  assign n9675 = ( x62 & n9393 ) | ( x62 & n9397 ) | ( n9393 & n9397 ) ;
  assign n9676 = ( n9393 & n9674 ) | ( n9393 & ~n9675 ) | ( n9674 & ~n9675 ) ;
  assign n9677 = n193 & n8859 ;
  assign n9678 = x62 & n9677 ;
  assign n9679 = x68 & n8866 ;
  assign n9680 = x67 & n8863 ;
  assign n9681 = n9679 | n9680 ;
  assign n9682 = x66 & n9125 ;
  assign n9683 = n9681 | n9682 ;
  assign n9684 = ( ~x62 & n9677 ) | ( ~x62 & n9683 ) | ( n9677 & n9683 ) ;
  assign n9685 = x62 & ~n9683 ;
  assign n9686 = ( ~n9678 & n9684 ) | ( ~n9678 & n9685 ) | ( n9684 & n9685 ) ;
  assign n9687 = ( x62 & x63 ) | ( x62 & x65 ) | ( x63 & x65 ) ;
  assign n9688 = ( x62 & x64 ) | ( x62 & ~n9394 ) | ( x64 & ~n9394 ) ;
  assign n9689 = ( x64 & n9687 ) | ( x64 & ~n9688 ) | ( n9687 & ~n9688 ) ;
  assign n9690 = ( ~n9676 & n9686 ) | ( ~n9676 & n9689 ) | ( n9686 & n9689 ) ;
  assign n9691 = ( n9676 & n9686 ) | ( n9676 & n9689 ) | ( n9686 & n9689 ) ;
  assign n9692 = ( n9676 & n9690 ) | ( n9676 & ~n9691 ) | ( n9690 & ~n9691 ) ;
  assign n9693 = n322 & n8067 ;
  assign n9694 = x59 & n9693 ;
  assign n9695 = x71 & n8074 ;
  assign n9696 = x70 & n8071 ;
  assign n9697 = n9695 | n9696 ;
  assign n9698 = x69 & n8298 ;
  assign n9699 = n9697 | n9698 ;
  assign n9700 = ( ~x59 & n9693 ) | ( ~x59 & n9699 ) | ( n9693 & n9699 ) ;
  assign n9701 = x59 & ~n9699 ;
  assign n9702 = ( ~n9694 & n9700 ) | ( ~n9694 & n9701 ) | ( n9700 & n9701 ) ;
  assign n9703 = ( n9410 & n9692 ) | ( n9410 & n9702 ) | ( n9692 & n9702 ) ;
  assign n9704 = ( ~n9410 & n9692 ) | ( ~n9410 & n9702 ) | ( n9692 & n9702 ) ;
  assign n9705 = ( n9410 & ~n9703 ) | ( n9410 & n9704 ) | ( ~n9703 & n9704 ) ;
  assign n9706 = n436 & n7277 ;
  assign n9707 = x56 & n9706 ;
  assign n9708 = x74 & n7545 ;
  assign n9709 = x73 & n7273 ;
  assign n9710 = n9708 | n9709 ;
  assign n9711 = x72 & n7552 ;
  assign n9712 = n9710 | n9711 ;
  assign n9713 = ( ~x56 & n9706 ) | ( ~x56 & n9712 ) | ( n9706 & n9712 ) ;
  assign n9714 = x56 & ~n9712 ;
  assign n9715 = ( ~n9707 & n9713 ) | ( ~n9707 & n9714 ) | ( n9713 & n9714 ) ;
  assign n9716 = ( n9424 & ~n9705 ) | ( n9424 & n9715 ) | ( ~n9705 & n9715 ) ;
  assign n9717 = ( n9424 & n9705 ) | ( n9424 & n9715 ) | ( n9705 & n9715 ) ;
  assign n9718 = ( n9705 & n9716 ) | ( n9705 & ~n9717 ) | ( n9716 & ~n9717 ) ;
  assign n9719 = ( n9426 & n9673 ) | ( n9426 & n9718 ) | ( n9673 & n9718 ) ;
  assign n9720 = ( ~n9426 & n9673 ) | ( ~n9426 & n9718 ) | ( n9673 & n9718 ) ;
  assign n9721 = ( n9426 & ~n9719 ) | ( n9426 & n9720 ) | ( ~n9719 & n9720 ) ;
  assign n9722 = n840 & n5858 ;
  assign n9723 = x50 & n9722 ;
  assign n9724 = x80 & n5865 ;
  assign n9725 = x79 & n5862 ;
  assign n9726 = n9724 | n9725 ;
  assign n9727 = x78 & n6092 ;
  assign n9728 = n9726 | n9727 ;
  assign n9729 = ( ~x50 & n9722 ) | ( ~x50 & n9728 ) | ( n9722 & n9728 ) ;
  assign n9730 = x50 & ~n9728 ;
  assign n9731 = ( ~n9723 & n9729 ) | ( ~n9723 & n9730 ) | ( n9729 & n9730 ) ;
  assign n9732 = ( n9440 & ~n9721 ) | ( n9440 & n9731 ) | ( ~n9721 & n9731 ) ;
  assign n9733 = ( n9440 & n9721 ) | ( n9440 & n9731 ) | ( n9721 & n9731 ) ;
  assign n9734 = ( n9721 & n9732 ) | ( n9721 & ~n9733 ) | ( n9732 & ~n9733 ) ;
  assign n9735 = ( n9442 & n9663 ) | ( n9442 & n9734 ) | ( n9663 & n9734 ) ;
  assign n9736 = ( ~n9442 & n9663 ) | ( ~n9442 & n9734 ) | ( n9663 & n9734 ) ;
  assign n9737 = ( n9442 & ~n9735 ) | ( n9442 & n9736 ) | ( ~n9735 & n9736 ) ;
  assign n9738 = n1384 & n4625 ;
  assign n9739 = x44 & n9738 ;
  assign n9740 = x86 & n4791 ;
  assign n9741 = x85 & n4621 ;
  assign n9742 = n9740 | n9741 ;
  assign n9743 = x84 & n4795 ;
  assign n9744 = n9742 | n9743 ;
  assign n9745 = ( ~x44 & n9738 ) | ( ~x44 & n9744 ) | ( n9738 & n9744 ) ;
  assign n9746 = x44 & ~n9744 ;
  assign n9747 = ( ~n9739 & n9745 ) | ( ~n9739 & n9746 ) | ( n9745 & n9746 ) ;
  assign n9748 = ( n9456 & ~n9737 ) | ( n9456 & n9747 ) | ( ~n9737 & n9747 ) ;
  assign n9749 = ( n9456 & n9737 ) | ( n9456 & n9747 ) | ( n9737 & n9747 ) ;
  assign n9750 = ( n9737 & n9748 ) | ( n9737 & ~n9749 ) | ( n9748 & ~n9749 ) ;
  assign n9751 = ( n9458 & n9653 ) | ( n9458 & n9750 ) | ( n9653 & n9750 ) ;
  assign n9752 = ( ~n9458 & n9653 ) | ( ~n9458 & n9750 ) | ( n9653 & n9750 ) ;
  assign n9753 = ( n9458 & ~n9751 ) | ( n9458 & n9752 ) | ( ~n9751 & n9752 ) ;
  assign n9754 = n2083 & n3492 ;
  assign n9755 = x38 & n9754 ;
  assign n9756 = x92 & n3499 ;
  assign n9757 = x91 & n3496 ;
  assign n9758 = n9756 | n9757 ;
  assign n9759 = x90 & n3662 ;
  assign n9760 = n9758 | n9759 ;
  assign n9761 = ( ~x38 & n9754 ) | ( ~x38 & n9760 ) | ( n9754 & n9760 ) ;
  assign n9762 = x38 & ~n9760 ;
  assign n9763 = ( ~n9755 & n9761 ) | ( ~n9755 & n9762 ) | ( n9761 & n9762 ) ;
  assign n9764 = ( n9471 & n9753 ) | ( n9471 & n9763 ) | ( n9753 & n9763 ) ;
  assign n9765 = ( n9471 & ~n9753 ) | ( n9471 & n9763 ) | ( ~n9753 & n9763 ) ;
  assign n9766 = ( n9753 & ~n9764 ) | ( n9753 & n9765 ) | ( ~n9764 & n9765 ) ;
  assign n9767 = ( n9474 & n9643 ) | ( n9474 & n9766 ) | ( n9643 & n9766 ) ;
  assign n9768 = ( ~n9474 & n9643 ) | ( ~n9474 & n9766 ) | ( n9643 & n9766 ) ;
  assign n9769 = ( n9474 & ~n9767 ) | ( n9474 & n9768 ) | ( ~n9767 & n9768 ) ;
  assign n9770 = n2545 & n2939 ;
  assign n9771 = x32 & n9770 ;
  assign n9772 = x98 & n2552 ;
  assign n9773 = x97 & n2549 ;
  assign n9774 = n9772 | n9773 ;
  assign n9775 = x96 & n2696 ;
  assign n9776 = n9774 | n9775 ;
  assign n9777 = ( ~x32 & n9770 ) | ( ~x32 & n9776 ) | ( n9770 & n9776 ) ;
  assign n9778 = x32 & ~n9776 ;
  assign n9779 = ( ~n9771 & n9777 ) | ( ~n9771 & n9778 ) | ( n9777 & n9778 ) ;
  assign n9780 = ( n9487 & ~n9769 ) | ( n9487 & n9779 ) | ( ~n9769 & n9779 ) ;
  assign n9781 = ( n9487 & n9769 ) | ( n9487 & n9779 ) | ( n9769 & n9779 ) ;
  assign n9782 = ( n9769 & n9780 ) | ( n9769 & ~n9781 ) | ( n9780 & ~n9781 ) ;
  assign n9783 = ( n9501 & n9633 ) | ( n9501 & n9782 ) | ( n9633 & n9782 ) ;
  assign n9784 = ( ~n9501 & n9633 ) | ( ~n9501 & n9782 ) | ( n9633 & n9782 ) ;
  assign n9785 = ( n9501 & ~n9783 ) | ( n9501 & n9784 ) | ( ~n9783 & n9784 ) ;
  assign n9786 = n1755 & n3957 ;
  assign n9787 = x26 & n9786 ;
  assign n9788 = x104 & n1762 ;
  assign n9789 = x103 & n1759 ;
  assign n9790 = n9788 | n9789 ;
  assign n9791 = x102 & n1895 ;
  assign n9792 = n9790 | n9791 ;
  assign n9793 = ( ~x26 & n9786 ) | ( ~x26 & n9792 ) | ( n9786 & n9792 ) ;
  assign n9794 = x26 & ~n9792 ;
  assign n9795 = ( ~n9787 & n9793 ) | ( ~n9787 & n9794 ) | ( n9793 & n9794 ) ;
  assign n9796 = ( n9503 & ~n9785 ) | ( n9503 & n9795 ) | ( ~n9785 & n9795 ) ;
  assign n9797 = ( n9503 & n9785 ) | ( n9503 & n9795 ) | ( n9785 & n9795 ) ;
  assign n9798 = ( n9785 & n9796 ) | ( n9785 & ~n9797 ) | ( n9796 & ~n9797 ) ;
  assign n9799 = ( n9613 & n9623 ) | ( n9613 & n9798 ) | ( n9623 & n9798 ) ;
  assign n9800 = ( ~n9613 & n9623 ) | ( ~n9613 & n9798 ) | ( n9623 & n9798 ) ;
  assign n9801 = ( n9613 & ~n9799 ) | ( n9613 & n9800 ) | ( ~n9799 & n9800 ) ;
  assign n9802 = ( n9249 & n9331 ) | ( n9249 & ~n9505 ) | ( n9331 & ~n9505 ) ;
  assign n9803 = ( n9505 & ~n9613 ) | ( n9505 & n9802 ) | ( ~n9613 & n9802 ) ;
  assign n9804 = ( n9251 & n9321 ) | ( n9251 & n9803 ) | ( n9321 & n9803 ) ;
  assign n9805 = n1146 & n5331 ;
  assign n9806 = x20 & n9805 ;
  assign n9807 = x110 & n1153 ;
  assign n9808 = x109 & n1150 ;
  assign n9809 = n9807 | n9808 ;
  assign n9810 = x108 & n1217 ;
  assign n9811 = n9809 | n9810 ;
  assign n9812 = ( ~x20 & n9805 ) | ( ~x20 & n9811 ) | ( n9805 & n9811 ) ;
  assign n9813 = x20 & ~n9811 ;
  assign n9814 = ( ~n9806 & n9812 ) | ( ~n9806 & n9813 ) | ( n9812 & n9813 ) ;
  assign n9815 = ( ~n9801 & n9804 ) | ( ~n9801 & n9814 ) | ( n9804 & n9814 ) ;
  assign n9816 = ( n9801 & n9804 ) | ( n9801 & n9814 ) | ( n9804 & n9814 ) ;
  assign n9817 = ( n9801 & n9815 ) | ( n9801 & ~n9816 ) | ( n9815 & ~n9816 ) ;
  assign n9818 = ( n9522 & n9612 ) | ( n9522 & n9817 ) | ( n9612 & n9817 ) ;
  assign n9819 = ( ~n9522 & n9612 ) | ( ~n9522 & n9817 ) | ( n9612 & n9817 ) ;
  assign n9820 = ( n9522 & ~n9818 ) | ( n9522 & n9819 ) | ( ~n9818 & n9819 ) ;
  assign n9821 = n649 & n6462 ;
  assign n9822 = x14 & n9821 ;
  assign n9823 = x116 & n656 ;
  assign n9824 = x115 & n653 ;
  assign n9825 = n9823 | n9824 ;
  assign n9826 = x114 & n744 ;
  assign n9827 = n9825 | n9826 ;
  assign n9828 = ( ~x14 & n9821 ) | ( ~x14 & n9827 ) | ( n9821 & n9827 ) ;
  assign n9829 = x14 & ~n9827 ;
  assign n9830 = ( ~n9822 & n9828 ) | ( ~n9822 & n9829 ) | ( n9828 & n9829 ) ;
  assign n9831 = ( n9536 & ~n9820 ) | ( n9536 & n9830 ) | ( ~n9820 & n9830 ) ;
  assign n9832 = ( n9536 & n9820 ) | ( n9536 & n9830 ) | ( n9820 & n9830 ) ;
  assign n9833 = ( n9820 & n9831 ) | ( n9820 & ~n9832 ) | ( n9831 & ~n9832 ) ;
  assign n9834 = ( n9549 & n9602 ) | ( n9549 & n9833 ) | ( n9602 & n9833 ) ;
  assign n9835 = ( ~n9549 & n9602 ) | ( ~n9549 & n9833 ) | ( n9602 & n9833 ) ;
  assign n9836 = ( n9549 & ~n9834 ) | ( n9549 & n9835 ) | ( ~n9834 & n9835 ) ;
  assign n9837 = n206 & n9009 ;
  assign n9838 = x5 & n9837 ;
  assign n9839 = x125 & n205 ;
  assign n9840 = x124 & n201 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = x123 & n221 ;
  assign n9843 = n9841 | n9842 ;
  assign n9844 = ( ~x5 & n9837 ) | ( ~x5 & n9843 ) | ( n9837 & n9843 ) ;
  assign n9845 = x5 & ~n9843 ;
  assign n9846 = ( ~n9838 & n9844 ) | ( ~n9838 & n9845 ) | ( n9844 & n9845 ) ;
  assign n9847 = n301 & n8207 ;
  assign n9848 = x8 & n9847 ;
  assign n9849 = x122 & n309 ;
  assign n9850 = x121 & n306 ;
  assign n9851 = n9849 | n9850 ;
  assign n9852 = x120 & n359 ;
  assign n9853 = n9851 | n9852 ;
  assign n9854 = ( ~x8 & n9847 ) | ( ~x8 & n9853 ) | ( n9847 & n9853 ) ;
  assign n9855 = x8 & ~n9853 ;
  assign n9856 = ( ~n9848 & n9854 ) | ( ~n9848 & n9855 ) | ( n9854 & n9855 ) ;
  assign n9857 = ( n9836 & n9846 ) | ( n9836 & n9856 ) | ( n9846 & n9856 ) ;
  assign n9858 = ( ~n9836 & n9846 ) | ( ~n9836 & n9856 ) | ( n9846 & n9856 ) ;
  assign n9859 = ( n9836 & ~n9857 ) | ( n9836 & n9858 ) | ( ~n9857 & n9858 ) ;
  assign n9860 = x126 & n136 ;
  assign n9861 = x127 & n172 ;
  assign n9862 = n146 | n9861 ;
  assign n9863 = ~x126 & x127 ;
  assign n9864 = x126 | n9036 ;
  assign n9865 = x127 & n9864 ;
  assign n9866 = ( ~n9036 & n9864 ) | ( ~n9036 & n9865 ) | ( n9864 & n9865 ) ;
  assign n9867 = ( x126 & n9863 ) | ( x126 & ~n9866 ) | ( n9863 & ~n9866 ) ;
  assign n9868 = ( n9861 & n9862 ) | ( n9861 & n9867 ) | ( n9862 & n9867 ) ;
  assign n9869 = ( x2 & ~n9860 ) | ( x2 & n9868 ) | ( ~n9860 & n9868 ) ;
  assign n9870 = ( x2 & n9860 ) | ( x2 & n9868 ) | ( n9860 & n9868 ) ;
  assign n9871 = n9869 & ~n9870 ;
  assign n9872 = ( n9571 & ~n9859 ) | ( n9571 & n9871 ) | ( ~n9859 & n9871 ) ;
  assign n9873 = ( n9571 & n9859 ) | ( n9571 & n9871 ) | ( n9859 & n9871 ) ;
  assign n9874 = ( n9859 & n9872 ) | ( n9859 & ~n9873 ) | ( n9872 & ~n9873 ) ;
  assign n9875 = ( n9587 & n9591 ) | ( n9587 & n9874 ) | ( n9591 & n9874 ) ;
  assign n9876 = ( n9587 & ~n9591 ) | ( n9587 & n9874 ) | ( ~n9591 & n9874 ) ;
  assign n9877 = ( n9591 & ~n9875 ) | ( n9591 & n9876 ) | ( ~n9875 & n9876 ) ;
  assign n9878 = n649 & n6924 ;
  assign n9879 = x14 & n9878 ;
  assign n9880 = x117 & n656 ;
  assign n9881 = x116 & n653 ;
  assign n9882 = n9880 | n9881 ;
  assign n9883 = x115 & n744 ;
  assign n9884 = n9882 | n9883 ;
  assign n9885 = ( ~x14 & n9878 ) | ( ~x14 & n9884 ) | ( n9878 & n9884 ) ;
  assign n9886 = x14 & ~n9884 ;
  assign n9887 = ( ~n9879 & n9885 ) | ( ~n9879 & n9886 ) | ( n9885 & n9886 ) ;
  assign n9888 = n1146 & n5347 ;
  assign n9889 = x20 & n9888 ;
  assign n9890 = x111 & n1153 ;
  assign n9891 = x110 & n1150 ;
  assign n9892 = n9890 | n9891 ;
  assign n9893 = x109 & n1217 ;
  assign n9894 = n9892 | n9893 ;
  assign n9895 = ( ~x20 & n9888 ) | ( ~x20 & n9894 ) | ( n9888 & n9894 ) ;
  assign n9896 = x20 & ~n9894 ;
  assign n9897 = ( ~n9889 & n9895 ) | ( ~n9889 & n9896 ) | ( n9895 & n9896 ) ;
  assign n9898 = n2137 & n3764 ;
  assign n9899 = x29 & n9898 ;
  assign n9900 = x102 & n2144 ;
  assign n9901 = x101 & n2141 ;
  assign n9902 = n9900 | n9901 ;
  assign n9903 = x100 & n2267 ;
  assign n9904 = n9902 | n9903 ;
  assign n9905 = ( ~x29 & n9898 ) | ( ~x29 & n9904 ) | ( n9898 & n9904 ) ;
  assign n9906 = x29 & ~n9904 ;
  assign n9907 = ( ~n9899 & n9905 ) | ( ~n9899 & n9906 ) | ( n9905 & n9906 ) ;
  assign n9908 = n2772 & n2982 ;
  assign n9909 = x35 & n9908 ;
  assign n9910 = x96 & n2989 ;
  assign n9911 = x95 & n2986 ;
  assign n9912 = n9910 | n9911 ;
  assign n9913 = x94 & n3159 ;
  assign n9914 = n9912 | n9913 ;
  assign n9915 = ( ~x35 & n9908 ) | ( ~x35 & n9914 ) | ( n9908 & n9914 ) ;
  assign n9916 = x35 & ~n9914 ;
  assign n9917 = ( ~n9909 & n9915 ) | ( ~n9909 & n9916 ) | ( n9915 & n9916 ) ;
  assign n9918 = n2220 & n3492 ;
  assign n9919 = x38 & n9918 ;
  assign n9920 = x93 & n3499 ;
  assign n9921 = x92 & n3496 ;
  assign n9922 = n9920 | n9921 ;
  assign n9923 = x91 & n3662 ;
  assign n9924 = n9922 | n9923 ;
  assign n9925 = ( ~x38 & n9918 ) | ( ~x38 & n9924 ) | ( n9918 & n9924 ) ;
  assign n9926 = x38 & ~n9924 ;
  assign n9927 = ( ~n9919 & n9925 ) | ( ~n9919 & n9926 ) | ( n9925 & n9926 ) ;
  assign n9928 = n1494 & n4625 ;
  assign n9929 = x44 & n9928 ;
  assign n9930 = x87 & n4791 ;
  assign n9931 = x86 & n4621 ;
  assign n9932 = n9930 | n9931 ;
  assign n9933 = x85 & n4795 ;
  assign n9934 = n9932 | n9933 ;
  assign n9935 = ( ~x44 & n9928 ) | ( ~x44 & n9934 ) | ( n9928 & n9934 ) ;
  assign n9936 = x44 & ~n9934 ;
  assign n9937 = ( ~n9929 & n9935 ) | ( ~n9929 & n9936 ) | ( n9935 & n9936 ) ;
  assign n9938 = n1190 & n5223 ;
  assign n9939 = x47 & n9938 ;
  assign n9940 = x84 & n5230 ;
  assign n9941 = x83 & n5227 ;
  assign n9942 = n9940 | n9941 ;
  assign n9943 = x82 & n5434 ;
  assign n9944 = n9942 | n9943 ;
  assign n9945 = ( ~x47 & n9938 ) | ( ~x47 & n9944 ) | ( n9938 & n9944 ) ;
  assign n9946 = x47 & ~n9944 ;
  assign n9947 = ( ~n9939 & n9945 ) | ( ~n9939 & n9946 ) | ( n9945 & n9946 ) ;
  assign n9948 = n697 & n6546 ;
  assign n9949 = x53 & n9948 ;
  assign n9950 = x78 & n6553 ;
  assign n9951 = x77 & n6550 ;
  assign n9952 = n9950 | n9951 ;
  assign n9953 = x76 & n6787 ;
  assign n9954 = n9952 | n9953 ;
  assign n9955 = ( ~x53 & n9948 ) | ( ~x53 & n9954 ) | ( n9948 & n9954 ) ;
  assign n9956 = x53 & ~n9954 ;
  assign n9957 = ( ~n9949 & n9955 ) | ( ~n9949 & n9956 ) | ( n9955 & n9956 ) ;
  assign n9958 = n508 & n7277 ;
  assign n9959 = x56 & n9958 ;
  assign n9960 = x75 & n7545 ;
  assign n9961 = x74 & n7273 ;
  assign n9962 = n9960 | n9961 ;
  assign n9963 = x73 & n7552 ;
  assign n9964 = n9962 | n9963 ;
  assign n9965 = ( ~x56 & n9958 ) | ( ~x56 & n9964 ) | ( n9958 & n9964 ) ;
  assign n9966 = x56 & ~n9964 ;
  assign n9967 = ( ~n9959 & n9965 ) | ( ~n9959 & n9966 ) | ( n9965 & n9966 ) ;
  assign n9968 = n240 & n8859 ;
  assign n9969 = x62 & n9968 ;
  assign n9970 = x69 & n8866 ;
  assign n9971 = x68 & n8863 ;
  assign n9972 = n9970 | n9971 ;
  assign n9973 = x67 & n9125 ;
  assign n9974 = n9972 | n9973 ;
  assign n9975 = ( ~x62 & n9968 ) | ( ~x62 & n9974 ) | ( n9968 & n9974 ) ;
  assign n9976 = x62 & ~n9974 ;
  assign n9977 = ( ~n9969 & n9975 ) | ( ~n9969 & n9976 ) | ( n9975 & n9976 ) ;
  assign n9978 = ( x62 & x63 ) | ( x62 & x66 ) | ( x63 & x66 ) ;
  assign n9979 = ( x62 & x65 ) | ( x62 & ~n9394 ) | ( x65 & ~n9394 ) ;
  assign n9980 = ( x65 & n9978 ) | ( x65 & ~n9979 ) | ( n9978 & ~n9979 ) ;
  assign n9981 = ( n9691 & n9977 ) | ( n9691 & n9980 ) | ( n9977 & n9980 ) ;
  assign n9982 = ( ~n9691 & n9977 ) | ( ~n9691 & n9980 ) | ( n9977 & n9980 ) ;
  assign n9983 = ( n9691 & ~n9981 ) | ( n9691 & n9982 ) | ( ~n9981 & n9982 ) ;
  assign n9984 = n372 & n8067 ;
  assign n9985 = x59 & n9984 ;
  assign n9986 = x72 & n8074 ;
  assign n9987 = x71 & n8071 ;
  assign n9988 = n9986 | n9987 ;
  assign n9989 = x70 & n8298 ;
  assign n9990 = n9988 | n9989 ;
  assign n9991 = ( ~x59 & n9984 ) | ( ~x59 & n9990 ) | ( n9984 & n9990 ) ;
  assign n9992 = x59 & ~n9990 ;
  assign n9993 = ( ~n9985 & n9991 ) | ( ~n9985 & n9992 ) | ( n9991 & n9992 ) ;
  assign n9994 = ( n9703 & ~n9983 ) | ( n9703 & n9993 ) | ( ~n9983 & n9993 ) ;
  assign n9995 = ( n9703 & n9983 ) | ( n9703 & n9993 ) | ( n9983 & n9993 ) ;
  assign n9996 = ( n9983 & n9994 ) | ( n9983 & ~n9995 ) | ( n9994 & ~n9995 ) ;
  assign n9997 = ( n9717 & n9967 ) | ( n9717 & n9996 ) | ( n9967 & n9996 ) ;
  assign n9998 = ( ~n9717 & n9967 ) | ( ~n9717 & n9996 ) | ( n9967 & n9996 ) ;
  assign n9999 = ( n9717 & ~n9997 ) | ( n9717 & n9998 ) | ( ~n9997 & n9998 ) ;
  assign n10000 = ( n9719 & n9957 ) | ( n9719 & n9999 ) | ( n9957 & n9999 ) ;
  assign n10001 = ( ~n9719 & n9957 ) | ( ~n9719 & n9999 ) | ( n9957 & n9999 ) ;
  assign n10002 = ( n9719 & ~n10000 ) | ( n9719 & n10001 ) | ( ~n10000 & n10001 ) ;
  assign n10003 = n990 & n5858 ;
  assign n10004 = x50 & n10003 ;
  assign n10005 = x81 & n5865 ;
  assign n10006 = x80 & n5862 ;
  assign n10007 = n10005 | n10006 ;
  assign n10008 = x79 & n6092 ;
  assign n10009 = n10007 | n10008 ;
  assign n10010 = ( ~x50 & n10003 ) | ( ~x50 & n10009 ) | ( n10003 & n10009 ) ;
  assign n10011 = x50 & ~n10009 ;
  assign n10012 = ( ~n10004 & n10010 ) | ( ~n10004 & n10011 ) | ( n10010 & n10011 ) ;
  assign n10013 = ( n9733 & ~n10002 ) | ( n9733 & n10012 ) | ( ~n10002 & n10012 ) ;
  assign n10014 = ( n9733 & n10002 ) | ( n9733 & n10012 ) | ( n10002 & n10012 ) ;
  assign n10015 = ( n10002 & n10013 ) | ( n10002 & ~n10014 ) | ( n10013 & ~n10014 ) ;
  assign n10016 = ( n9735 & n9947 ) | ( n9735 & n10015 ) | ( n9947 & n10015 ) ;
  assign n10017 = ( ~n9735 & n9947 ) | ( ~n9735 & n10015 ) | ( n9947 & n10015 ) ;
  assign n10018 = ( n9735 & ~n10016 ) | ( n9735 & n10017 ) | ( ~n10016 & n10017 ) ;
  assign n10019 = ( n9749 & n9937 ) | ( n9749 & n10018 ) | ( n9937 & n10018 ) ;
  assign n10020 = ( ~n9749 & n9937 ) | ( ~n9749 & n10018 ) | ( n9937 & n10018 ) ;
  assign n10021 = ( n9749 & ~n10019 ) | ( n9749 & n10020 ) | ( ~n10019 & n10020 ) ;
  assign n10022 = n1838 & n4020 ;
  assign n10023 = x41 & n10022 ;
  assign n10024 = x90 & n4027 ;
  assign n10025 = x89 & n4024 ;
  assign n10026 = n10024 | n10025 ;
  assign n10027 = x88 & n4223 ;
  assign n10028 = n10026 | n10027 ;
  assign n10029 = ( ~x41 & n10022 ) | ( ~x41 & n10028 ) | ( n10022 & n10028 ) ;
  assign n10030 = x41 & ~n10028 ;
  assign n10031 = ( ~n10023 & n10029 ) | ( ~n10023 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10032 = ( n9751 & ~n10021 ) | ( n9751 & n10031 ) | ( ~n10021 & n10031 ) ;
  assign n10033 = ( n9751 & n10021 ) | ( n9751 & n10031 ) | ( n10021 & n10031 ) ;
  assign n10034 = ( n10021 & n10032 ) | ( n10021 & ~n10033 ) | ( n10032 & ~n10033 ) ;
  assign n10035 = ( ~n9764 & n9927 ) | ( ~n9764 & n10034 ) | ( n9927 & n10034 ) ;
  assign n10036 = ( n9764 & n9927 ) | ( n9764 & n10034 ) | ( n9927 & n10034 ) ;
  assign n10037 = ( n9764 & n10035 ) | ( n9764 & ~n10036 ) | ( n10035 & ~n10036 ) ;
  assign n10038 = ( n9767 & n9917 ) | ( n9767 & n10037 ) | ( n9917 & n10037 ) ;
  assign n10039 = ( ~n9767 & n9917 ) | ( ~n9767 & n10037 ) | ( n9917 & n10037 ) ;
  assign n10040 = ( n9767 & ~n10038 ) | ( n9767 & n10039 ) | ( ~n10038 & n10039 ) ;
  assign n10041 = n2545 & n3248 ;
  assign n10042 = x32 & n10041 ;
  assign n10043 = x99 & n2552 ;
  assign n10044 = x98 & n2549 ;
  assign n10045 = n10043 | n10044 ;
  assign n10046 = x97 & n2696 ;
  assign n10047 = n10045 | n10046 ;
  assign n10048 = ( ~x32 & n10041 ) | ( ~x32 & n10047 ) | ( n10041 & n10047 ) ;
  assign n10049 = x32 & ~n10047 ;
  assign n10050 = ( ~n10042 & n10048 ) | ( ~n10042 & n10049 ) | ( n10048 & n10049 ) ;
  assign n10051 = ( n9781 & ~n10040 ) | ( n9781 & n10050 ) | ( ~n10040 & n10050 ) ;
  assign n10052 = ( n9781 & n10040 ) | ( n9781 & n10050 ) | ( n10040 & n10050 ) ;
  assign n10053 = ( n10040 & n10051 ) | ( n10040 & ~n10052 ) | ( n10051 & ~n10052 ) ;
  assign n10054 = ( n9783 & n9907 ) | ( n9783 & n10053 ) | ( n9907 & n10053 ) ;
  assign n10055 = ( ~n9783 & n9907 ) | ( ~n9783 & n10053 ) | ( n9907 & n10053 ) ;
  assign n10056 = ( n9783 & ~n10054 ) | ( n9783 & n10055 ) | ( ~n10054 & n10055 ) ;
  assign n10057 = n1755 & n4145 ;
  assign n10058 = x26 & n10057 ;
  assign n10059 = x105 & n1762 ;
  assign n10060 = x104 & n1759 ;
  assign n10061 = n10059 | n10060 ;
  assign n10062 = x103 & n1895 ;
  assign n10063 = n10061 | n10062 ;
  assign n10064 = ( ~x26 & n10057 ) | ( ~x26 & n10063 ) | ( n10057 & n10063 ) ;
  assign n10065 = x26 & ~n10063 ;
  assign n10066 = ( ~n10058 & n10064 ) | ( ~n10058 & n10065 ) | ( n10064 & n10065 ) ;
  assign n10067 = ( n9797 & n10056 ) | ( n9797 & n10066 ) | ( n10056 & n10066 ) ;
  assign n10068 = ( ~n9797 & n10056 ) | ( ~n9797 & n10066 ) | ( n10056 & n10066 ) ;
  assign n10069 = ( n9797 & ~n10067 ) | ( n9797 & n10068 ) | ( ~n10067 & n10068 ) ;
  assign n10070 = n1427 & n4914 ;
  assign n10071 = x23 & n10070 ;
  assign n10072 = x108 & n1434 ;
  assign n10073 = x107 & n1431 ;
  assign n10074 = n10072 | n10073 ;
  assign n10075 = x106 & n1531 ;
  assign n10076 = n10074 | n10075 ;
  assign n10077 = ( ~x23 & n10070 ) | ( ~x23 & n10076 ) | ( n10070 & n10076 ) ;
  assign n10078 = x23 & ~n10076 ;
  assign n10079 = ( ~n10071 & n10077 ) | ( ~n10071 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10080 = ( n9799 & ~n10069 ) | ( n9799 & n10079 ) | ( ~n10069 & n10079 ) ;
  assign n10081 = ( n9799 & n10069 ) | ( n9799 & n10079 ) | ( n10069 & n10079 ) ;
  assign n10082 = ( n10069 & n10080 ) | ( n10069 & ~n10081 ) | ( n10080 & ~n10081 ) ;
  assign n10083 = ( n9816 & n9897 ) | ( n9816 & n10082 ) | ( n9897 & n10082 ) ;
  assign n10084 = ( ~n9816 & n9897 ) | ( ~n9816 & n10082 ) | ( n9897 & n10082 ) ;
  assign n10085 = ( n9816 & ~n10083 ) | ( n9816 & n10084 ) | ( ~n10083 & n10084 ) ;
  assign n10086 = n874 & n6002 ;
  assign n10087 = x17 & n10086 ;
  assign n10088 = x114 & n881 ;
  assign n10089 = x113 & n878 ;
  assign n10090 = n10088 | n10089 ;
  assign n10091 = x112 & n959 ;
  assign n10092 = n10090 | n10091 ;
  assign n10093 = ( ~x17 & n10086 ) | ( ~x17 & n10092 ) | ( n10086 & n10092 ) ;
  assign n10094 = x17 & ~n10092 ;
  assign n10095 = ( ~n10087 & n10093 ) | ( ~n10087 & n10094 ) | ( n10093 & n10094 ) ;
  assign n10096 = ( n9818 & ~n10085 ) | ( n9818 & n10095 ) | ( ~n10085 & n10095 ) ;
  assign n10097 = ( n9818 & n10085 ) | ( n9818 & n10095 ) | ( n10085 & n10095 ) ;
  assign n10098 = ( n10085 & n10096 ) | ( n10085 & ~n10097 ) | ( n10096 & ~n10097 ) ;
  assign n10099 = ( n9832 & n9887 ) | ( n9832 & n10098 ) | ( n9887 & n10098 ) ;
  assign n10100 = ( ~n9832 & n9887 ) | ( ~n9832 & n10098 ) | ( n9887 & n10098 ) ;
  assign n10101 = ( n9832 & ~n10099 ) | ( n9832 & n10100 ) | ( ~n10099 & n10100 ) ;
  assign n10102 = n301 & n8461 ;
  assign n10103 = x8 & n10102 ;
  assign n10104 = x123 & n309 ;
  assign n10105 = x122 & n306 ;
  assign n10106 = n10104 | n10105 ;
  assign n10107 = x121 & n359 ;
  assign n10108 = n10106 | n10107 ;
  assign n10109 = ( ~x8 & n10102 ) | ( ~x8 & n10108 ) | ( n10102 & n10108 ) ;
  assign n10110 = x8 & ~n10108 ;
  assign n10111 = ( ~n10103 & n10109 ) | ( ~n10103 & n10110 ) | ( n10109 & n10110 ) ;
  assign n10112 = n449 & n7444 ;
  assign n10113 = x11 & n10112 ;
  assign n10114 = x120 & n456 ;
  assign n10115 = x119 & n453 ;
  assign n10116 = n10114 | n10115 ;
  assign n10117 = x118 & n536 ;
  assign n10118 = n10116 | n10117 ;
  assign n10119 = ( ~x11 & n10112 ) | ( ~x11 & n10118 ) | ( n10112 & n10118 ) ;
  assign n10120 = x11 & ~n10118 ;
  assign n10121 = ( ~n10113 & n10119 ) | ( ~n10113 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10122 = ( ~n10101 & n10111 ) | ( ~n10101 & n10121 ) | ( n10111 & n10121 ) ;
  assign n10123 = ( n10101 & n10111 ) | ( n10101 & n10121 ) | ( n10111 & n10121 ) ;
  assign n10124 = ( n10101 & n10122 ) | ( n10101 & ~n10123 ) | ( n10122 & ~n10123 ) ;
  assign n10125 = n206 & n9038 ;
  assign n10126 = x5 & n10125 ;
  assign n10127 = x126 & n205 ;
  assign n10128 = x125 & n201 ;
  assign n10129 = n10127 | n10128 ;
  assign n10130 = x124 & n221 ;
  assign n10131 = n10129 | n10130 ;
  assign n10132 = ( ~x5 & n10125 ) | ( ~x5 & n10131 ) | ( n10125 & n10131 ) ;
  assign n10133 = x5 & ~n10131 ;
  assign n10134 = ( ~n10126 & n10132 ) | ( ~n10126 & n10133 ) | ( n10132 & n10133 ) ;
  assign n10135 = ( n9834 & n10124 ) | ( n9834 & n10134 ) | ( n10124 & n10134 ) ;
  assign n10136 = ( ~n9834 & n10124 ) | ( ~n9834 & n10134 ) | ( n10124 & n10134 ) ;
  assign n10137 = ( n9834 & ~n10135 ) | ( n9834 & n10136 ) | ( ~n10135 & n10136 ) ;
  assign n10138 = x0 & x1 ;
  assign n10139 = n9865 & n10138 ;
  assign n10140 = ( ~x0 & x127 ) | ( ~x0 & n9865 ) | ( x127 & n9865 ) ;
  assign n10141 = ( x2 & n144 ) | ( x2 & ~n10140 ) | ( n144 & ~n10140 ) ;
  assign n10142 = n10139 | n10141 ;
  assign n10143 = ( n9857 & ~n10137 ) | ( n9857 & n10142 ) | ( ~n10137 & n10142 ) ;
  assign n10144 = ( n9857 & n10137 ) | ( n9857 & n10142 ) | ( n10137 & n10142 ) ;
  assign n10145 = ( n10137 & n10143 ) | ( n10137 & ~n10144 ) | ( n10143 & ~n10144 ) ;
  assign n10146 = ( n9873 & ~n9875 ) | ( n9873 & n10145 ) | ( ~n9875 & n10145 ) ;
  assign n10147 = ( n9873 & n9875 ) | ( n9873 & n10145 ) | ( n9875 & n10145 ) ;
  assign n10148 = ( n9875 & n10146 ) | ( n9875 & ~n10147 ) | ( n10146 & ~n10147 ) ;
  assign n10149 = n206 & n9576 ;
  assign n10150 = x5 & n10149 ;
  assign n10151 = x127 & n205 ;
  assign n10152 = x126 & n201 ;
  assign n10153 = n10151 | n10152 ;
  assign n10154 = x125 & n221 ;
  assign n10155 = n10153 | n10154 ;
  assign n10156 = ( ~x5 & n10149 ) | ( ~x5 & n10155 ) | ( n10149 & n10155 ) ;
  assign n10157 = x5 & ~n10155 ;
  assign n10158 = ( ~n10150 & n10156 ) | ( ~n10150 & n10157 ) | ( n10156 & n10157 ) ;
  assign n10159 = n449 & n7696 ;
  assign n10160 = x11 & n10159 ;
  assign n10161 = x121 & n456 ;
  assign n10162 = x120 & n453 ;
  assign n10163 = n10161 | n10162 ;
  assign n10164 = x119 & n536 ;
  assign n10165 = n10163 | n10164 ;
  assign n10166 = ( ~x11 & n10159 ) | ( ~x11 & n10165 ) | ( n10159 & n10165 ) ;
  assign n10167 = x11 & ~n10165 ;
  assign n10168 = ( ~n10160 & n10166 ) | ( ~n10160 & n10167 ) | ( n10166 & n10167 ) ;
  assign n10169 = n649 & n6940 ;
  assign n10170 = x14 & n10169 ;
  assign n10171 = x118 & n656 ;
  assign n10172 = x117 & n653 ;
  assign n10173 = n10171 | n10172 ;
  assign n10174 = x116 & n744 ;
  assign n10175 = n10173 | n10174 ;
  assign n10176 = ( ~x14 & n10169 ) | ( ~x14 & n10175 ) | ( n10169 & n10175 ) ;
  assign n10177 = x14 & ~n10175 ;
  assign n10178 = ( ~n10170 & n10176 ) | ( ~n10170 & n10177 ) | ( n10176 & n10177 ) ;
  assign n10179 = n874 & n6446 ;
  assign n10180 = x17 & n10179 ;
  assign n10181 = x115 & n881 ;
  assign n10182 = x114 & n878 ;
  assign n10183 = n10181 | n10182 ;
  assign n10184 = x113 & n959 ;
  assign n10185 = n10183 | n10184 ;
  assign n10186 = ( ~x17 & n10179 ) | ( ~x17 & n10185 ) | ( n10179 & n10185 ) ;
  assign n10187 = x17 & ~n10185 ;
  assign n10188 = ( ~n10180 & n10186 ) | ( ~n10180 & n10187 ) | ( n10186 & n10187 ) ;
  assign n10189 = n1427 & n4930 ;
  assign n10190 = x23 & n10189 ;
  assign n10191 = x109 & n1434 ;
  assign n10192 = x108 & n1431 ;
  assign n10193 = n10191 | n10192 ;
  assign n10194 = x107 & n1531 ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = ( ~x23 & n10189 ) | ( ~x23 & n10195 ) | ( n10189 & n10195 ) ;
  assign n10197 = x23 & ~n10195 ;
  assign n10198 = ( ~n10190 & n10196 ) | ( ~n10190 & n10197 ) | ( n10196 & n10197 ) ;
  assign n10199 = n1755 & n4331 ;
  assign n10200 = x26 & n10199 ;
  assign n10201 = x106 & n1762 ;
  assign n10202 = x105 & n1759 ;
  assign n10203 = n10201 | n10202 ;
  assign n10204 = x104 & n1895 ;
  assign n10205 = n10203 | n10204 ;
  assign n10206 = ( ~x26 & n10199 ) | ( ~x26 & n10205 ) | ( n10199 & n10205 ) ;
  assign n10207 = x26 & ~n10205 ;
  assign n10208 = ( ~n10200 & n10206 ) | ( ~n10200 & n10207 ) | ( n10206 & n10207 ) ;
  assign n10209 = n2545 & n3264 ;
  assign n10210 = x32 & n10209 ;
  assign n10211 = x100 & n2552 ;
  assign n10212 = x99 & n2549 ;
  assign n10213 = n10211 | n10212 ;
  assign n10214 = x98 & n2696 ;
  assign n10215 = n10213 | n10214 ;
  assign n10216 = ( ~x32 & n10209 ) | ( ~x32 & n10215 ) | ( n10209 & n10215 ) ;
  assign n10217 = x32 & ~n10215 ;
  assign n10218 = ( ~n10210 & n10216 ) | ( ~n10210 & n10217 ) | ( n10216 & n10217 ) ;
  assign n10219 = n2788 & n2982 ;
  assign n10220 = x35 & n10219 ;
  assign n10221 = x97 & n2989 ;
  assign n10222 = x96 & n2986 ;
  assign n10223 = n10221 | n10222 ;
  assign n10224 = x95 & n3159 ;
  assign n10225 = n10223 | n10224 ;
  assign n10226 = ( ~x35 & n10219 ) | ( ~x35 & n10225 ) | ( n10219 & n10225 ) ;
  assign n10227 = x35 & ~n10225 ;
  assign n10228 = ( ~n10220 & n10226 ) | ( ~n10220 & n10227 ) | ( n10226 & n10227 ) ;
  assign n10229 = n2476 & n3492 ;
  assign n10230 = x38 & n10229 ;
  assign n10231 = x94 & n3499 ;
  assign n10232 = x93 & n3496 ;
  assign n10233 = n10231 | n10232 ;
  assign n10234 = x92 & n3662 ;
  assign n10235 = n10233 | n10234 ;
  assign n10236 = ( ~x38 & n10229 ) | ( ~x38 & n10235 ) | ( n10229 & n10235 ) ;
  assign n10237 = x38 & ~n10235 ;
  assign n10238 = ( ~n10230 & n10236 ) | ( ~n10230 & n10237 ) | ( n10236 & n10237 ) ;
  assign n10239 = n1959 & n4020 ;
  assign n10240 = x41 & n10239 ;
  assign n10241 = x91 & n4027 ;
  assign n10242 = x90 & n4024 ;
  assign n10243 = n10241 | n10242 ;
  assign n10244 = x89 & n4223 ;
  assign n10245 = n10243 | n10244 ;
  assign n10246 = ( ~x41 & n10239 ) | ( ~x41 & n10245 ) | ( n10239 & n10245 ) ;
  assign n10247 = x41 & ~n10245 ;
  assign n10248 = ( ~n10240 & n10246 ) | ( ~n10240 & n10247 ) | ( n10246 & n10247 ) ;
  assign n10249 = n1368 & n5223 ;
  assign n10250 = x47 & n10249 ;
  assign n10251 = x85 & n5230 ;
  assign n10252 = x84 & n5227 ;
  assign n10253 = n10251 | n10252 ;
  assign n10254 = x83 & n5434 ;
  assign n10255 = n10253 | n10254 ;
  assign n10256 = ( ~x47 & n10249 ) | ( ~x47 & n10255 ) | ( n10249 & n10255 ) ;
  assign n10257 = x47 & ~n10255 ;
  assign n10258 = ( ~n10250 & n10256 ) | ( ~n10250 & n10257 ) | ( n10256 & n10257 ) ;
  assign n10259 = n1006 & n5858 ;
  assign n10260 = x50 & n10259 ;
  assign n10261 = x82 & n5865 ;
  assign n10262 = x81 & n5862 ;
  assign n10263 = n10261 | n10262 ;
  assign n10264 = x80 & n6092 ;
  assign n10265 = n10263 | n10264 ;
  assign n10266 = ( ~x50 & n10259 ) | ( ~x50 & n10265 ) | ( n10259 & n10265 ) ;
  assign n10267 = x50 & ~n10265 ;
  assign n10268 = ( ~n10260 & n10266 ) | ( ~n10260 & n10267 ) | ( n10266 & n10267 ) ;
  assign n10269 = n823 & n6546 ;
  assign n10270 = x53 & n10269 ;
  assign n10271 = x79 & n6553 ;
  assign n10272 = x78 & n6550 ;
  assign n10273 = n10271 | n10272 ;
  assign n10274 = x77 & n6787 ;
  assign n10275 = n10273 | n10274 ;
  assign n10276 = ( ~x53 & n10269 ) | ( ~x53 & n10275 ) | ( n10269 & n10275 ) ;
  assign n10277 = x53 & ~n10275 ;
  assign n10278 = ( ~n10270 & n10276 ) | ( ~n10270 & n10277 ) | ( n10276 & n10277 ) ;
  assign n10279 = n565 & n7277 ;
  assign n10280 = x56 & n10279 ;
  assign n10281 = x76 & n7545 ;
  assign n10282 = x75 & n7273 ;
  assign n10283 = n10281 | n10282 ;
  assign n10284 = x74 & n7552 ;
  assign n10285 = n10283 | n10284 ;
  assign n10286 = ( ~x56 & n10279 ) | ( ~x56 & n10285 ) | ( n10279 & n10285 ) ;
  assign n10287 = x56 & ~n10285 ;
  assign n10288 = ( ~n10280 & n10286 ) | ( ~n10280 & n10287 ) | ( n10286 & n10287 ) ;
  assign n10289 = n388 & n8067 ;
  assign n10290 = x59 & n10289 ;
  assign n10291 = x73 & n8074 ;
  assign n10292 = x72 & n8071 ;
  assign n10293 = n10291 | n10292 ;
  assign n10294 = x71 & n8298 ;
  assign n10295 = n10293 | n10294 ;
  assign n10296 = ( ~x59 & n10289 ) | ( ~x59 & n10295 ) | ( n10289 & n10295 ) ;
  assign n10297 = x59 & ~n10295 ;
  assign n10298 = ( ~n10290 & n10296 ) | ( ~n10290 & n10297 ) | ( n10296 & n10297 ) ;
  assign n10299 = ( x62 & x63 ) | ( x62 & x67 ) | ( x63 & x67 ) ;
  assign n10300 = ( x62 & x66 ) | ( x62 & ~n9394 ) | ( x66 & ~n9394 ) ;
  assign n10301 = ( x66 & n10299 ) | ( x66 & ~n10300 ) | ( n10299 & ~n10300 ) ;
  assign n10302 = n276 & n8859 ;
  assign n10303 = x62 & n10302 ;
  assign n10304 = x70 & n8866 ;
  assign n10305 = x69 & n8863 ;
  assign n10306 = n10304 | n10305 ;
  assign n10307 = x68 & n9125 ;
  assign n10308 = n10306 | n10307 ;
  assign n10309 = ( ~x62 & n10302 ) | ( ~x62 & n10308 ) | ( n10302 & n10308 ) ;
  assign n10310 = x62 & ~n10308 ;
  assign n10311 = ( ~n10303 & n10309 ) | ( ~n10303 & n10310 ) | ( n10309 & n10310 ) ;
  assign n10312 = ( x2 & ~n10301 ) | ( x2 & n10311 ) | ( ~n10301 & n10311 ) ;
  assign n10313 = ( x2 & n10301 ) | ( x2 & n10311 ) | ( n10301 & n10311 ) ;
  assign n10314 = ( n10301 & n10312 ) | ( n10301 & ~n10313 ) | ( n10312 & ~n10313 ) ;
  assign n10315 = ( n9981 & n10298 ) | ( n9981 & n10314 ) | ( n10298 & n10314 ) ;
  assign n10316 = ( ~n9981 & n10298 ) | ( ~n9981 & n10314 ) | ( n10298 & n10314 ) ;
  assign n10317 = ( n9981 & ~n10315 ) | ( n9981 & n10316 ) | ( ~n10315 & n10316 ) ;
  assign n10318 = ( ~n9995 & n10288 ) | ( ~n9995 & n10317 ) | ( n10288 & n10317 ) ;
  assign n10319 = ( n9995 & n10288 ) | ( n9995 & n10317 ) | ( n10288 & n10317 ) ;
  assign n10320 = ( n9995 & n10318 ) | ( n9995 & ~n10319 ) | ( n10318 & ~n10319 ) ;
  assign n10321 = ( n9997 & n10278 ) | ( n9997 & n10320 ) | ( n10278 & n10320 ) ;
  assign n10322 = ( ~n9997 & n10278 ) | ( ~n9997 & n10320 ) | ( n10278 & n10320 ) ;
  assign n10323 = ( n9997 & ~n10321 ) | ( n9997 & n10322 ) | ( ~n10321 & n10322 ) ;
  assign n10324 = ( n10000 & n10268 ) | ( n10000 & n10323 ) | ( n10268 & n10323 ) ;
  assign n10325 = ( ~n10000 & n10268 ) | ( ~n10000 & n10323 ) | ( n10268 & n10323 ) ;
  assign n10326 = ( n10000 & ~n10324 ) | ( n10000 & n10325 ) | ( ~n10324 & n10325 ) ;
  assign n10327 = ( n10014 & n10258 ) | ( n10014 & n10326 ) | ( n10258 & n10326 ) ;
  assign n10328 = ( ~n10014 & n10258 ) | ( ~n10014 & n10326 ) | ( n10258 & n10326 ) ;
  assign n10329 = ( n10014 & ~n10327 ) | ( n10014 & n10328 ) | ( ~n10327 & n10328 ) ;
  assign n10330 = n1602 & n4625 ;
  assign n10331 = x44 & n10330 ;
  assign n10332 = x88 & n4791 ;
  assign n10333 = x87 & n4621 ;
  assign n10334 = n10332 | n10333 ;
  assign n10335 = x86 & n4795 ;
  assign n10336 = n10334 | n10335 ;
  assign n10337 = ( ~x44 & n10330 ) | ( ~x44 & n10336 ) | ( n10330 & n10336 ) ;
  assign n10338 = x44 & ~n10336 ;
  assign n10339 = ( ~n10331 & n10337 ) | ( ~n10331 & n10338 ) | ( n10337 & n10338 ) ;
  assign n10340 = ( n10016 & n10329 ) | ( n10016 & n10339 ) | ( n10329 & n10339 ) ;
  assign n10341 = ( ~n10016 & n10329 ) | ( ~n10016 & n10339 ) | ( n10329 & n10339 ) ;
  assign n10342 = ( n10016 & ~n10340 ) | ( n10016 & n10341 ) | ( ~n10340 & n10341 ) ;
  assign n10343 = ( n10019 & n10248 ) | ( n10019 & n10342 ) | ( n10248 & n10342 ) ;
  assign n10344 = ( ~n10019 & n10248 ) | ( ~n10019 & n10342 ) | ( n10248 & n10342 ) ;
  assign n10345 = ( n10019 & ~n10343 ) | ( n10019 & n10344 ) | ( ~n10343 & n10344 ) ;
  assign n10346 = ( n10033 & n10238 ) | ( n10033 & n10345 ) | ( n10238 & n10345 ) ;
  assign n10347 = ( ~n10033 & n10238 ) | ( ~n10033 & n10345 ) | ( n10238 & n10345 ) ;
  assign n10348 = ( n10033 & ~n10346 ) | ( n10033 & n10347 ) | ( ~n10346 & n10347 ) ;
  assign n10349 = ( n10036 & n10228 ) | ( n10036 & n10348 ) | ( n10228 & n10348 ) ;
  assign n10350 = ( ~n10036 & n10228 ) | ( ~n10036 & n10348 ) | ( n10228 & n10348 ) ;
  assign n10351 = ( n10036 & ~n10349 ) | ( n10036 & n10350 ) | ( ~n10349 & n10350 ) ;
  assign n10352 = ( n10038 & n10218 ) | ( n10038 & n10351 ) | ( n10218 & n10351 ) ;
  assign n10353 = ( ~n10038 & n10218 ) | ( ~n10038 & n10351 ) | ( n10218 & n10351 ) ;
  assign n10354 = ( n10038 & ~n10352 ) | ( n10038 & n10353 ) | ( ~n10352 & n10353 ) ;
  assign n10355 = n2137 & n3941 ;
  assign n10356 = x29 & n10355 ;
  assign n10357 = x103 & n2144 ;
  assign n10358 = x102 & n2141 ;
  assign n10359 = n10357 | n10358 ;
  assign n10360 = x101 & n2267 ;
  assign n10361 = n10359 | n10360 ;
  assign n10362 = ( ~x29 & n10355 ) | ( ~x29 & n10361 ) | ( n10355 & n10361 ) ;
  assign n10363 = x29 & ~n10361 ;
  assign n10364 = ( ~n10356 & n10362 ) | ( ~n10356 & n10363 ) | ( n10362 & n10363 ) ;
  assign n10365 = ( n10052 & n10354 ) | ( n10052 & n10364 ) | ( n10354 & n10364 ) ;
  assign n10366 = ( ~n10052 & n10354 ) | ( ~n10052 & n10364 ) | ( n10354 & n10364 ) ;
  assign n10367 = ( n10052 & ~n10365 ) | ( n10052 & n10366 ) | ( ~n10365 & n10366 ) ;
  assign n10368 = ( n10054 & n10208 ) | ( n10054 & n10367 ) | ( n10208 & n10367 ) ;
  assign n10369 = ( ~n10054 & n10208 ) | ( ~n10054 & n10367 ) | ( n10208 & n10367 ) ;
  assign n10370 = ( n10054 & ~n10368 ) | ( n10054 & n10369 ) | ( ~n10368 & n10369 ) ;
  assign n10371 = ( n10067 & n10198 ) | ( n10067 & n10370 ) | ( n10198 & n10370 ) ;
  assign n10372 = ( ~n10067 & n10198 ) | ( ~n10067 & n10370 ) | ( n10198 & n10370 ) ;
  assign n10373 = ( n10067 & ~n10371 ) | ( n10067 & n10372 ) | ( ~n10371 & n10372 ) ;
  assign n10374 = n1146 & n5558 ;
  assign n10375 = x20 & n10374 ;
  assign n10376 = x112 & n1153 ;
  assign n10377 = x111 & n1150 ;
  assign n10378 = n10376 | n10377 ;
  assign n10379 = x110 & n1217 ;
  assign n10380 = n10378 | n10379 ;
  assign n10381 = ( ~x20 & n10374 ) | ( ~x20 & n10380 ) | ( n10374 & n10380 ) ;
  assign n10382 = x20 & ~n10380 ;
  assign n10383 = ( ~n10375 & n10381 ) | ( ~n10375 & n10382 ) | ( n10381 & n10382 ) ;
  assign n10384 = ( n10081 & n10373 ) | ( n10081 & n10383 ) | ( n10373 & n10383 ) ;
  assign n10385 = ( ~n10081 & n10373 ) | ( ~n10081 & n10383 ) | ( n10373 & n10383 ) ;
  assign n10386 = ( n10081 & ~n10384 ) | ( n10081 & n10385 ) | ( ~n10384 & n10385 ) ;
  assign n10387 = ( n10083 & n10188 ) | ( n10083 & n10386 ) | ( n10188 & n10386 ) ;
  assign n10388 = ( ~n10083 & n10188 ) | ( ~n10083 & n10386 ) | ( n10188 & n10386 ) ;
  assign n10389 = ( n10083 & ~n10387 ) | ( n10083 & n10388 ) | ( ~n10387 & n10388 ) ;
  assign n10390 = ( n10097 & n10178 ) | ( n10097 & n10389 ) | ( n10178 & n10389 ) ;
  assign n10391 = ( ~n10097 & n10178 ) | ( ~n10097 & n10389 ) | ( n10178 & n10389 ) ;
  assign n10392 = ( n10097 & ~n10390 ) | ( n10097 & n10391 ) | ( ~n10390 & n10391 ) ;
  assign n10393 = ( n10099 & n10168 ) | ( n10099 & n10392 ) | ( n10168 & n10392 ) ;
  assign n10394 = ( ~n10099 & n10168 ) | ( ~n10099 & n10392 ) | ( n10168 & n10392 ) ;
  assign n10395 = ( n10099 & ~n10393 ) | ( n10099 & n10394 ) | ( ~n10393 & n10394 ) ;
  assign n10396 = n301 & n8729 ;
  assign n10397 = x8 & n10396 ;
  assign n10398 = x124 & n309 ;
  assign n10399 = x123 & n306 ;
  assign n10400 = n10398 | n10399 ;
  assign n10401 = x122 & n359 ;
  assign n10402 = n10400 | n10401 ;
  assign n10403 = ( ~x8 & n10396 ) | ( ~x8 & n10402 ) | ( n10396 & n10402 ) ;
  assign n10404 = x8 & ~n10402 ;
  assign n10405 = ( ~n10397 & n10403 ) | ( ~n10397 & n10404 ) | ( n10403 & n10404 ) ;
  assign n10406 = ( n10123 & n10395 ) | ( n10123 & n10405 ) | ( n10395 & n10405 ) ;
  assign n10407 = ( ~n10123 & n10395 ) | ( ~n10123 & n10405 ) | ( n10395 & n10405 ) ;
  assign n10408 = ( n10123 & ~n10406 ) | ( n10123 & n10407 ) | ( ~n10406 & n10407 ) ;
  assign n10409 = ( n10135 & n10158 ) | ( n10135 & n10408 ) | ( n10158 & n10408 ) ;
  assign n10410 = ( ~n10135 & n10158 ) | ( ~n10135 & n10408 ) | ( n10158 & n10408 ) ;
  assign n10411 = ( n10135 & ~n10409 ) | ( n10135 & n10410 ) | ( ~n10409 & n10410 ) ;
  assign n10412 = ( n10144 & ~n10147 ) | ( n10144 & n10411 ) | ( ~n10147 & n10411 ) ;
  assign n10413 = ( n10144 & n10147 ) | ( n10144 & n10411 ) | ( n10147 & n10411 ) ;
  assign n10414 = ( n10147 & n10412 ) | ( n10147 & ~n10413 ) | ( n10412 & ~n10413 ) ;
  assign n10415 = n301 & n9009 ;
  assign n10416 = x8 & n10415 ;
  assign n10417 = x125 & n309 ;
  assign n10418 = x124 & n306 ;
  assign n10419 = n10417 | n10418 ;
  assign n10420 = x123 & n359 ;
  assign n10421 = n10419 | n10420 ;
  assign n10422 = ( ~x8 & n10415 ) | ( ~x8 & n10421 ) | ( n10415 & n10421 ) ;
  assign n10423 = x8 & ~n10421 ;
  assign n10424 = ( ~n10416 & n10422 ) | ( ~n10416 & n10423 ) | ( n10422 & n10423 ) ;
  assign n10425 = n449 & n8207 ;
  assign n10426 = x11 & n10425 ;
  assign n10427 = x122 & n456 ;
  assign n10428 = x121 & n453 ;
  assign n10429 = n10427 | n10428 ;
  assign n10430 = x120 & n536 ;
  assign n10431 = n10429 | n10430 ;
  assign n10432 = ( ~x11 & n10425 ) | ( ~x11 & n10431 ) | ( n10425 & n10431 ) ;
  assign n10433 = x11 & ~n10431 ;
  assign n10434 = ( ~n10426 & n10432 ) | ( ~n10426 & n10433 ) | ( n10432 & n10433 ) ;
  assign n10435 = n649 & n7181 ;
  assign n10436 = x14 & n10435 ;
  assign n10437 = x119 & n656 ;
  assign n10438 = x118 & n653 ;
  assign n10439 = n10437 | n10438 ;
  assign n10440 = x117 & n744 ;
  assign n10441 = n10439 | n10440 ;
  assign n10442 = ( ~x14 & n10435 ) | ( ~x14 & n10441 ) | ( n10435 & n10441 ) ;
  assign n10443 = x14 & ~n10441 ;
  assign n10444 = ( ~n10436 & n10442 ) | ( ~n10436 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10445 = n874 & n6462 ;
  assign n10446 = x17 & n10445 ;
  assign n10447 = x116 & n881 ;
  assign n10448 = x115 & n878 ;
  assign n10449 = n10447 | n10448 ;
  assign n10450 = x114 & n959 ;
  assign n10451 = n10449 | n10450 ;
  assign n10452 = ( ~x17 & n10445 ) | ( ~x17 & n10451 ) | ( n10445 & n10451 ) ;
  assign n10453 = x17 & ~n10451 ;
  assign n10454 = ( ~n10446 & n10452 ) | ( ~n10446 & n10453 ) | ( n10452 & n10453 ) ;
  assign n10455 = n1146 & n5774 ;
  assign n10456 = x20 & n10455 ;
  assign n10457 = x113 & n1153 ;
  assign n10458 = x112 & n1150 ;
  assign n10459 = n10457 | n10458 ;
  assign n10460 = x111 & n1217 ;
  assign n10461 = n10459 | n10460 ;
  assign n10462 = ( ~x20 & n10455 ) | ( ~x20 & n10461 ) | ( n10455 & n10461 ) ;
  assign n10463 = x20 & ~n10461 ;
  assign n10464 = ( ~n10456 & n10462 ) | ( ~n10456 & n10463 ) | ( n10462 & n10463 ) ;
  assign n10465 = n1427 & n5331 ;
  assign n10466 = x23 & n10465 ;
  assign n10467 = x110 & n1434 ;
  assign n10468 = x109 & n1431 ;
  assign n10469 = n10467 | n10468 ;
  assign n10470 = x108 & n1531 ;
  assign n10471 = n10469 | n10470 ;
  assign n10472 = ( ~x23 & n10465 ) | ( ~x23 & n10471 ) | ( n10465 & n10471 ) ;
  assign n10473 = x23 & ~n10471 ;
  assign n10474 = ( ~n10466 & n10472 ) | ( ~n10466 & n10473 ) | ( n10472 & n10473 ) ;
  assign n10475 = n1755 & n4523 ;
  assign n10476 = x26 & n10475 ;
  assign n10477 = x107 & n1762 ;
  assign n10478 = x106 & n1759 ;
  assign n10479 = n10477 | n10478 ;
  assign n10480 = x105 & n1895 ;
  assign n10481 = n10479 | n10480 ;
  assign n10482 = ( ~x26 & n10475 ) | ( ~x26 & n10481 ) | ( n10475 & n10481 ) ;
  assign n10483 = x26 & ~n10481 ;
  assign n10484 = ( ~n10476 & n10482 ) | ( ~n10476 & n10483 ) | ( n10482 & n10483 ) ;
  assign n10485 = n2137 & n3957 ;
  assign n10486 = x29 & n10485 ;
  assign n10487 = x104 & n2144 ;
  assign n10488 = x103 & n2141 ;
  assign n10489 = n10487 | n10488 ;
  assign n10490 = x102 & n2267 ;
  assign n10491 = n10489 | n10490 ;
  assign n10492 = ( ~x29 & n10485 ) | ( ~x29 & n10491 ) | ( n10485 & n10491 ) ;
  assign n10493 = x29 & ~n10491 ;
  assign n10494 = ( ~n10486 & n10492 ) | ( ~n10486 & n10493 ) | ( n10492 & n10493 ) ;
  assign n10495 = n2939 & n2982 ;
  assign n10496 = x35 & n10495 ;
  assign n10497 = x98 & n2989 ;
  assign n10498 = x97 & n2986 ;
  assign n10499 = n10497 | n10498 ;
  assign n10500 = x96 & n3159 ;
  assign n10501 = n10499 | n10500 ;
  assign n10502 = ( ~x35 & n10495 ) | ( ~x35 & n10501 ) | ( n10495 & n10501 ) ;
  assign n10503 = x35 & ~n10501 ;
  assign n10504 = ( ~n10496 & n10502 ) | ( ~n10496 & n10503 ) | ( n10502 & n10503 ) ;
  assign n10505 = n1822 & n4625 ;
  assign n10506 = x44 & n10505 ;
  assign n10507 = x89 & n4791 ;
  assign n10508 = x88 & n4621 ;
  assign n10509 = n10507 | n10508 ;
  assign n10510 = x87 & n4795 ;
  assign n10511 = n10509 | n10510 ;
  assign n10512 = ( ~x44 & n10505 ) | ( ~x44 & n10511 ) | ( n10505 & n10511 ) ;
  assign n10513 = x44 & ~n10511 ;
  assign n10514 = ( ~n10506 & n10512 ) | ( ~n10506 & n10513 ) | ( n10512 & n10513 ) ;
  assign n10515 = n1384 & n5223 ;
  assign n10516 = x47 & n10515 ;
  assign n10517 = x86 & n5230 ;
  assign n10518 = x85 & n5227 ;
  assign n10519 = n10517 | n10518 ;
  assign n10520 = x84 & n5434 ;
  assign n10521 = n10519 | n10520 ;
  assign n10522 = ( ~x47 & n10515 ) | ( ~x47 & n10521 ) | ( n10515 & n10521 ) ;
  assign n10523 = x47 & ~n10521 ;
  assign n10524 = ( ~n10516 & n10522 ) | ( ~n10516 & n10523 ) | ( n10522 & n10523 ) ;
  assign n10525 = n1093 & n5858 ;
  assign n10526 = x50 & n10525 ;
  assign n10527 = x83 & n5865 ;
  assign n10528 = x82 & n5862 ;
  assign n10529 = n10527 | n10528 ;
  assign n10530 = x81 & n6092 ;
  assign n10531 = n10529 | n10530 ;
  assign n10532 = ( ~x50 & n10525 ) | ( ~x50 & n10531 ) | ( n10525 & n10531 ) ;
  assign n10533 = x50 & ~n10531 ;
  assign n10534 = ( ~n10526 & n10532 ) | ( ~n10526 & n10533 ) | ( n10532 & n10533 ) ;
  assign n10535 = n840 & n6546 ;
  assign n10536 = x53 & n10535 ;
  assign n10537 = x80 & n6553 ;
  assign n10538 = x79 & n6550 ;
  assign n10539 = n10537 | n10538 ;
  assign n10540 = x78 & n6787 ;
  assign n10541 = n10539 | n10540 ;
  assign n10542 = ( ~x53 & n10535 ) | ( ~x53 & n10541 ) | ( n10535 & n10541 ) ;
  assign n10543 = x53 & ~n10541 ;
  assign n10544 = ( ~n10536 & n10542 ) | ( ~n10536 & n10543 ) | ( n10542 & n10543 ) ;
  assign n10545 = n436 & n8067 ;
  assign n10546 = x59 & n10545 ;
  assign n10547 = x74 & n8074 ;
  assign n10548 = x73 & n8071 ;
  assign n10549 = n10547 | n10548 ;
  assign n10550 = x72 & n8298 ;
  assign n10551 = n10549 | n10550 ;
  assign n10552 = ( ~x59 & n10545 ) | ( ~x59 & n10551 ) | ( n10545 & n10551 ) ;
  assign n10553 = x59 & ~n10551 ;
  assign n10554 = ( ~n10546 & n10552 ) | ( ~n10546 & n10553 ) | ( n10552 & n10553 ) ;
  assign n10555 = n322 & n8859 ;
  assign n10556 = x62 & n10555 ;
  assign n10557 = x71 & n8866 ;
  assign n10558 = x70 & n8863 ;
  assign n10559 = n10557 | n10558 ;
  assign n10560 = x69 & n9125 ;
  assign n10561 = n10559 | n10560 ;
  assign n10562 = ( ~x62 & n10555 ) | ( ~x62 & n10561 ) | ( n10555 & n10561 ) ;
  assign n10563 = x62 & ~n10561 ;
  assign n10564 = ( ~n10556 & n10562 ) | ( ~n10556 & n10563 ) | ( n10562 & n10563 ) ;
  assign n10565 = ( x62 & x63 ) | ( x62 & x68 ) | ( x63 & x68 ) ;
  assign n10566 = ( x62 & x67 ) | ( x62 & ~n9394 ) | ( x67 & ~n9394 ) ;
  assign n10567 = ( x67 & n10565 ) | ( x67 & ~n10566 ) | ( n10565 & ~n10566 ) ;
  assign n10568 = ( x2 & n10564 ) | ( x2 & n10567 ) | ( n10564 & n10567 ) ;
  assign n10569 = ( ~x2 & n10564 ) | ( ~x2 & n10567 ) | ( n10564 & n10567 ) ;
  assign n10570 = ( x2 & ~n10568 ) | ( x2 & n10569 ) | ( ~n10568 & n10569 ) ;
  assign n10571 = ( n10313 & n10554 ) | ( n10313 & n10570 ) | ( n10554 & n10570 ) ;
  assign n10572 = ( n10313 & ~n10554 ) | ( n10313 & n10570 ) | ( ~n10554 & n10570 ) ;
  assign n10573 = ( n10554 & ~n10571 ) | ( n10554 & n10572 ) | ( ~n10571 & n10572 ) ;
  assign n10574 = n626 & n7277 ;
  assign n10575 = x56 & n10574 ;
  assign n10576 = x77 & n7545 ;
  assign n10577 = x76 & n7273 ;
  assign n10578 = n10576 | n10577 ;
  assign n10579 = x75 & n7552 ;
  assign n10580 = n10578 | n10579 ;
  assign n10581 = ( ~x56 & n10574 ) | ( ~x56 & n10580 ) | ( n10574 & n10580 ) ;
  assign n10582 = x56 & ~n10580 ;
  assign n10583 = ( ~n10575 & n10581 ) | ( ~n10575 & n10582 ) | ( n10581 & n10582 ) ;
  assign n10584 = ( n10315 & ~n10573 ) | ( n10315 & n10583 ) | ( ~n10573 & n10583 ) ;
  assign n10585 = ( n10315 & n10573 ) | ( n10315 & n10583 ) | ( n10573 & n10583 ) ;
  assign n10586 = ( n10573 & n10584 ) | ( n10573 & ~n10585 ) | ( n10584 & ~n10585 ) ;
  assign n10587 = ( ~n10319 & n10544 ) | ( ~n10319 & n10586 ) | ( n10544 & n10586 ) ;
  assign n10588 = ( n10319 & n10544 ) | ( n10319 & n10586 ) | ( n10544 & n10586 ) ;
  assign n10589 = ( n10319 & n10587 ) | ( n10319 & ~n10588 ) | ( n10587 & ~n10588 ) ;
  assign n10590 = ( n10321 & ~n10534 ) | ( n10321 & n10589 ) | ( ~n10534 & n10589 ) ;
  assign n10591 = ( n10321 & n10534 ) | ( n10321 & n10589 ) | ( n10534 & n10589 ) ;
  assign n10592 = ( n10534 & n10590 ) | ( n10534 & ~n10591 ) | ( n10590 & ~n10591 ) ;
  assign n10593 = ( n10324 & ~n10524 ) | ( n10324 & n10592 ) | ( ~n10524 & n10592 ) ;
  assign n10594 = ( n10324 & n10524 ) | ( n10324 & n10592 ) | ( n10524 & n10592 ) ;
  assign n10595 = ( n10524 & n10593 ) | ( n10524 & ~n10594 ) | ( n10593 & ~n10594 ) ;
  assign n10596 = ( n10327 & n10514 ) | ( n10327 & n10595 ) | ( n10514 & n10595 ) ;
  assign n10597 = ( ~n10327 & n10514 ) | ( ~n10327 & n10595 ) | ( n10514 & n10595 ) ;
  assign n10598 = ( n10327 & ~n10596 ) | ( n10327 & n10597 ) | ( ~n10596 & n10597 ) ;
  assign n10599 = n2083 & n4020 ;
  assign n10600 = x41 & n10599 ;
  assign n10601 = x92 & n4027 ;
  assign n10602 = x91 & n4024 ;
  assign n10603 = n10601 | n10602 ;
  assign n10604 = x90 & n4223 ;
  assign n10605 = n10603 | n10604 ;
  assign n10606 = ( ~x41 & n10599 ) | ( ~x41 & n10605 ) | ( n10599 & n10605 ) ;
  assign n10607 = x41 & ~n10605 ;
  assign n10608 = ( ~n10600 & n10606 ) | ( ~n10600 & n10607 ) | ( n10606 & n10607 ) ;
  assign n10609 = ( n10340 & n10598 ) | ( n10340 & n10608 ) | ( n10598 & n10608 ) ;
  assign n10610 = ( ~n10340 & n10598 ) | ( ~n10340 & n10608 ) | ( n10598 & n10608 ) ;
  assign n10611 = ( n10340 & ~n10609 ) | ( n10340 & n10610 ) | ( ~n10609 & n10610 ) ;
  assign n10612 = n2492 & n3492 ;
  assign n10613 = x38 & n10612 ;
  assign n10614 = x95 & n3499 ;
  assign n10615 = x94 & n3496 ;
  assign n10616 = n10614 | n10615 ;
  assign n10617 = x93 & n3662 ;
  assign n10618 = n10616 | n10617 ;
  assign n10619 = ( ~x38 & n10612 ) | ( ~x38 & n10618 ) | ( n10612 & n10618 ) ;
  assign n10620 = x38 & ~n10618 ;
  assign n10621 = ( ~n10613 & n10619 ) | ( ~n10613 & n10620 ) | ( n10619 & n10620 ) ;
  assign n10622 = ( n10343 & ~n10611 ) | ( n10343 & n10621 ) | ( ~n10611 & n10621 ) ;
  assign n10623 = ( n10343 & n10611 ) | ( n10343 & n10621 ) | ( n10611 & n10621 ) ;
  assign n10624 = ( n10611 & n10622 ) | ( n10611 & ~n10623 ) | ( n10622 & ~n10623 ) ;
  assign n10625 = ( ~n10346 & n10504 ) | ( ~n10346 & n10624 ) | ( n10504 & n10624 ) ;
  assign n10626 = ( n10346 & n10504 ) | ( n10346 & n10624 ) | ( n10504 & n10624 ) ;
  assign n10627 = ( n10346 & n10625 ) | ( n10346 & ~n10626 ) | ( n10625 & ~n10626 ) ;
  assign n10628 = n2545 & n3591 ;
  assign n10629 = x32 & n10628 ;
  assign n10630 = x101 & n2552 ;
  assign n10631 = x100 & n2549 ;
  assign n10632 = n10630 | n10631 ;
  assign n10633 = x99 & n2696 ;
  assign n10634 = n10632 | n10633 ;
  assign n10635 = ( ~x32 & n10628 ) | ( ~x32 & n10634 ) | ( n10628 & n10634 ) ;
  assign n10636 = x32 & ~n10634 ;
  assign n10637 = ( ~n10629 & n10635 ) | ( ~n10629 & n10636 ) | ( n10635 & n10636 ) ;
  assign n10638 = ( n10349 & ~n10627 ) | ( n10349 & n10637 ) | ( ~n10627 & n10637 ) ;
  assign n10639 = ( n10349 & n10627 ) | ( n10349 & n10637 ) | ( n10627 & n10637 ) ;
  assign n10640 = ( n10627 & n10638 ) | ( n10627 & ~n10639 ) | ( n10638 & ~n10639 ) ;
  assign n10641 = ( n10352 & ~n10494 ) | ( n10352 & n10640 ) | ( ~n10494 & n10640 ) ;
  assign n10642 = ( n10352 & n10494 ) | ( n10352 & n10640 ) | ( n10494 & n10640 ) ;
  assign n10643 = ( n10494 & n10641 ) | ( n10494 & ~n10642 ) | ( n10641 & ~n10642 ) ;
  assign n10644 = ( n10365 & n10484 ) | ( n10365 & n10643 ) | ( n10484 & n10643 ) ;
  assign n10645 = ( ~n10365 & n10484 ) | ( ~n10365 & n10643 ) | ( n10484 & n10643 ) ;
  assign n10646 = ( n10365 & ~n10644 ) | ( n10365 & n10645 ) | ( ~n10644 & n10645 ) ;
  assign n10647 = ( n10368 & ~n10474 ) | ( n10368 & n10646 ) | ( ~n10474 & n10646 ) ;
  assign n10648 = ( n10368 & n10474 ) | ( n10368 & n10646 ) | ( n10474 & n10646 ) ;
  assign n10649 = ( n10474 & n10647 ) | ( n10474 & ~n10648 ) | ( n10647 & ~n10648 ) ;
  assign n10650 = ( n10371 & ~n10464 ) | ( n10371 & n10649 ) | ( ~n10464 & n10649 ) ;
  assign n10651 = ( n10371 & n10464 ) | ( n10371 & n10649 ) | ( n10464 & n10649 ) ;
  assign n10652 = ( n10464 & n10650 ) | ( n10464 & ~n10651 ) | ( n10650 & ~n10651 ) ;
  assign n10653 = ( n10384 & ~n10454 ) | ( n10384 & n10652 ) | ( ~n10454 & n10652 ) ;
  assign n10654 = ( n10384 & n10454 ) | ( n10384 & n10652 ) | ( n10454 & n10652 ) ;
  assign n10655 = ( n10454 & n10653 ) | ( n10454 & ~n10654 ) | ( n10653 & ~n10654 ) ;
  assign n10656 = ( n10387 & ~n10444 ) | ( n10387 & n10655 ) | ( ~n10444 & n10655 ) ;
  assign n10657 = ( n10387 & n10444 ) | ( n10387 & n10655 ) | ( n10444 & n10655 ) ;
  assign n10658 = ( n10444 & n10656 ) | ( n10444 & ~n10657 ) | ( n10656 & ~n10657 ) ;
  assign n10659 = ( n10390 & ~n10434 ) | ( n10390 & n10658 ) | ( ~n10434 & n10658 ) ;
  assign n10660 = ( n10390 & n10434 ) | ( n10390 & n10658 ) | ( n10434 & n10658 ) ;
  assign n10661 = ( n10434 & n10659 ) | ( n10434 & ~n10660 ) | ( n10659 & ~n10660 ) ;
  assign n10662 = ( n10393 & n10424 ) | ( n10393 & n10661 ) | ( n10424 & n10661 ) ;
  assign n10663 = ( ~n10393 & n10424 ) | ( ~n10393 & n10661 ) | ( n10424 & n10661 ) ;
  assign n10664 = ( n10393 & ~n10662 ) | ( n10393 & n10663 ) | ( ~n10662 & n10663 ) ;
  assign n10665 = x127 & n201 ;
  assign n10666 = n206 | n10665 ;
  assign n10667 = ( n9867 & n10665 ) | ( n9867 & n10666 ) | ( n10665 & n10666 ) ;
  assign n10668 = x126 & n221 ;
  assign n10669 = ( ~x5 & n10667 ) | ( ~x5 & n10668 ) | ( n10667 & n10668 ) ;
  assign n10670 = ( x5 & ~n10667 ) | ( x5 & n10668 ) | ( ~n10667 & n10668 ) ;
  assign n10671 = ~n10668 & n10670 ;
  assign n10672 = n10669 | n10671 ;
  assign n10673 = ( n10406 & n10664 ) | ( n10406 & n10672 ) | ( n10664 & n10672 ) ;
  assign n10674 = ( n10406 & ~n10664 ) | ( n10406 & n10672 ) | ( ~n10664 & n10672 ) ;
  assign n10675 = ( n10664 & ~n10673 ) | ( n10664 & n10674 ) | ( ~n10673 & n10674 ) ;
  assign n10676 = ( n10409 & ~n10413 ) | ( n10409 & n10675 ) | ( ~n10413 & n10675 ) ;
  assign n10677 = ( n10409 & n10413 ) | ( n10409 & n10675 ) | ( n10413 & n10675 ) ;
  assign n10678 = ( n10413 & n10676 ) | ( n10413 & ~n10677 ) | ( n10676 & ~n10677 ) ;
  assign n10679 = x127 & n221 ;
  assign n10680 = n206 | n10679 ;
  assign n10681 = ( n9865 & n10679 ) | ( n9865 & n10680 ) | ( n10679 & n10680 ) ;
  assign n10682 = x5 & ~n10681 ;
  assign n10683 = ~x5 & n10681 ;
  assign n10684 = n10682 | n10683 ;
  assign n10685 = n301 & n9038 ;
  assign n10686 = x8 & n10685 ;
  assign n10687 = x126 & n309 ;
  assign n10688 = x125 & n306 ;
  assign n10689 = n10687 | n10688 ;
  assign n10690 = x124 & n359 ;
  assign n10691 = n10689 | n10690 ;
  assign n10692 = ( ~x8 & n10685 ) | ( ~x8 & n10691 ) | ( n10685 & n10691 ) ;
  assign n10693 = x8 & ~n10691 ;
  assign n10694 = ( ~n10686 & n10692 ) | ( ~n10686 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10695 = n449 & n8461 ;
  assign n10696 = x11 & n10695 ;
  assign n10697 = x123 & n456 ;
  assign n10698 = x122 & n453 ;
  assign n10699 = n10697 | n10698 ;
  assign n10700 = x121 & n536 ;
  assign n10701 = n10699 | n10700 ;
  assign n10702 = ( ~x11 & n10695 ) | ( ~x11 & n10701 ) | ( n10695 & n10701 ) ;
  assign n10703 = x11 & ~n10701 ;
  assign n10704 = ( ~n10696 & n10702 ) | ( ~n10696 & n10703 ) | ( n10702 & n10703 ) ;
  assign n10705 = n649 & n7444 ;
  assign n10706 = x14 & n10705 ;
  assign n10707 = x120 & n656 ;
  assign n10708 = x119 & n653 ;
  assign n10709 = n10707 | n10708 ;
  assign n10710 = x118 & n744 ;
  assign n10711 = n10709 | n10710 ;
  assign n10712 = ( ~x14 & n10705 ) | ( ~x14 & n10711 ) | ( n10705 & n10711 ) ;
  assign n10713 = x14 & ~n10711 ;
  assign n10714 = ( ~n10706 & n10712 ) | ( ~n10706 & n10713 ) | ( n10712 & n10713 ) ;
  assign n10715 = n874 & n6924 ;
  assign n10716 = x17 & n10715 ;
  assign n10717 = x117 & n881 ;
  assign n10718 = x116 & n878 ;
  assign n10719 = n10717 | n10718 ;
  assign n10720 = x115 & n959 ;
  assign n10721 = n10719 | n10720 ;
  assign n10722 = ( ~x17 & n10715 ) | ( ~x17 & n10721 ) | ( n10715 & n10721 ) ;
  assign n10723 = x17 & ~n10721 ;
  assign n10724 = ( ~n10716 & n10722 ) | ( ~n10716 & n10723 ) | ( n10722 & n10723 ) ;
  assign n10725 = n1146 & n6002 ;
  assign n10726 = x20 & n10725 ;
  assign n10727 = x114 & n1153 ;
  assign n10728 = x113 & n1150 ;
  assign n10729 = n10727 | n10728 ;
  assign n10730 = x112 & n1217 ;
  assign n10731 = n10729 | n10730 ;
  assign n10732 = ( ~x20 & n10725 ) | ( ~x20 & n10731 ) | ( n10725 & n10731 ) ;
  assign n10733 = x20 & ~n10731 ;
  assign n10734 = ( ~n10726 & n10732 ) | ( ~n10726 & n10733 ) | ( n10732 & n10733 ) ;
  assign n10735 = n1427 & n5347 ;
  assign n10736 = x23 & n10735 ;
  assign n10737 = x111 & n1434 ;
  assign n10738 = x110 & n1431 ;
  assign n10739 = n10737 | n10738 ;
  assign n10740 = x109 & n1531 ;
  assign n10741 = n10739 | n10740 ;
  assign n10742 = ( ~x23 & n10735 ) | ( ~x23 & n10741 ) | ( n10735 & n10741 ) ;
  assign n10743 = x23 & ~n10741 ;
  assign n10744 = ( ~n10736 & n10742 ) | ( ~n10736 & n10743 ) | ( n10742 & n10743 ) ;
  assign n10745 = n1755 & n4914 ;
  assign n10746 = x26 & n10745 ;
  assign n10747 = x108 & n1762 ;
  assign n10748 = x107 & n1759 ;
  assign n10749 = n10747 | n10748 ;
  assign n10750 = x106 & n1895 ;
  assign n10751 = n10749 | n10750 ;
  assign n10752 = ( ~x26 & n10745 ) | ( ~x26 & n10751 ) | ( n10745 & n10751 ) ;
  assign n10753 = x26 & ~n10751 ;
  assign n10754 = ( ~n10746 & n10752 ) | ( ~n10746 & n10753 ) | ( n10752 & n10753 ) ;
  assign n10755 = n2137 & n4145 ;
  assign n10756 = x29 & n10755 ;
  assign n10757 = x105 & n2144 ;
  assign n10758 = x104 & n2141 ;
  assign n10759 = n10757 | n10758 ;
  assign n10760 = x103 & n2267 ;
  assign n10761 = n10759 | n10760 ;
  assign n10762 = ( ~x29 & n10755 ) | ( ~x29 & n10761 ) | ( n10755 & n10761 ) ;
  assign n10763 = x29 & ~n10761 ;
  assign n10764 = ( ~n10756 & n10762 ) | ( ~n10756 & n10763 ) | ( n10762 & n10763 ) ;
  assign n10765 = n2545 & n3764 ;
  assign n10766 = x32 & n10765 ;
  assign n10767 = x102 & n2552 ;
  assign n10768 = x101 & n2549 ;
  assign n10769 = n10767 | n10768 ;
  assign n10770 = x100 & n2696 ;
  assign n10771 = n10769 | n10770 ;
  assign n10772 = ( ~x32 & n10765 ) | ( ~x32 & n10771 ) | ( n10765 & n10771 ) ;
  assign n10773 = x32 & ~n10771 ;
  assign n10774 = ( ~n10766 & n10772 ) | ( ~n10766 & n10773 ) | ( n10772 & n10773 ) ;
  assign n10775 = n2982 & n3248 ;
  assign n10776 = x35 & n10775 ;
  assign n10777 = x99 & n2989 ;
  assign n10778 = x98 & n2986 ;
  assign n10779 = n10777 | n10778 ;
  assign n10780 = x97 & n3159 ;
  assign n10781 = n10779 | n10780 ;
  assign n10782 = ( ~x35 & n10775 ) | ( ~x35 & n10781 ) | ( n10775 & n10781 ) ;
  assign n10783 = x35 & ~n10781 ;
  assign n10784 = ( ~n10776 & n10782 ) | ( ~n10776 & n10783 ) | ( n10782 & n10783 ) ;
  assign n10785 = n2772 & n3492 ;
  assign n10786 = x38 & n10785 ;
  assign n10787 = x96 & n3499 ;
  assign n10788 = x95 & n3496 ;
  assign n10789 = n10787 | n10788 ;
  assign n10790 = x94 & n3662 ;
  assign n10791 = n10789 | n10790 ;
  assign n10792 = ( ~x38 & n10785 ) | ( ~x38 & n10791 ) | ( n10785 & n10791 ) ;
  assign n10793 = x38 & ~n10791 ;
  assign n10794 = ( ~n10786 & n10792 ) | ( ~n10786 & n10793 ) | ( n10792 & n10793 ) ;
  assign n10795 = n2220 & n4020 ;
  assign n10796 = x41 & n10795 ;
  assign n10797 = x93 & n4027 ;
  assign n10798 = x92 & n4024 ;
  assign n10799 = n10797 | n10798 ;
  assign n10800 = x91 & n4223 ;
  assign n10801 = n10799 | n10800 ;
  assign n10802 = ( ~x41 & n10795 ) | ( ~x41 & n10801 ) | ( n10795 & n10801 ) ;
  assign n10803 = x41 & ~n10801 ;
  assign n10804 = ( ~n10796 & n10802 ) | ( ~n10796 & n10803 ) | ( n10802 & n10803 ) ;
  assign n10805 = n1838 & n4625 ;
  assign n10806 = x44 & n10805 ;
  assign n10807 = x90 & n4791 ;
  assign n10808 = x89 & n4621 ;
  assign n10809 = n10807 | n10808 ;
  assign n10810 = x88 & n4795 ;
  assign n10811 = n10809 | n10810 ;
  assign n10812 = ( ~x44 & n10805 ) | ( ~x44 & n10811 ) | ( n10805 & n10811 ) ;
  assign n10813 = x44 & ~n10811 ;
  assign n10814 = ( ~n10806 & n10812 ) | ( ~n10806 & n10813 ) | ( n10812 & n10813 ) ;
  assign n10815 = x86 & n5227 ;
  assign n10816 = x85 | n10815 ;
  assign n10817 = ( n5434 & n10815 ) | ( n5434 & n10816 ) | ( n10815 & n10816 ) ;
  assign n10818 = n1494 & n5223 ;
  assign n10819 = n10817 | n10818 ;
  assign n10820 = x87 & n5230 ;
  assign n10821 = ( ~x47 & n10819 ) | ( ~x47 & n10820 ) | ( n10819 & n10820 ) ;
  assign n10822 = ( x47 & ~n10819 ) | ( x47 & n10820 ) | ( ~n10819 & n10820 ) ;
  assign n10823 = ~n10820 & n10822 ;
  assign n10824 = n10821 | n10823 ;
  assign n10825 = n1190 & n5858 ;
  assign n10826 = x50 & n10825 ;
  assign n10827 = x84 & n5865 ;
  assign n10828 = x83 & n5862 ;
  assign n10829 = n10827 | n10828 ;
  assign n10830 = x82 & n6092 ;
  assign n10831 = n10829 | n10830 ;
  assign n10832 = ( ~x50 & n10825 ) | ( ~x50 & n10831 ) | ( n10825 & n10831 ) ;
  assign n10833 = x50 & ~n10831 ;
  assign n10834 = ( ~n10826 & n10832 ) | ( ~n10826 & n10833 ) | ( n10832 & n10833 ) ;
  assign n10835 = n990 & n6546 ;
  assign n10836 = x53 & n10835 ;
  assign n10837 = x81 & n6553 ;
  assign n10838 = x80 & n6550 ;
  assign n10839 = n10837 | n10838 ;
  assign n10840 = x79 & n6787 ;
  assign n10841 = n10839 | n10840 ;
  assign n10842 = ( ~x53 & n10835 ) | ( ~x53 & n10841 ) | ( n10835 & n10841 ) ;
  assign n10843 = x53 & ~n10841 ;
  assign n10844 = ( ~n10836 & n10842 ) | ( ~n10836 & n10843 ) | ( n10842 & n10843 ) ;
  assign n10845 = n508 & n8067 ;
  assign n10846 = x59 & n10845 ;
  assign n10847 = x75 & n8074 ;
  assign n10848 = x74 & n8071 ;
  assign n10849 = n10847 | n10848 ;
  assign n10850 = x73 & n8298 ;
  assign n10851 = n10849 | n10850 ;
  assign n10852 = ( ~x59 & n10845 ) | ( ~x59 & n10851 ) | ( n10845 & n10851 ) ;
  assign n10853 = x59 & ~n10851 ;
  assign n10854 = ( ~n10846 & n10852 ) | ( ~n10846 & n10853 ) | ( n10852 & n10853 ) ;
  assign n10855 = n372 & n8859 ;
  assign n10856 = x62 & n10855 ;
  assign n10857 = x72 & n8866 ;
  assign n10858 = x71 & n8863 ;
  assign n10859 = n10857 | n10858 ;
  assign n10860 = x70 & n9125 ;
  assign n10861 = n10859 | n10860 ;
  assign n10862 = ( ~x62 & n10855 ) | ( ~x62 & n10861 ) | ( n10855 & n10861 ) ;
  assign n10863 = x62 & ~n10861 ;
  assign n10864 = ( ~n10856 & n10862 ) | ( ~n10856 & n10863 ) | ( n10862 & n10863 ) ;
  assign n10865 = ( x62 & x63 ) | ( x62 & x69 ) | ( x63 & x69 ) ;
  assign n10866 = ( x62 & x68 ) | ( x62 & ~n9394 ) | ( x68 & ~n9394 ) ;
  assign n10867 = ( x68 & n10865 ) | ( x68 & ~n10866 ) | ( n10865 & ~n10866 ) ;
  assign n10868 = ( x2 & n10864 ) | ( x2 & n10867 ) | ( n10864 & n10867 ) ;
  assign n10869 = ( ~x2 & n10864 ) | ( ~x2 & n10867 ) | ( n10864 & n10867 ) ;
  assign n10870 = ( x2 & ~n10868 ) | ( x2 & n10869 ) | ( ~n10868 & n10869 ) ;
  assign n10871 = ( n10568 & n10854 ) | ( n10568 & n10870 ) | ( n10854 & n10870 ) ;
  assign n10872 = ( n10568 & ~n10854 ) | ( n10568 & n10870 ) | ( ~n10854 & n10870 ) ;
  assign n10873 = ( n10854 & ~n10871 ) | ( n10854 & n10872 ) | ( ~n10871 & n10872 ) ;
  assign n10874 = n697 & n7277 ;
  assign n10875 = x56 & n10874 ;
  assign n10876 = x78 & n7545 ;
  assign n10877 = x77 & n7273 ;
  assign n10878 = n10876 | n10877 ;
  assign n10879 = x76 & n7552 ;
  assign n10880 = n10878 | n10879 ;
  assign n10881 = ( ~x56 & n10874 ) | ( ~x56 & n10880 ) | ( n10874 & n10880 ) ;
  assign n10882 = x56 & ~n10880 ;
  assign n10883 = ( ~n10875 & n10881 ) | ( ~n10875 & n10882 ) | ( n10881 & n10882 ) ;
  assign n10884 = ( n10571 & ~n10873 ) | ( n10571 & n10883 ) | ( ~n10873 & n10883 ) ;
  assign n10885 = ( n10571 & n10873 ) | ( n10571 & n10883 ) | ( n10873 & n10883 ) ;
  assign n10886 = ( n10873 & n10884 ) | ( n10873 & ~n10885 ) | ( n10884 & ~n10885 ) ;
  assign n10887 = ( n10585 & n10844 ) | ( n10585 & n10886 ) | ( n10844 & n10886 ) ;
  assign n10888 = ( n10585 & ~n10844 ) | ( n10585 & n10886 ) | ( ~n10844 & n10886 ) ;
  assign n10889 = ( n10844 & ~n10887 ) | ( n10844 & n10888 ) | ( ~n10887 & n10888 ) ;
  assign n10890 = ( n10588 & n10834 ) | ( n10588 & n10889 ) | ( n10834 & n10889 ) ;
  assign n10891 = ( n10588 & ~n10834 ) | ( n10588 & n10889 ) | ( ~n10834 & n10889 ) ;
  assign n10892 = ( n10834 & ~n10890 ) | ( n10834 & n10891 ) | ( ~n10890 & n10891 ) ;
  assign n10893 = ( n10591 & n10824 ) | ( n10591 & n10892 ) | ( n10824 & n10892 ) ;
  assign n10894 = ( n10591 & ~n10824 ) | ( n10591 & n10892 ) | ( ~n10824 & n10892 ) ;
  assign n10895 = ( n10824 & ~n10893 ) | ( n10824 & n10894 ) | ( ~n10893 & n10894 ) ;
  assign n10896 = ( n10594 & n10814 ) | ( n10594 & n10895 ) | ( n10814 & n10895 ) ;
  assign n10897 = ( n10594 & ~n10814 ) | ( n10594 & n10895 ) | ( ~n10814 & n10895 ) ;
  assign n10898 = ( n10814 & ~n10896 ) | ( n10814 & n10897 ) | ( ~n10896 & n10897 ) ;
  assign n10899 = ( n10596 & ~n10804 ) | ( n10596 & n10898 ) | ( ~n10804 & n10898 ) ;
  assign n10900 = ( n10596 & n10804 ) | ( n10596 & n10898 ) | ( n10804 & n10898 ) ;
  assign n10901 = ( n10804 & n10899 ) | ( n10804 & ~n10900 ) | ( n10899 & ~n10900 ) ;
  assign n10902 = ( n10609 & n10794 ) | ( n10609 & n10901 ) | ( n10794 & n10901 ) ;
  assign n10903 = ( n10609 & ~n10794 ) | ( n10609 & n10901 ) | ( ~n10794 & n10901 ) ;
  assign n10904 = ( n10794 & ~n10902 ) | ( n10794 & n10903 ) | ( ~n10902 & n10903 ) ;
  assign n10905 = ( n10623 & ~n10784 ) | ( n10623 & n10904 ) | ( ~n10784 & n10904 ) ;
  assign n10906 = ( n10623 & n10784 ) | ( n10623 & n10904 ) | ( n10784 & n10904 ) ;
  assign n10907 = ( n10784 & n10905 ) | ( n10784 & ~n10906 ) | ( n10905 & ~n10906 ) ;
  assign n10908 = ( n10626 & ~n10774 ) | ( n10626 & n10907 ) | ( ~n10774 & n10907 ) ;
  assign n10909 = ( n10626 & n10774 ) | ( n10626 & n10907 ) | ( n10774 & n10907 ) ;
  assign n10910 = ( n10774 & n10908 ) | ( n10774 & ~n10909 ) | ( n10908 & ~n10909 ) ;
  assign n10911 = ( n10639 & n10764 ) | ( n10639 & n10910 ) | ( n10764 & n10910 ) ;
  assign n10912 = ( n10639 & ~n10764 ) | ( n10639 & n10910 ) | ( ~n10764 & n10910 ) ;
  assign n10913 = ( n10764 & ~n10911 ) | ( n10764 & n10912 ) | ( ~n10911 & n10912 ) ;
  assign n10914 = ( n10642 & ~n10754 ) | ( n10642 & n10913 ) | ( ~n10754 & n10913 ) ;
  assign n10915 = ( n10642 & n10754 ) | ( n10642 & n10913 ) | ( n10754 & n10913 ) ;
  assign n10916 = ( n10754 & n10914 ) | ( n10754 & ~n10915 ) | ( n10914 & ~n10915 ) ;
  assign n10917 = ( n10644 & n10744 ) | ( n10644 & n10916 ) | ( n10744 & n10916 ) ;
  assign n10918 = ( n10644 & ~n10744 ) | ( n10644 & n10916 ) | ( ~n10744 & n10916 ) ;
  assign n10919 = ( n10744 & ~n10917 ) | ( n10744 & n10918 ) | ( ~n10917 & n10918 ) ;
  assign n10920 = ( n10648 & n10734 ) | ( n10648 & n10919 ) | ( n10734 & n10919 ) ;
  assign n10921 = ( n10648 & ~n10734 ) | ( n10648 & n10919 ) | ( ~n10734 & n10919 ) ;
  assign n10922 = ( n10734 & ~n10920 ) | ( n10734 & n10921 ) | ( ~n10920 & n10921 ) ;
  assign n10923 = ( n10651 & n10724 ) | ( n10651 & n10922 ) | ( n10724 & n10922 ) ;
  assign n10924 = ( n10651 & ~n10724 ) | ( n10651 & n10922 ) | ( ~n10724 & n10922 ) ;
  assign n10925 = ( n10724 & ~n10923 ) | ( n10724 & n10924 ) | ( ~n10923 & n10924 ) ;
  assign n10926 = ( n10654 & n10714 ) | ( n10654 & n10925 ) | ( n10714 & n10925 ) ;
  assign n10927 = ( n10654 & ~n10714 ) | ( n10654 & n10925 ) | ( ~n10714 & n10925 ) ;
  assign n10928 = ( n10714 & ~n10926 ) | ( n10714 & n10927 ) | ( ~n10926 & n10927 ) ;
  assign n10929 = ( n10657 & n10704 ) | ( n10657 & n10928 ) | ( n10704 & n10928 ) ;
  assign n10930 = ( n10657 & ~n10704 ) | ( n10657 & n10928 ) | ( ~n10704 & n10928 ) ;
  assign n10931 = ( n10704 & ~n10929 ) | ( n10704 & n10930 ) | ( ~n10929 & n10930 ) ;
  assign n10932 = ( n10660 & n10694 ) | ( n10660 & n10931 ) | ( n10694 & n10931 ) ;
  assign n10933 = ( n10660 & ~n10694 ) | ( n10660 & n10931 ) | ( ~n10694 & n10931 ) ;
  assign n10934 = ( n10694 & ~n10932 ) | ( n10694 & n10933 ) | ( ~n10932 & n10933 ) ;
  assign n10935 = ( n10662 & ~n10684 ) | ( n10662 & n10934 ) | ( ~n10684 & n10934 ) ;
  assign n10936 = ( n10662 & n10684 ) | ( n10662 & n10934 ) | ( n10684 & n10934 ) ;
  assign n10937 = ( n10684 & n10935 ) | ( n10684 & ~n10936 ) | ( n10935 & ~n10936 ) ;
  assign n10938 = ( n10673 & ~n10677 ) | ( n10673 & n10937 ) | ( ~n10677 & n10937 ) ;
  assign n10939 = ( n10673 & n10677 ) | ( n10673 & n10937 ) | ( n10677 & n10937 ) ;
  assign n10940 = ( n10677 & n10938 ) | ( n10677 & ~n10939 ) | ( n10938 & ~n10939 ) ;
  assign n10941 = n301 & n9576 ;
  assign n10942 = x8 & n10941 ;
  assign n10943 = x127 & n309 ;
  assign n10944 = x126 & n306 ;
  assign n10945 = n10943 | n10944 ;
  assign n10946 = x125 & n359 ;
  assign n10947 = n10945 | n10946 ;
  assign n10948 = ( ~x8 & n10941 ) | ( ~x8 & n10947 ) | ( n10941 & n10947 ) ;
  assign n10949 = x8 & ~n10947 ;
  assign n10950 = ( ~n10942 & n10948 ) | ( ~n10942 & n10949 ) | ( n10948 & n10949 ) ;
  assign n10951 = n449 & n8729 ;
  assign n10952 = x11 & n10951 ;
  assign n10953 = x123 & n453 ;
  assign n10954 = x122 & n536 ;
  assign n10955 = n10953 | n10954 ;
  assign n10956 = x124 & n456 ;
  assign n10957 = n10955 | n10956 ;
  assign n10958 = ( ~x11 & n10951 ) | ( ~x11 & n10957 ) | ( n10951 & n10957 ) ;
  assign n10959 = x11 & ~n10957 ;
  assign n10960 = ( ~n10952 & n10958 ) | ( ~n10952 & n10959 ) | ( n10958 & n10959 ) ;
  assign n10961 = n649 & n7696 ;
  assign n10962 = x14 & n10961 ;
  assign n10963 = x121 & n656 ;
  assign n10964 = x120 & n653 ;
  assign n10965 = n10963 | n10964 ;
  assign n10966 = x119 & n744 ;
  assign n10967 = n10965 | n10966 ;
  assign n10968 = ( ~x14 & n10961 ) | ( ~x14 & n10967 ) | ( n10961 & n10967 ) ;
  assign n10969 = x14 & ~n10967 ;
  assign n10970 = ( ~n10962 & n10968 ) | ( ~n10962 & n10969 ) | ( n10968 & n10969 ) ;
  assign n10971 = n874 & n6940 ;
  assign n10972 = x17 & n10971 ;
  assign n10973 = x118 & n881 ;
  assign n10974 = x117 & n878 ;
  assign n10975 = n10973 | n10974 ;
  assign n10976 = x116 & n959 ;
  assign n10977 = n10975 | n10976 ;
  assign n10978 = ( ~x17 & n10971 ) | ( ~x17 & n10977 ) | ( n10971 & n10977 ) ;
  assign n10979 = x17 & ~n10977 ;
  assign n10980 = ( ~n10972 & n10978 ) | ( ~n10972 & n10979 ) | ( n10978 & n10979 ) ;
  assign n10981 = n1146 & n6446 ;
  assign n10982 = x20 & n10981 ;
  assign n10983 = x115 & n1153 ;
  assign n10984 = x114 & n1150 ;
  assign n10985 = n10983 | n10984 ;
  assign n10986 = x113 & n1217 ;
  assign n10987 = n10985 | n10986 ;
  assign n10988 = ( ~x20 & n10981 ) | ( ~x20 & n10987 ) | ( n10981 & n10987 ) ;
  assign n10989 = x20 & ~n10987 ;
  assign n10990 = ( ~n10982 & n10988 ) | ( ~n10982 & n10989 ) | ( n10988 & n10989 ) ;
  assign n10991 = n1427 & n5558 ;
  assign n10992 = x23 & n10991 ;
  assign n10993 = x112 & n1434 ;
  assign n10994 = x111 & n1431 ;
  assign n10995 = n10993 | n10994 ;
  assign n10996 = x110 & n1531 ;
  assign n10997 = n10995 | n10996 ;
  assign n10998 = ( ~x23 & n10991 ) | ( ~x23 & n10997 ) | ( n10991 & n10997 ) ;
  assign n10999 = x23 & ~n10997 ;
  assign n11000 = ( ~n10992 & n10998 ) | ( ~n10992 & n10999 ) | ( n10998 & n10999 ) ;
  assign n11001 = n1755 & n4930 ;
  assign n11002 = x26 & n11001 ;
  assign n11003 = x109 & n1762 ;
  assign n11004 = x108 & n1759 ;
  assign n11005 = n11003 | n11004 ;
  assign n11006 = x107 & n1895 ;
  assign n11007 = n11005 | n11006 ;
  assign n11008 = ( ~x26 & n11001 ) | ( ~x26 & n11007 ) | ( n11001 & n11007 ) ;
  assign n11009 = x26 & ~n11007 ;
  assign n11010 = ( ~n11002 & n11008 ) | ( ~n11002 & n11009 ) | ( n11008 & n11009 ) ;
  assign n11011 = n2137 & n4331 ;
  assign n11012 = x29 & n11011 ;
  assign n11013 = x106 & n2144 ;
  assign n11014 = x105 & n2141 ;
  assign n11015 = n11013 | n11014 ;
  assign n11016 = x104 & n2267 ;
  assign n11017 = n11015 | n11016 ;
  assign n11018 = ( ~x29 & n11011 ) | ( ~x29 & n11017 ) | ( n11011 & n11017 ) ;
  assign n11019 = x29 & ~n11017 ;
  assign n11020 = ( ~n11012 & n11018 ) | ( ~n11012 & n11019 ) | ( n11018 & n11019 ) ;
  assign n11021 = n2545 & n3941 ;
  assign n11022 = x32 & n11021 ;
  assign n11023 = x103 & n2552 ;
  assign n11024 = x102 & n2549 ;
  assign n11025 = n11023 | n11024 ;
  assign n11026 = x101 & n2696 ;
  assign n11027 = n11025 | n11026 ;
  assign n11028 = ( ~x32 & n11021 ) | ( ~x32 & n11027 ) | ( n11021 & n11027 ) ;
  assign n11029 = x32 & ~n11027 ;
  assign n11030 = ( ~n11022 & n11028 ) | ( ~n11022 & n11029 ) | ( n11028 & n11029 ) ;
  assign n11031 = n2982 & n3264 ;
  assign n11032 = x35 & n11031 ;
  assign n11033 = x100 & n2989 ;
  assign n11034 = x99 & n2986 ;
  assign n11035 = n11033 | n11034 ;
  assign n11036 = x98 & n3159 ;
  assign n11037 = n11035 | n11036 ;
  assign n11038 = ( ~x35 & n11031 ) | ( ~x35 & n11037 ) | ( n11031 & n11037 ) ;
  assign n11039 = x35 & ~n11037 ;
  assign n11040 = ( ~n11032 & n11038 ) | ( ~n11032 & n11039 ) | ( n11038 & n11039 ) ;
  assign n11041 = n2788 & n3492 ;
  assign n11042 = x38 & n11041 ;
  assign n11043 = x97 & n3499 ;
  assign n11044 = x96 & n3496 ;
  assign n11045 = n11043 | n11044 ;
  assign n11046 = x95 & n3662 ;
  assign n11047 = n11045 | n11046 ;
  assign n11048 = ( ~x38 & n11041 ) | ( ~x38 & n11047 ) | ( n11041 & n11047 ) ;
  assign n11049 = x38 & ~n11047 ;
  assign n11050 = ( ~n11042 & n11048 ) | ( ~n11042 & n11049 ) | ( n11048 & n11049 ) ;
  assign n11051 = n2476 & n4020 ;
  assign n11052 = x41 & n11051 ;
  assign n11053 = x94 & n4027 ;
  assign n11054 = x93 & n4024 ;
  assign n11055 = n11053 | n11054 ;
  assign n11056 = x92 & n4223 ;
  assign n11057 = n11055 | n11056 ;
  assign n11058 = ( ~x41 & n11051 ) | ( ~x41 & n11057 ) | ( n11051 & n11057 ) ;
  assign n11059 = x41 & ~n11057 ;
  assign n11060 = ( ~n11052 & n11058 ) | ( ~n11052 & n11059 ) | ( n11058 & n11059 ) ;
  assign n11061 = n1602 & n5223 ;
  assign n11062 = x47 & n11061 ;
  assign n11063 = x88 & n5230 ;
  assign n11064 = x87 & n5227 ;
  assign n11065 = n11063 | n11064 ;
  assign n11066 = x86 & n5434 ;
  assign n11067 = n11065 | n11066 ;
  assign n11068 = ( ~x47 & n11061 ) | ( ~x47 & n11067 ) | ( n11061 & n11067 ) ;
  assign n11069 = x47 & ~n11067 ;
  assign n11070 = ( ~n11062 & n11068 ) | ( ~n11062 & n11069 ) | ( n11068 & n11069 ) ;
  assign n11071 = n1368 & n5858 ;
  assign n11072 = x50 & n11071 ;
  assign n11073 = x85 & n5865 ;
  assign n11074 = x84 & n5862 ;
  assign n11075 = n11073 | n11074 ;
  assign n11076 = x83 & n6092 ;
  assign n11077 = n11075 | n11076 ;
  assign n11078 = ( ~x50 & n11071 ) | ( ~x50 & n11077 ) | ( n11071 & n11077 ) ;
  assign n11079 = x50 & ~n11077 ;
  assign n11080 = ( ~n11072 & n11078 ) | ( ~n11072 & n11079 ) | ( n11078 & n11079 ) ;
  assign n11081 = n1006 & n6546 ;
  assign n11082 = x53 & n11081 ;
  assign n11083 = x82 & n6553 ;
  assign n11084 = x81 & n6550 ;
  assign n11085 = n11083 | n11084 ;
  assign n11086 = x80 & n6787 ;
  assign n11087 = n11085 | n11086 ;
  assign n11088 = ( ~x53 & n11081 ) | ( ~x53 & n11087 ) | ( n11081 & n11087 ) ;
  assign n11089 = x53 & ~n11087 ;
  assign n11090 = ( ~n11082 & n11088 ) | ( ~n11082 & n11089 ) | ( n11088 & n11089 ) ;
  assign n11091 = n823 & n7277 ;
  assign n11092 = x56 & n11091 ;
  assign n11093 = x79 & n7545 ;
  assign n11094 = x78 & n7273 ;
  assign n11095 = n11093 | n11094 ;
  assign n11096 = x77 & n7552 ;
  assign n11097 = n11095 | n11096 ;
  assign n11098 = ( ~x56 & n11091 ) | ( ~x56 & n11097 ) | ( n11091 & n11097 ) ;
  assign n11099 = x56 & ~n11097 ;
  assign n11100 = ( ~n11092 & n11098 ) | ( ~n11092 & n11099 ) | ( n11098 & n11099 ) ;
  assign n11101 = n565 & n8067 ;
  assign n11102 = x59 & n11101 ;
  assign n11103 = x76 & n8074 ;
  assign n11104 = x75 & n8071 ;
  assign n11105 = n11103 | n11104 ;
  assign n11106 = x74 & n8298 ;
  assign n11107 = n11105 | n11106 ;
  assign n11108 = ( ~x59 & n11101 ) | ( ~x59 & n11107 ) | ( n11101 & n11107 ) ;
  assign n11109 = x59 & ~n11107 ;
  assign n11110 = ( ~n11102 & n11108 ) | ( ~n11102 & n11109 ) | ( n11108 & n11109 ) ;
  assign n11111 = ( x62 & x63 ) | ( x62 & x70 ) | ( x63 & x70 ) ;
  assign n11112 = ( x62 & x69 ) | ( x62 & ~n9394 ) | ( x69 & ~n9394 ) ;
  assign n11113 = ( x69 & n11111 ) | ( x69 & ~n11112 ) | ( n11111 & ~n11112 ) ;
  assign n11114 = ( x2 & ~x5 ) | ( x2 & n11113 ) | ( ~x5 & n11113 ) ;
  assign n11115 = ( x2 & x5 ) | ( x2 & ~n11113 ) | ( x5 & ~n11113 ) ;
  assign n11116 = ( ~x2 & n11114 ) | ( ~x2 & n11115 ) | ( n11114 & n11115 ) ;
  assign n11117 = n388 & n8859 ;
  assign n11118 = x62 & n11117 ;
  assign n11119 = x73 & n8866 ;
  assign n11120 = x72 & n8863 ;
  assign n11121 = n11119 | n11120 ;
  assign n11122 = x71 & n9125 ;
  assign n11123 = n11121 | n11122 ;
  assign n11124 = ( ~x62 & n11117 ) | ( ~x62 & n11123 ) | ( n11117 & n11123 ) ;
  assign n11125 = x62 & ~n11123 ;
  assign n11126 = ( ~n11118 & n11124 ) | ( ~n11118 & n11125 ) | ( n11124 & n11125 ) ;
  assign n11127 = ( n10868 & ~n11116 ) | ( n10868 & n11126 ) | ( ~n11116 & n11126 ) ;
  assign n11128 = ( n10868 & n11116 ) | ( n10868 & n11126 ) | ( n11116 & n11126 ) ;
  assign n11129 = ( n11116 & n11127 ) | ( n11116 & ~n11128 ) | ( n11127 & ~n11128 ) ;
  assign n11130 = ( n10871 & n11110 ) | ( n10871 & n11129 ) | ( n11110 & n11129 ) ;
  assign n11131 = ( ~n10871 & n11110 ) | ( ~n10871 & n11129 ) | ( n11110 & n11129 ) ;
  assign n11132 = ( n10871 & ~n11130 ) | ( n10871 & n11131 ) | ( ~n11130 & n11131 ) ;
  assign n11133 = ( n10885 & n11100 ) | ( n10885 & n11132 ) | ( n11100 & n11132 ) ;
  assign n11134 = ( n10885 & ~n11100 ) | ( n10885 & n11132 ) | ( ~n11100 & n11132 ) ;
  assign n11135 = ( n11100 & ~n11133 ) | ( n11100 & n11134 ) | ( ~n11133 & n11134 ) ;
  assign n11136 = ( n10887 & n11090 ) | ( n10887 & n11135 ) | ( n11090 & n11135 ) ;
  assign n11137 = ( n10887 & ~n11090 ) | ( n10887 & n11135 ) | ( ~n11090 & n11135 ) ;
  assign n11138 = ( n11090 & ~n11136 ) | ( n11090 & n11137 ) | ( ~n11136 & n11137 ) ;
  assign n11139 = ( ~n10890 & n11080 ) | ( ~n10890 & n11138 ) | ( n11080 & n11138 ) ;
  assign n11140 = ( n10890 & n11080 ) | ( n10890 & n11138 ) | ( n11080 & n11138 ) ;
  assign n11141 = ( n10890 & n11139 ) | ( n10890 & ~n11140 ) | ( n11139 & ~n11140 ) ;
  assign n11142 = ( n10893 & n11070 ) | ( n10893 & n11141 ) | ( n11070 & n11141 ) ;
  assign n11143 = ( ~n10893 & n11070 ) | ( ~n10893 & n11141 ) | ( n11070 & n11141 ) ;
  assign n11144 = ( n10893 & ~n11142 ) | ( n10893 & n11143 ) | ( ~n11142 & n11143 ) ;
  assign n11145 = n1959 & n4625 ;
  assign n11146 = x44 & n11145 ;
  assign n11147 = x91 & n4791 ;
  assign n11148 = x90 & n4621 ;
  assign n11149 = n11147 | n11148 ;
  assign n11150 = x89 & n4795 ;
  assign n11151 = n11149 | n11150 ;
  assign n11152 = ( ~x44 & n11145 ) | ( ~x44 & n11151 ) | ( n11145 & n11151 ) ;
  assign n11153 = x44 & ~n11151 ;
  assign n11154 = ( ~n11146 & n11152 ) | ( ~n11146 & n11153 ) | ( n11152 & n11153 ) ;
  assign n11155 = ( n10896 & ~n11144 ) | ( n10896 & n11154 ) | ( ~n11144 & n11154 ) ;
  assign n11156 = ( n10896 & n11144 ) | ( n10896 & n11154 ) | ( n11144 & n11154 ) ;
  assign n11157 = ( n11144 & n11155 ) | ( n11144 & ~n11156 ) | ( n11155 & ~n11156 ) ;
  assign n11158 = ( n10900 & n11060 ) | ( n10900 & n11157 ) | ( n11060 & n11157 ) ;
  assign n11159 = ( ~n10900 & n11060 ) | ( ~n10900 & n11157 ) | ( n11060 & n11157 ) ;
  assign n11160 = ( n10900 & ~n11158 ) | ( n10900 & n11159 ) | ( ~n11158 & n11159 ) ;
  assign n11161 = ( n10902 & n11050 ) | ( n10902 & n11160 ) | ( n11050 & n11160 ) ;
  assign n11162 = ( n10902 & ~n11050 ) | ( n10902 & n11160 ) | ( ~n11050 & n11160 ) ;
  assign n11163 = ( n11050 & ~n11161 ) | ( n11050 & n11162 ) | ( ~n11161 & n11162 ) ;
  assign n11164 = ( n10906 & n11040 ) | ( n10906 & n11163 ) | ( n11040 & n11163 ) ;
  assign n11165 = ( ~n10906 & n11040 ) | ( ~n10906 & n11163 ) | ( n11040 & n11163 ) ;
  assign n11166 = ( n10906 & ~n11164 ) | ( n10906 & n11165 ) | ( ~n11164 & n11165 ) ;
  assign n11167 = ( ~n10909 & n11030 ) | ( ~n10909 & n11166 ) | ( n11030 & n11166 ) ;
  assign n11168 = ( n10909 & n11030 ) | ( n10909 & n11166 ) | ( n11030 & n11166 ) ;
  assign n11169 = ( n10909 & n11167 ) | ( n10909 & ~n11168 ) | ( n11167 & ~n11168 ) ;
  assign n11170 = ( n10911 & n11020 ) | ( n10911 & n11169 ) | ( n11020 & n11169 ) ;
  assign n11171 = ( ~n10911 & n11020 ) | ( ~n10911 & n11169 ) | ( n11020 & n11169 ) ;
  assign n11172 = ( n10911 & ~n11170 ) | ( n10911 & n11171 ) | ( ~n11170 & n11171 ) ;
  assign n11173 = ( n10915 & n11010 ) | ( n10915 & n11172 ) | ( n11010 & n11172 ) ;
  assign n11174 = ( n10915 & ~n11010 ) | ( n10915 & n11172 ) | ( ~n11010 & n11172 ) ;
  assign n11175 = ( n11010 & ~n11173 ) | ( n11010 & n11174 ) | ( ~n11173 & n11174 ) ;
  assign n11176 = ( n10917 & n11000 ) | ( n10917 & n11175 ) | ( n11000 & n11175 ) ;
  assign n11177 = ( ~n10917 & n11000 ) | ( ~n10917 & n11175 ) | ( n11000 & n11175 ) ;
  assign n11178 = ( n10917 & ~n11176 ) | ( n10917 & n11177 ) | ( ~n11176 & n11177 ) ;
  assign n11179 = ( n10920 & n10990 ) | ( n10920 & n11178 ) | ( n10990 & n11178 ) ;
  assign n11180 = ( ~n10920 & n10990 ) | ( ~n10920 & n11178 ) | ( n10990 & n11178 ) ;
  assign n11181 = ( n10920 & ~n11179 ) | ( n10920 & n11180 ) | ( ~n11179 & n11180 ) ;
  assign n11182 = ( n10923 & n10980 ) | ( n10923 & n11181 ) | ( n10980 & n11181 ) ;
  assign n11183 = ( ~n10923 & n10980 ) | ( ~n10923 & n11181 ) | ( n10980 & n11181 ) ;
  assign n11184 = ( n10923 & ~n11182 ) | ( n10923 & n11183 ) | ( ~n11182 & n11183 ) ;
  assign n11185 = ( n10926 & n10970 ) | ( n10926 & n11184 ) | ( n10970 & n11184 ) ;
  assign n11186 = ( ~n10926 & n10970 ) | ( ~n10926 & n11184 ) | ( n10970 & n11184 ) ;
  assign n11187 = ( n10926 & ~n11185 ) | ( n10926 & n11186 ) | ( ~n11185 & n11186 ) ;
  assign n11188 = ( n10929 & n10960 ) | ( n10929 & n11187 ) | ( n10960 & n11187 ) ;
  assign n11189 = ( ~n10929 & n10960 ) | ( ~n10929 & n11187 ) | ( n10960 & n11187 ) ;
  assign n11190 = ( n10929 & ~n11188 ) | ( n10929 & n11189 ) | ( ~n11188 & n11189 ) ;
  assign n11191 = ( n10932 & n10950 ) | ( n10932 & n11190 ) | ( n10950 & n11190 ) ;
  assign n11192 = ( ~n10932 & n10950 ) | ( ~n10932 & n11190 ) | ( n10950 & n11190 ) ;
  assign n11193 = ( n10932 & ~n11191 ) | ( n10932 & n11192 ) | ( ~n11191 & n11192 ) ;
  assign n11194 = ( n10936 & ~n10939 ) | ( n10936 & n11193 ) | ( ~n10939 & n11193 ) ;
  assign n11195 = ( n10936 & n10939 ) | ( n10936 & n11193 ) | ( n10939 & n11193 ) ;
  assign n11196 = ( n10939 & n11194 ) | ( n10939 & ~n11195 ) | ( n11194 & ~n11195 ) ;
  assign n11197 = x127 & n306 ;
  assign n11198 = n301 | n11197 ;
  assign n11199 = ( n9867 & n11197 ) | ( n9867 & n11198 ) | ( n11197 & n11198 ) ;
  assign n11200 = x126 & n359 ;
  assign n11201 = ( ~x8 & n11199 ) | ( ~x8 & n11200 ) | ( n11199 & n11200 ) ;
  assign n11202 = ( x8 & ~n11199 ) | ( x8 & n11200 ) | ( ~n11199 & n11200 ) ;
  assign n11203 = ~n11200 & n11202 ;
  assign n11204 = n11201 | n11203 ;
  assign n11205 = n449 & n9009 ;
  assign n11206 = x11 & n11205 ;
  assign n11207 = x125 & n456 ;
  assign n11208 = x124 & n453 ;
  assign n11209 = n11207 | n11208 ;
  assign n11210 = x123 & n536 ;
  assign n11211 = n11209 | n11210 ;
  assign n11212 = ( ~x11 & n11205 ) | ( ~x11 & n11211 ) | ( n11205 & n11211 ) ;
  assign n11213 = x11 & ~n11211 ;
  assign n11214 = ( ~n11206 & n11212 ) | ( ~n11206 & n11213 ) | ( n11212 & n11213 ) ;
  assign n11215 = n649 & n8207 ;
  assign n11216 = x14 & n11215 ;
  assign n11217 = x122 & n656 ;
  assign n11218 = x121 & n653 ;
  assign n11219 = n11217 | n11218 ;
  assign n11220 = x120 & n744 ;
  assign n11221 = n11219 | n11220 ;
  assign n11222 = ( ~x14 & n11215 ) | ( ~x14 & n11221 ) | ( n11215 & n11221 ) ;
  assign n11223 = x14 & ~n11221 ;
  assign n11224 = ( ~n11216 & n11222 ) | ( ~n11216 & n11223 ) | ( n11222 & n11223 ) ;
  assign n11225 = n874 & n7181 ;
  assign n11226 = x17 & n11225 ;
  assign n11227 = x119 & n881 ;
  assign n11228 = x118 & n878 ;
  assign n11229 = n11227 | n11228 ;
  assign n11230 = x117 & n959 ;
  assign n11231 = n11229 | n11230 ;
  assign n11232 = ( ~x17 & n11225 ) | ( ~x17 & n11231 ) | ( n11225 & n11231 ) ;
  assign n11233 = x17 & ~n11231 ;
  assign n11234 = ( ~n11226 & n11232 ) | ( ~n11226 & n11233 ) | ( n11232 & n11233 ) ;
  assign n11235 = n1146 & n6462 ;
  assign n11236 = x20 & n11235 ;
  assign n11237 = x116 & n1153 ;
  assign n11238 = x115 & n1150 ;
  assign n11239 = n11237 | n11238 ;
  assign n11240 = x114 & n1217 ;
  assign n11241 = n11239 | n11240 ;
  assign n11242 = ( ~x20 & n11235 ) | ( ~x20 & n11241 ) | ( n11235 & n11241 ) ;
  assign n11243 = x20 & ~n11241 ;
  assign n11244 = ( ~n11236 & n11242 ) | ( ~n11236 & n11243 ) | ( n11242 & n11243 ) ;
  assign n11245 = n1427 & n5774 ;
  assign n11246 = x23 & n11245 ;
  assign n11247 = x113 & n1434 ;
  assign n11248 = x112 & n1431 ;
  assign n11249 = n11247 | n11248 ;
  assign n11250 = x111 & n1531 ;
  assign n11251 = n11249 | n11250 ;
  assign n11252 = ( ~x23 & n11245 ) | ( ~x23 & n11251 ) | ( n11245 & n11251 ) ;
  assign n11253 = x23 & ~n11251 ;
  assign n11254 = ( ~n11246 & n11252 ) | ( ~n11246 & n11253 ) | ( n11252 & n11253 ) ;
  assign n11255 = n1755 & n5331 ;
  assign n11256 = x26 & n11255 ;
  assign n11257 = x110 & n1762 ;
  assign n11258 = x109 & n1759 ;
  assign n11259 = n11257 | n11258 ;
  assign n11260 = x108 & n1895 ;
  assign n11261 = n11259 | n11260 ;
  assign n11262 = ( ~x26 & n11255 ) | ( ~x26 & n11261 ) | ( n11255 & n11261 ) ;
  assign n11263 = x26 & ~n11261 ;
  assign n11264 = ( ~n11256 & n11262 ) | ( ~n11256 & n11263 ) | ( n11262 & n11263 ) ;
  assign n11265 = n2137 & n4523 ;
  assign n11266 = x29 & n11265 ;
  assign n11267 = x107 & n2144 ;
  assign n11268 = x106 & n2141 ;
  assign n11269 = n11267 | n11268 ;
  assign n11270 = x105 & n2267 ;
  assign n11271 = n11269 | n11270 ;
  assign n11272 = ( ~x29 & n11265 ) | ( ~x29 & n11271 ) | ( n11265 & n11271 ) ;
  assign n11273 = x29 & ~n11271 ;
  assign n11274 = ( ~n11266 & n11272 ) | ( ~n11266 & n11273 ) | ( n11272 & n11273 ) ;
  assign n11275 = n2545 & n3957 ;
  assign n11276 = x32 & n11275 ;
  assign n11277 = x104 & n2552 ;
  assign n11278 = x103 & n2549 ;
  assign n11279 = n11277 | n11278 ;
  assign n11280 = x102 & n2696 ;
  assign n11281 = n11279 | n11280 ;
  assign n11282 = ( ~x32 & n11275 ) | ( ~x32 & n11281 ) | ( n11275 & n11281 ) ;
  assign n11283 = x32 & ~n11281 ;
  assign n11284 = ( ~n11276 & n11282 ) | ( ~n11276 & n11283 ) | ( n11282 & n11283 ) ;
  assign n11285 = n2982 & n3591 ;
  assign n11286 = x35 & n11285 ;
  assign n11287 = x101 & n2989 ;
  assign n11288 = x100 & n2986 ;
  assign n11289 = n11287 | n11288 ;
  assign n11290 = x99 & n3159 ;
  assign n11291 = n11289 | n11290 ;
  assign n11292 = ( ~x35 & n11285 ) | ( ~x35 & n11291 ) | ( n11285 & n11291 ) ;
  assign n11293 = x35 & ~n11291 ;
  assign n11294 = ( ~n11286 & n11292 ) | ( ~n11286 & n11293 ) | ( n11292 & n11293 ) ;
  assign n11295 = n2939 & n3492 ;
  assign n11296 = x38 & n11295 ;
  assign n11297 = x98 & n3499 ;
  assign n11298 = x97 & n3496 ;
  assign n11299 = n11297 | n11298 ;
  assign n11300 = x96 & n3662 ;
  assign n11301 = n11299 | n11300 ;
  assign n11302 = ( ~x38 & n11295 ) | ( ~x38 & n11301 ) | ( n11295 & n11301 ) ;
  assign n11303 = x38 & ~n11301 ;
  assign n11304 = ( ~n11296 & n11302 ) | ( ~n11296 & n11303 ) | ( n11302 & n11303 ) ;
  assign n11305 = n2492 & n4020 ;
  assign n11306 = x41 & n11305 ;
  assign n11307 = x95 & n4027 ;
  assign n11308 = x94 & n4024 ;
  assign n11309 = n11307 | n11308 ;
  assign n11310 = x93 & n4223 ;
  assign n11311 = n11309 | n11310 ;
  assign n11312 = ( ~x41 & n11305 ) | ( ~x41 & n11311 ) | ( n11305 & n11311 ) ;
  assign n11313 = x41 & ~n11311 ;
  assign n11314 = ( ~n11306 & n11312 ) | ( ~n11306 & n11313 ) | ( n11312 & n11313 ) ;
  assign n11315 = n2083 & n4625 ;
  assign n11316 = x44 & n11315 ;
  assign n11317 = x92 & n4791 ;
  assign n11318 = x91 & n4621 ;
  assign n11319 = n11317 | n11318 ;
  assign n11320 = x90 & n4795 ;
  assign n11321 = n11319 | n11320 ;
  assign n11322 = ( ~x44 & n11315 ) | ( ~x44 & n11321 ) | ( n11315 & n11321 ) ;
  assign n11323 = x44 & ~n11321 ;
  assign n11324 = ( ~n11316 & n11322 ) | ( ~n11316 & n11323 ) | ( n11322 & n11323 ) ;
  assign n11325 = n1822 & n5223 ;
  assign n11326 = x47 & n11325 ;
  assign n11327 = x89 & n5230 ;
  assign n11328 = x88 & n5227 ;
  assign n11329 = n11327 | n11328 ;
  assign n11330 = x87 & n5434 ;
  assign n11331 = n11329 | n11330 ;
  assign n11332 = ( ~x47 & n11325 ) | ( ~x47 & n11331 ) | ( n11325 & n11331 ) ;
  assign n11333 = x47 & ~n11331 ;
  assign n11334 = ( ~n11326 & n11332 ) | ( ~n11326 & n11333 ) | ( n11332 & n11333 ) ;
  assign n11335 = n1384 & n5858 ;
  assign n11336 = x50 & n11335 ;
  assign n11337 = x86 & n5865 ;
  assign n11338 = x85 & n5862 ;
  assign n11339 = n11337 | n11338 ;
  assign n11340 = x84 & n6092 ;
  assign n11341 = n11339 | n11340 ;
  assign n11342 = ( ~x50 & n11335 ) | ( ~x50 & n11341 ) | ( n11335 & n11341 ) ;
  assign n11343 = x50 & ~n11341 ;
  assign n11344 = ( ~n11336 & n11342 ) | ( ~n11336 & n11343 ) | ( n11342 & n11343 ) ;
  assign n11345 = n1093 & n6546 ;
  assign n11346 = x53 & n11345 ;
  assign n11347 = x83 & n6553 ;
  assign n11348 = x82 & n6550 ;
  assign n11349 = n11347 | n11348 ;
  assign n11350 = x81 & n6787 ;
  assign n11351 = n11349 | n11350 ;
  assign n11352 = ( ~x53 & n11345 ) | ( ~x53 & n11351 ) | ( n11345 & n11351 ) ;
  assign n11353 = x53 & ~n11351 ;
  assign n11354 = ( ~n11346 & n11352 ) | ( ~n11346 & n11353 ) | ( n11352 & n11353 ) ;
  assign n11355 = n840 & n7277 ;
  assign n11356 = x56 & n11355 ;
  assign n11357 = x80 & n7545 ;
  assign n11358 = x79 & n7273 ;
  assign n11359 = n11357 | n11358 ;
  assign n11360 = x78 & n7552 ;
  assign n11361 = n11359 | n11360 ;
  assign n11362 = ( ~x56 & n11355 ) | ( ~x56 & n11361 ) | ( n11355 & n11361 ) ;
  assign n11363 = x56 & ~n11361 ;
  assign n11364 = ( ~n11356 & n11362 ) | ( ~n11356 & n11363 ) | ( n11362 & n11363 ) ;
  assign n11365 = n626 & n8067 ;
  assign n11366 = x59 & n11365 ;
  assign n11367 = x77 & n8074 ;
  assign n11368 = x76 & n8071 ;
  assign n11369 = n11367 | n11368 ;
  assign n11370 = x75 & n8298 ;
  assign n11371 = n11369 | n11370 ;
  assign n11372 = ( ~x59 & n11365 ) | ( ~x59 & n11371 ) | ( n11365 & n11371 ) ;
  assign n11373 = x59 & ~n11371 ;
  assign n11374 = ( ~n11366 & n11372 ) | ( ~n11366 & n11373 ) | ( n11372 & n11373 ) ;
  assign n11375 = n436 & n8859 ;
  assign n11376 = x62 & n11375 ;
  assign n11377 = x74 & n8866 ;
  assign n11378 = x73 & n8863 ;
  assign n11379 = n11377 | n11378 ;
  assign n11380 = x72 & n9125 ;
  assign n11381 = n11379 | n11380 ;
  assign n11382 = ( ~x62 & n11375 ) | ( ~x62 & n11381 ) | ( n11375 & n11381 ) ;
  assign n11383 = x62 & ~n11381 ;
  assign n11384 = ( ~n11376 & n11382 ) | ( ~n11376 & n11383 ) | ( n11382 & n11383 ) ;
  assign n11385 = ( x62 & x63 ) | ( x62 & x71 ) | ( x63 & x71 ) ;
  assign n11386 = ( x62 & x70 ) | ( x62 & ~n9394 ) | ( x70 & ~n9394 ) ;
  assign n11387 = ( x70 & n11385 ) | ( x70 & ~n11386 ) | ( n11385 & ~n11386 ) ;
  assign n11388 = ( n11115 & ~n11384 ) | ( n11115 & n11387 ) | ( ~n11384 & n11387 ) ;
  assign n11389 = ( n11115 & n11384 ) | ( n11115 & n11387 ) | ( n11384 & n11387 ) ;
  assign n11390 = ( n11384 & n11388 ) | ( n11384 & ~n11389 ) | ( n11388 & ~n11389 ) ;
  assign n11391 = ( n11128 & n11374 ) | ( n11128 & n11390 ) | ( n11374 & n11390 ) ;
  assign n11392 = ( n11128 & ~n11374 ) | ( n11128 & n11390 ) | ( ~n11374 & n11390 ) ;
  assign n11393 = ( n11374 & ~n11391 ) | ( n11374 & n11392 ) | ( ~n11391 & n11392 ) ;
  assign n11394 = ( n11130 & n11364 ) | ( n11130 & n11393 ) | ( n11364 & n11393 ) ;
  assign n11395 = ( n11130 & ~n11364 ) | ( n11130 & n11393 ) | ( ~n11364 & n11393 ) ;
  assign n11396 = ( n11364 & ~n11394 ) | ( n11364 & n11395 ) | ( ~n11394 & n11395 ) ;
  assign n11397 = ( n11133 & n11354 ) | ( n11133 & n11396 ) | ( n11354 & n11396 ) ;
  assign n11398 = ( n11133 & ~n11354 ) | ( n11133 & n11396 ) | ( ~n11354 & n11396 ) ;
  assign n11399 = ( n11354 & ~n11397 ) | ( n11354 & n11398 ) | ( ~n11397 & n11398 ) ;
  assign n11400 = ( n11136 & n11344 ) | ( n11136 & n11399 ) | ( n11344 & n11399 ) ;
  assign n11401 = ( n11136 & ~n11344 ) | ( n11136 & n11399 ) | ( ~n11344 & n11399 ) ;
  assign n11402 = ( n11344 & ~n11400 ) | ( n11344 & n11401 ) | ( ~n11400 & n11401 ) ;
  assign n11403 = ( n11140 & ~n11334 ) | ( n11140 & n11402 ) | ( ~n11334 & n11402 ) ;
  assign n11404 = ( n11140 & n11334 ) | ( n11140 & n11402 ) | ( n11334 & n11402 ) ;
  assign n11405 = ( n11334 & n11403 ) | ( n11334 & ~n11404 ) | ( n11403 & ~n11404 ) ;
  assign n11406 = ( n11142 & n11324 ) | ( n11142 & n11405 ) | ( n11324 & n11405 ) ;
  assign n11407 = ( n11142 & ~n11324 ) | ( n11142 & n11405 ) | ( ~n11324 & n11405 ) ;
  assign n11408 = ( n11324 & ~n11406 ) | ( n11324 & n11407 ) | ( ~n11406 & n11407 ) ;
  assign n11409 = ( n11156 & n11314 ) | ( n11156 & n11408 ) | ( n11314 & n11408 ) ;
  assign n11410 = ( n11156 & ~n11314 ) | ( n11156 & n11408 ) | ( ~n11314 & n11408 ) ;
  assign n11411 = ( n11314 & ~n11409 ) | ( n11314 & n11410 ) | ( ~n11409 & n11410 ) ;
  assign n11412 = ( n11158 & n11304 ) | ( n11158 & n11411 ) | ( n11304 & n11411 ) ;
  assign n11413 = ( n11158 & ~n11304 ) | ( n11158 & n11411 ) | ( ~n11304 & n11411 ) ;
  assign n11414 = ( n11304 & ~n11412 ) | ( n11304 & n11413 ) | ( ~n11412 & n11413 ) ;
  assign n11415 = ( n11161 & n11294 ) | ( n11161 & n11414 ) | ( n11294 & n11414 ) ;
  assign n11416 = ( n11161 & ~n11294 ) | ( n11161 & n11414 ) | ( ~n11294 & n11414 ) ;
  assign n11417 = ( n11294 & ~n11415 ) | ( n11294 & n11416 ) | ( ~n11415 & n11416 ) ;
  assign n11418 = ( n11164 & n11284 ) | ( n11164 & n11417 ) | ( n11284 & n11417 ) ;
  assign n11419 = ( n11164 & ~n11284 ) | ( n11164 & n11417 ) | ( ~n11284 & n11417 ) ;
  assign n11420 = ( n11284 & ~n11418 ) | ( n11284 & n11419 ) | ( ~n11418 & n11419 ) ;
  assign n11421 = ( n11168 & n11274 ) | ( n11168 & n11420 ) | ( n11274 & n11420 ) ;
  assign n11422 = ( n11168 & ~n11274 ) | ( n11168 & n11420 ) | ( ~n11274 & n11420 ) ;
  assign n11423 = ( n11274 & ~n11421 ) | ( n11274 & n11422 ) | ( ~n11421 & n11422 ) ;
  assign n11424 = ( n11170 & n11264 ) | ( n11170 & n11423 ) | ( n11264 & n11423 ) ;
  assign n11425 = ( n11170 & ~n11264 ) | ( n11170 & n11423 ) | ( ~n11264 & n11423 ) ;
  assign n11426 = ( n11264 & ~n11424 ) | ( n11264 & n11425 ) | ( ~n11424 & n11425 ) ;
  assign n11427 = ( n11173 & n11254 ) | ( n11173 & n11426 ) | ( n11254 & n11426 ) ;
  assign n11428 = ( n11173 & ~n11254 ) | ( n11173 & n11426 ) | ( ~n11254 & n11426 ) ;
  assign n11429 = ( n11254 & ~n11427 ) | ( n11254 & n11428 ) | ( ~n11427 & n11428 ) ;
  assign n11430 = ( n11176 & n11244 ) | ( n11176 & n11429 ) | ( n11244 & n11429 ) ;
  assign n11431 = ( n11176 & ~n11244 ) | ( n11176 & n11429 ) | ( ~n11244 & n11429 ) ;
  assign n11432 = ( n11244 & ~n11430 ) | ( n11244 & n11431 ) | ( ~n11430 & n11431 ) ;
  assign n11433 = ( n11179 & n11234 ) | ( n11179 & n11432 ) | ( n11234 & n11432 ) ;
  assign n11434 = ( n11179 & ~n11234 ) | ( n11179 & n11432 ) | ( ~n11234 & n11432 ) ;
  assign n11435 = ( n11234 & ~n11433 ) | ( n11234 & n11434 ) | ( ~n11433 & n11434 ) ;
  assign n11436 = ( n11182 & n11224 ) | ( n11182 & n11435 ) | ( n11224 & n11435 ) ;
  assign n11437 = ( n11182 & ~n11224 ) | ( n11182 & n11435 ) | ( ~n11224 & n11435 ) ;
  assign n11438 = ( n11224 & ~n11436 ) | ( n11224 & n11437 ) | ( ~n11436 & n11437 ) ;
  assign n11439 = ( n11185 & n11214 ) | ( n11185 & n11438 ) | ( n11214 & n11438 ) ;
  assign n11440 = ( n11185 & ~n11214 ) | ( n11185 & n11438 ) | ( ~n11214 & n11438 ) ;
  assign n11441 = ( n11214 & ~n11439 ) | ( n11214 & n11440 ) | ( ~n11439 & n11440 ) ;
  assign n11442 = ( n11188 & n11204 ) | ( n11188 & n11441 ) | ( n11204 & n11441 ) ;
  assign n11443 = ( n11188 & ~n11204 ) | ( n11188 & n11441 ) | ( ~n11204 & n11441 ) ;
  assign n11444 = ( n11204 & ~n11442 ) | ( n11204 & n11443 ) | ( ~n11442 & n11443 ) ;
  assign n11445 = ( n11191 & ~n11195 ) | ( n11191 & n11444 ) | ( ~n11195 & n11444 ) ;
  assign n11446 = ( n11191 & n11195 ) | ( n11191 & n11444 ) | ( n11195 & n11444 ) ;
  assign n11447 = ( n11195 & n11445 ) | ( n11195 & ~n11446 ) | ( n11445 & ~n11446 ) ;
  assign n11448 = n449 & n9038 ;
  assign n11449 = x11 & n11448 ;
  assign n11450 = x126 & n456 ;
  assign n11451 = x125 & n453 ;
  assign n11452 = n11450 | n11451 ;
  assign n11453 = x124 & n536 ;
  assign n11454 = n11452 | n11453 ;
  assign n11455 = ( ~x11 & n11448 ) | ( ~x11 & n11454 ) | ( n11448 & n11454 ) ;
  assign n11456 = x11 & ~n11454 ;
  assign n11457 = ( ~n11449 & n11455 ) | ( ~n11449 & n11456 ) | ( n11455 & n11456 ) ;
  assign n11458 = n649 & n8461 ;
  assign n11459 = x14 & n11458 ;
  assign n11460 = x123 & n656 ;
  assign n11461 = x122 & n653 ;
  assign n11462 = n11460 | n11461 ;
  assign n11463 = x121 & n744 ;
  assign n11464 = n11462 | n11463 ;
  assign n11465 = ( ~x14 & n11458 ) | ( ~x14 & n11464 ) | ( n11458 & n11464 ) ;
  assign n11466 = x14 & ~n11464 ;
  assign n11467 = ( ~n11459 & n11465 ) | ( ~n11459 & n11466 ) | ( n11465 & n11466 ) ;
  assign n11468 = n874 & n7444 ;
  assign n11469 = x17 & n11468 ;
  assign n11470 = x120 & n881 ;
  assign n11471 = x119 & n878 ;
  assign n11472 = n11470 | n11471 ;
  assign n11473 = x118 & n959 ;
  assign n11474 = n11472 | n11473 ;
  assign n11475 = ( ~x17 & n11468 ) | ( ~x17 & n11474 ) | ( n11468 & n11474 ) ;
  assign n11476 = x17 & ~n11474 ;
  assign n11477 = ( ~n11469 & n11475 ) | ( ~n11469 & n11476 ) | ( n11475 & n11476 ) ;
  assign n11478 = n1146 & n6924 ;
  assign n11479 = x20 & n11478 ;
  assign n11480 = x117 & n1153 ;
  assign n11481 = x116 & n1150 ;
  assign n11482 = n11480 | n11481 ;
  assign n11483 = x115 & n1217 ;
  assign n11484 = n11482 | n11483 ;
  assign n11485 = ( ~x20 & n11478 ) | ( ~x20 & n11484 ) | ( n11478 & n11484 ) ;
  assign n11486 = x20 & ~n11484 ;
  assign n11487 = ( ~n11479 & n11485 ) | ( ~n11479 & n11486 ) | ( n11485 & n11486 ) ;
  assign n11488 = n1427 & n6002 ;
  assign n11489 = x23 & n11488 ;
  assign n11490 = x114 & n1434 ;
  assign n11491 = x113 & n1431 ;
  assign n11492 = n11490 | n11491 ;
  assign n11493 = x112 & n1531 ;
  assign n11494 = n11492 | n11493 ;
  assign n11495 = ( ~x23 & n11488 ) | ( ~x23 & n11494 ) | ( n11488 & n11494 ) ;
  assign n11496 = x23 & ~n11494 ;
  assign n11497 = ( ~n11489 & n11495 ) | ( ~n11489 & n11496 ) | ( n11495 & n11496 ) ;
  assign n11498 = n1755 & n5347 ;
  assign n11499 = x26 & n11498 ;
  assign n11500 = x111 & n1762 ;
  assign n11501 = x110 & n1759 ;
  assign n11502 = n11500 | n11501 ;
  assign n11503 = x109 & n1895 ;
  assign n11504 = n11502 | n11503 ;
  assign n11505 = ( ~x26 & n11498 ) | ( ~x26 & n11504 ) | ( n11498 & n11504 ) ;
  assign n11506 = x26 & ~n11504 ;
  assign n11507 = ( ~n11499 & n11505 ) | ( ~n11499 & n11506 ) | ( n11505 & n11506 ) ;
  assign n11508 = n2137 & n4914 ;
  assign n11509 = x29 & n11508 ;
  assign n11510 = x108 & n2144 ;
  assign n11511 = x107 & n2141 ;
  assign n11512 = n11510 | n11511 ;
  assign n11513 = x106 & n2267 ;
  assign n11514 = n11512 | n11513 ;
  assign n11515 = ( ~x29 & n11508 ) | ( ~x29 & n11514 ) | ( n11508 & n11514 ) ;
  assign n11516 = x29 & ~n11514 ;
  assign n11517 = ( ~n11509 & n11515 ) | ( ~n11509 & n11516 ) | ( n11515 & n11516 ) ;
  assign n11518 = n2545 & n4145 ;
  assign n11519 = x32 & n11518 ;
  assign n11520 = x105 & n2552 ;
  assign n11521 = x104 & n2549 ;
  assign n11522 = n11520 | n11521 ;
  assign n11523 = x103 & n2696 ;
  assign n11524 = n11522 | n11523 ;
  assign n11525 = ( ~x32 & n11518 ) | ( ~x32 & n11524 ) | ( n11518 & n11524 ) ;
  assign n11526 = x32 & ~n11524 ;
  assign n11527 = ( ~n11519 & n11525 ) | ( ~n11519 & n11526 ) | ( n11525 & n11526 ) ;
  assign n11528 = n2982 & n3764 ;
  assign n11529 = x35 & n11528 ;
  assign n11530 = x102 & n2989 ;
  assign n11531 = x101 & n2986 ;
  assign n11532 = n11530 | n11531 ;
  assign n11533 = x100 & n3159 ;
  assign n11534 = n11532 | n11533 ;
  assign n11535 = ( ~x35 & n11528 ) | ( ~x35 & n11534 ) | ( n11528 & n11534 ) ;
  assign n11536 = x35 & ~n11534 ;
  assign n11537 = ( ~n11529 & n11535 ) | ( ~n11529 & n11536 ) | ( n11535 & n11536 ) ;
  assign n11538 = n3248 & n3492 ;
  assign n11539 = x38 & n11538 ;
  assign n11540 = x99 & n3499 ;
  assign n11541 = x98 & n3496 ;
  assign n11542 = n11540 | n11541 ;
  assign n11543 = x97 & n3662 ;
  assign n11544 = n11542 | n11543 ;
  assign n11545 = ( ~x38 & n11538 ) | ( ~x38 & n11544 ) | ( n11538 & n11544 ) ;
  assign n11546 = x38 & ~n11544 ;
  assign n11547 = ( ~n11539 & n11545 ) | ( ~n11539 & n11546 ) | ( n11545 & n11546 ) ;
  assign n11548 = n2772 & n4020 ;
  assign n11549 = x41 & n11548 ;
  assign n11550 = x96 & n4027 ;
  assign n11551 = x95 & n4024 ;
  assign n11552 = n11550 | n11551 ;
  assign n11553 = x94 & n4223 ;
  assign n11554 = n11552 | n11553 ;
  assign n11555 = ( ~x41 & n11548 ) | ( ~x41 & n11554 ) | ( n11548 & n11554 ) ;
  assign n11556 = x41 & ~n11554 ;
  assign n11557 = ( ~n11549 & n11555 ) | ( ~n11549 & n11556 ) | ( n11555 & n11556 ) ;
  assign n11558 = x93 & n4791 ;
  assign n11559 = x44 & n11558 ;
  assign n11560 = x92 & n4621 ;
  assign n11561 = x91 | n11560 ;
  assign n11562 = ( n4795 & n11560 ) | ( n4795 & n11561 ) | ( n11560 & n11561 ) ;
  assign n11563 = n2220 & n4625 ;
  assign n11564 = n11562 | n11563 ;
  assign n11565 = ( ~x44 & n11558 ) | ( ~x44 & n11564 ) | ( n11558 & n11564 ) ;
  assign n11566 = x44 & ~n11564 ;
  assign n11567 = ( ~n11559 & n11565 ) | ( ~n11559 & n11566 ) | ( n11565 & n11566 ) ;
  assign n11568 = n1838 & n5223 ;
  assign n11569 = x47 & n11568 ;
  assign n11570 = x90 & n5230 ;
  assign n11571 = x89 & n5227 ;
  assign n11572 = n11570 | n11571 ;
  assign n11573 = x88 & n5434 ;
  assign n11574 = n11572 | n11573 ;
  assign n11575 = ( ~x47 & n11568 ) | ( ~x47 & n11574 ) | ( n11568 & n11574 ) ;
  assign n11576 = x47 & ~n11574 ;
  assign n11577 = ( ~n11569 & n11575 ) | ( ~n11569 & n11576 ) | ( n11575 & n11576 ) ;
  assign n11578 = n1494 & n5858 ;
  assign n11579 = x50 & n11578 ;
  assign n11580 = x87 & n5865 ;
  assign n11581 = x86 & n5862 ;
  assign n11582 = n11580 | n11581 ;
  assign n11583 = x85 & n6092 ;
  assign n11584 = n11582 | n11583 ;
  assign n11585 = ( ~x50 & n11578 ) | ( ~x50 & n11584 ) | ( n11578 & n11584 ) ;
  assign n11586 = x50 & ~n11584 ;
  assign n11587 = ( ~n11579 & n11585 ) | ( ~n11579 & n11586 ) | ( n11585 & n11586 ) ;
  assign n11588 = n1190 & n6546 ;
  assign n11589 = x53 & n11588 ;
  assign n11590 = x84 & n6553 ;
  assign n11591 = x83 & n6550 ;
  assign n11592 = n11590 | n11591 ;
  assign n11593 = x82 & n6787 ;
  assign n11594 = n11592 | n11593 ;
  assign n11595 = ( ~x53 & n11588 ) | ( ~x53 & n11594 ) | ( n11588 & n11594 ) ;
  assign n11596 = x53 & ~n11594 ;
  assign n11597 = ( ~n11589 & n11595 ) | ( ~n11589 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11598 = x78 & n8074 ;
  assign n11599 = x59 & n11598 ;
  assign n11600 = x77 & n8071 ;
  assign n11601 = x76 | n11600 ;
  assign n11602 = ( n8298 & n11600 ) | ( n8298 & n11601 ) | ( n11600 & n11601 ) ;
  assign n11603 = n697 & n8067 ;
  assign n11604 = n11602 | n11603 ;
  assign n11605 = ( ~x59 & n11598 ) | ( ~x59 & n11604 ) | ( n11598 & n11604 ) ;
  assign n11606 = x59 & ~n11604 ;
  assign n11607 = ( ~n11599 & n11605 ) | ( ~n11599 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11608 = n508 & n8859 ;
  assign n11609 = x62 & n11608 ;
  assign n11610 = x75 & n8866 ;
  assign n11611 = x74 & n8863 ;
  assign n11612 = n11610 | n11611 ;
  assign n11613 = x73 & n9125 ;
  assign n11614 = n11612 | n11613 ;
  assign n11615 = ( ~x62 & n11608 ) | ( ~x62 & n11614 ) | ( n11608 & n11614 ) ;
  assign n11616 = x62 & ~n11614 ;
  assign n11617 = ( ~n11609 & n11615 ) | ( ~n11609 & n11616 ) | ( n11615 & n11616 ) ;
  assign n11618 = ( x62 & x63 ) | ( x62 & x72 ) | ( x63 & x72 ) ;
  assign n11619 = ( x62 & x71 ) | ( x62 & ~n9394 ) | ( x71 & ~n9394 ) ;
  assign n11620 = ( x71 & n11618 ) | ( x71 & ~n11619 ) | ( n11618 & ~n11619 ) ;
  assign n11621 = ( n11387 & n11388 ) | ( n11387 & n11620 ) | ( n11388 & n11620 ) ;
  assign n11622 = ( n11115 & ~n11389 ) | ( n11115 & n11620 ) | ( ~n11389 & n11620 ) ;
  assign n11623 = ( n11387 & ~n11621 ) | ( n11387 & n11622 ) | ( ~n11621 & n11622 ) ;
  assign n11624 = ( n11607 & n11617 ) | ( n11607 & n11623 ) | ( n11617 & n11623 ) ;
  assign n11625 = ( ~n11607 & n11617 ) | ( ~n11607 & n11623 ) | ( n11617 & n11623 ) ;
  assign n11626 = ( n11607 & ~n11624 ) | ( n11607 & n11625 ) | ( ~n11624 & n11625 ) ;
  assign n11627 = n990 & n7277 ;
  assign n11628 = x56 & n11627 ;
  assign n11629 = x81 & n7545 ;
  assign n11630 = x80 & n7273 ;
  assign n11631 = n11629 | n11630 ;
  assign n11632 = x79 & n7552 ;
  assign n11633 = n11631 | n11632 ;
  assign n11634 = ( ~x56 & n11627 ) | ( ~x56 & n11633 ) | ( n11627 & n11633 ) ;
  assign n11635 = x56 & ~n11633 ;
  assign n11636 = ( ~n11628 & n11634 ) | ( ~n11628 & n11635 ) | ( n11634 & n11635 ) ;
  assign n11637 = ( n11391 & n11626 ) | ( n11391 & n11636 ) | ( n11626 & n11636 ) ;
  assign n11638 = ( n11391 & ~n11626 ) | ( n11391 & n11636 ) | ( ~n11626 & n11636 ) ;
  assign n11639 = ( n11626 & ~n11637 ) | ( n11626 & n11638 ) | ( ~n11637 & n11638 ) ;
  assign n11640 = ( n11394 & ~n11597 ) | ( n11394 & n11639 ) | ( ~n11597 & n11639 ) ;
  assign n11641 = ( n11394 & n11597 ) | ( n11394 & n11639 ) | ( n11597 & n11639 ) ;
  assign n11642 = ( n11597 & n11640 ) | ( n11597 & ~n11641 ) | ( n11640 & ~n11641 ) ;
  assign n11643 = ( n11397 & n11587 ) | ( n11397 & n11642 ) | ( n11587 & n11642 ) ;
  assign n11644 = ( n11397 & ~n11587 ) | ( n11397 & n11642 ) | ( ~n11587 & n11642 ) ;
  assign n11645 = ( n11587 & ~n11643 ) | ( n11587 & n11644 ) | ( ~n11643 & n11644 ) ;
  assign n11646 = ( n11400 & n11577 ) | ( n11400 & n11645 ) | ( n11577 & n11645 ) ;
  assign n11647 = ( n11400 & ~n11577 ) | ( n11400 & n11645 ) | ( ~n11577 & n11645 ) ;
  assign n11648 = ( n11577 & ~n11646 ) | ( n11577 & n11647 ) | ( ~n11646 & n11647 ) ;
  assign n11649 = ( n11404 & n11567 ) | ( n11404 & n11648 ) | ( n11567 & n11648 ) ;
  assign n11650 = ( n11404 & ~n11567 ) | ( n11404 & n11648 ) | ( ~n11567 & n11648 ) ;
  assign n11651 = ( n11567 & ~n11649 ) | ( n11567 & n11650 ) | ( ~n11649 & n11650 ) ;
  assign n11652 = ( n11406 & n11557 ) | ( n11406 & n11651 ) | ( n11557 & n11651 ) ;
  assign n11653 = ( n11406 & ~n11557 ) | ( n11406 & n11651 ) | ( ~n11557 & n11651 ) ;
  assign n11654 = ( n11557 & ~n11652 ) | ( n11557 & n11653 ) | ( ~n11652 & n11653 ) ;
  assign n11655 = ( n11409 & n11547 ) | ( n11409 & n11654 ) | ( n11547 & n11654 ) ;
  assign n11656 = ( n11409 & ~n11547 ) | ( n11409 & n11654 ) | ( ~n11547 & n11654 ) ;
  assign n11657 = ( n11547 & ~n11655 ) | ( n11547 & n11656 ) | ( ~n11655 & n11656 ) ;
  assign n11658 = ( n11412 & n11537 ) | ( n11412 & n11657 ) | ( n11537 & n11657 ) ;
  assign n11659 = ( n11412 & ~n11537 ) | ( n11412 & n11657 ) | ( ~n11537 & n11657 ) ;
  assign n11660 = ( n11537 & ~n11658 ) | ( n11537 & n11659 ) | ( ~n11658 & n11659 ) ;
  assign n11661 = ( n11415 & n11527 ) | ( n11415 & n11660 ) | ( n11527 & n11660 ) ;
  assign n11662 = ( n11415 & ~n11527 ) | ( n11415 & n11660 ) | ( ~n11527 & n11660 ) ;
  assign n11663 = ( n11527 & ~n11661 ) | ( n11527 & n11662 ) | ( ~n11661 & n11662 ) ;
  assign n11664 = ( n11418 & n11517 ) | ( n11418 & n11663 ) | ( n11517 & n11663 ) ;
  assign n11665 = ( n11418 & ~n11517 ) | ( n11418 & n11663 ) | ( ~n11517 & n11663 ) ;
  assign n11666 = ( n11517 & ~n11664 ) | ( n11517 & n11665 ) | ( ~n11664 & n11665 ) ;
  assign n11667 = ( n11421 & n11507 ) | ( n11421 & n11666 ) | ( n11507 & n11666 ) ;
  assign n11668 = ( n11421 & ~n11507 ) | ( n11421 & n11666 ) | ( ~n11507 & n11666 ) ;
  assign n11669 = ( n11507 & ~n11667 ) | ( n11507 & n11668 ) | ( ~n11667 & n11668 ) ;
  assign n11670 = ( n11424 & n11497 ) | ( n11424 & n11669 ) | ( n11497 & n11669 ) ;
  assign n11671 = ( n11424 & ~n11497 ) | ( n11424 & n11669 ) | ( ~n11497 & n11669 ) ;
  assign n11672 = ( n11497 & ~n11670 ) | ( n11497 & n11671 ) | ( ~n11670 & n11671 ) ;
  assign n11673 = ( n11427 & n11487 ) | ( n11427 & n11672 ) | ( n11487 & n11672 ) ;
  assign n11674 = ( n11427 & ~n11487 ) | ( n11427 & n11672 ) | ( ~n11487 & n11672 ) ;
  assign n11675 = ( n11487 & ~n11673 ) | ( n11487 & n11674 ) | ( ~n11673 & n11674 ) ;
  assign n11676 = ( n11430 & n11477 ) | ( n11430 & n11675 ) | ( n11477 & n11675 ) ;
  assign n11677 = ( n11430 & ~n11477 ) | ( n11430 & n11675 ) | ( ~n11477 & n11675 ) ;
  assign n11678 = ( n11477 & ~n11676 ) | ( n11477 & n11677 ) | ( ~n11676 & n11677 ) ;
  assign n11679 = ( n11433 & n11467 ) | ( n11433 & n11678 ) | ( n11467 & n11678 ) ;
  assign n11680 = ( n11433 & ~n11467 ) | ( n11433 & n11678 ) | ( ~n11467 & n11678 ) ;
  assign n11681 = ( n11467 & ~n11679 ) | ( n11467 & n11680 ) | ( ~n11679 & n11680 ) ;
  assign n11682 = ( n11436 & n11457 ) | ( n11436 & n11681 ) | ( n11457 & n11681 ) ;
  assign n11683 = ( n11436 & ~n11457 ) | ( n11436 & n11681 ) | ( ~n11457 & n11681 ) ;
  assign n11684 = ( n11457 & ~n11682 ) | ( n11457 & n11683 ) | ( ~n11682 & n11683 ) ;
  assign n11685 = x127 & n359 ;
  assign n11686 = n301 | n11685 ;
  assign n11687 = ( n9865 & n11685 ) | ( n9865 & n11686 ) | ( n11685 & n11686 ) ;
  assign n11688 = x8 & ~n11687 ;
  assign n11689 = ~x8 & n11687 ;
  assign n11690 = n11688 | n11689 ;
  assign n11691 = ( n11439 & n11684 ) | ( n11439 & n11690 ) | ( n11684 & n11690 ) ;
  assign n11692 = ( n11439 & ~n11684 ) | ( n11439 & n11690 ) | ( ~n11684 & n11690 ) ;
  assign n11693 = ( n11684 & ~n11691 ) | ( n11684 & n11692 ) | ( ~n11691 & n11692 ) ;
  assign n11694 = ( n11442 & ~n11446 ) | ( n11442 & n11693 ) | ( ~n11446 & n11693 ) ;
  assign n11695 = ( n11442 & n11446 ) | ( n11442 & n11693 ) | ( n11446 & n11693 ) ;
  assign n11696 = ( n11446 & n11694 ) | ( n11446 & ~n11695 ) | ( n11694 & ~n11695 ) ;
  assign n11697 = n449 & n9576 ;
  assign n11698 = x11 & n11697 ;
  assign n11699 = x127 & n456 ;
  assign n11700 = x126 & n453 ;
  assign n11701 = n11699 | n11700 ;
  assign n11702 = x125 & n536 ;
  assign n11703 = n11701 | n11702 ;
  assign n11704 = ( ~x11 & n11697 ) | ( ~x11 & n11703 ) | ( n11697 & n11703 ) ;
  assign n11705 = x11 & ~n11703 ;
  assign n11706 = ( ~n11698 & n11704 ) | ( ~n11698 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11707 = n649 & n8729 ;
  assign n11708 = x14 & n11707 ;
  assign n11709 = x124 & n656 ;
  assign n11710 = x123 & n653 ;
  assign n11711 = n11709 | n11710 ;
  assign n11712 = x122 & n744 ;
  assign n11713 = n11711 | n11712 ;
  assign n11714 = ( ~x14 & n11707 ) | ( ~x14 & n11713 ) | ( n11707 & n11713 ) ;
  assign n11715 = x14 & ~n11713 ;
  assign n11716 = ( ~n11708 & n11714 ) | ( ~n11708 & n11715 ) | ( n11714 & n11715 ) ;
  assign n11717 = n874 & n7696 ;
  assign n11718 = x17 & n11717 ;
  assign n11719 = x121 & n881 ;
  assign n11720 = x120 & n878 ;
  assign n11721 = n11719 | n11720 ;
  assign n11722 = x119 & n959 ;
  assign n11723 = n11721 | n11722 ;
  assign n11724 = ( ~x17 & n11717 ) | ( ~x17 & n11723 ) | ( n11717 & n11723 ) ;
  assign n11725 = x17 & ~n11723 ;
  assign n11726 = ( ~n11718 & n11724 ) | ( ~n11718 & n11725 ) | ( n11724 & n11725 ) ;
  assign n11727 = n1146 & n6940 ;
  assign n11728 = x20 & n11727 ;
  assign n11729 = x118 & n1153 ;
  assign n11730 = x117 & n1150 ;
  assign n11731 = n11729 | n11730 ;
  assign n11732 = x116 & n1217 ;
  assign n11733 = n11731 | n11732 ;
  assign n11734 = ( ~x20 & n11727 ) | ( ~x20 & n11733 ) | ( n11727 & n11733 ) ;
  assign n11735 = x20 & ~n11733 ;
  assign n11736 = ( ~n11728 & n11734 ) | ( ~n11728 & n11735 ) | ( n11734 & n11735 ) ;
  assign n11737 = n1427 & n6446 ;
  assign n11738 = x23 & n11737 ;
  assign n11739 = x115 & n1434 ;
  assign n11740 = x114 & n1431 ;
  assign n11741 = n11739 | n11740 ;
  assign n11742 = x113 & n1531 ;
  assign n11743 = n11741 | n11742 ;
  assign n11744 = ( ~x23 & n11737 ) | ( ~x23 & n11743 ) | ( n11737 & n11743 ) ;
  assign n11745 = x23 & ~n11743 ;
  assign n11746 = ( ~n11738 & n11744 ) | ( ~n11738 & n11745 ) | ( n11744 & n11745 ) ;
  assign n11747 = n1755 & n5558 ;
  assign n11748 = x26 & n11747 ;
  assign n11749 = x112 & n1762 ;
  assign n11750 = x111 & n1759 ;
  assign n11751 = n11749 | n11750 ;
  assign n11752 = x110 & n1895 ;
  assign n11753 = n11751 | n11752 ;
  assign n11754 = ( ~x26 & n11747 ) | ( ~x26 & n11753 ) | ( n11747 & n11753 ) ;
  assign n11755 = x26 & ~n11753 ;
  assign n11756 = ( ~n11748 & n11754 ) | ( ~n11748 & n11755 ) | ( n11754 & n11755 ) ;
  assign n11757 = n2137 & n4930 ;
  assign n11758 = x29 & n11757 ;
  assign n11759 = x109 & n2144 ;
  assign n11760 = x108 & n2141 ;
  assign n11761 = n11759 | n11760 ;
  assign n11762 = x107 & n2267 ;
  assign n11763 = n11761 | n11762 ;
  assign n11764 = ( ~x29 & n11757 ) | ( ~x29 & n11763 ) | ( n11757 & n11763 ) ;
  assign n11765 = x29 & ~n11763 ;
  assign n11766 = ( ~n11758 & n11764 ) | ( ~n11758 & n11765 ) | ( n11764 & n11765 ) ;
  assign n11767 = n2545 & n4331 ;
  assign n11768 = x32 & n11767 ;
  assign n11769 = x106 & n2552 ;
  assign n11770 = x105 & n2549 ;
  assign n11771 = n11769 | n11770 ;
  assign n11772 = x104 & n2696 ;
  assign n11773 = n11771 | n11772 ;
  assign n11774 = ( ~x32 & n11767 ) | ( ~x32 & n11773 ) | ( n11767 & n11773 ) ;
  assign n11775 = x32 & ~n11773 ;
  assign n11776 = ( ~n11768 & n11774 ) | ( ~n11768 & n11775 ) | ( n11774 & n11775 ) ;
  assign n11777 = n2982 & n3941 ;
  assign n11778 = x35 & n11777 ;
  assign n11779 = x103 & n2989 ;
  assign n11780 = x102 & n2986 ;
  assign n11781 = n11779 | n11780 ;
  assign n11782 = x101 & n3159 ;
  assign n11783 = n11781 | n11782 ;
  assign n11784 = ( ~x35 & n11777 ) | ( ~x35 & n11783 ) | ( n11777 & n11783 ) ;
  assign n11785 = x35 & ~n11783 ;
  assign n11786 = ( ~n11778 & n11784 ) | ( ~n11778 & n11785 ) | ( n11784 & n11785 ) ;
  assign n11787 = n3264 & n3492 ;
  assign n11788 = x38 & n11787 ;
  assign n11789 = x100 & n3499 ;
  assign n11790 = x99 & n3496 ;
  assign n11791 = n11789 | n11790 ;
  assign n11792 = x98 & n3662 ;
  assign n11793 = n11791 | n11792 ;
  assign n11794 = ( ~x38 & n11787 ) | ( ~x38 & n11793 ) | ( n11787 & n11793 ) ;
  assign n11795 = x38 & ~n11793 ;
  assign n11796 = ( ~n11788 & n11794 ) | ( ~n11788 & n11795 ) | ( n11794 & n11795 ) ;
  assign n11797 = n2788 & n4020 ;
  assign n11798 = x41 & n11797 ;
  assign n11799 = x97 & n4027 ;
  assign n11800 = x96 & n4024 ;
  assign n11801 = n11799 | n11800 ;
  assign n11802 = x95 & n4223 ;
  assign n11803 = n11801 | n11802 ;
  assign n11804 = ( ~x41 & n11797 ) | ( ~x41 & n11803 ) | ( n11797 & n11803 ) ;
  assign n11805 = x41 & ~n11803 ;
  assign n11806 = ( ~n11798 & n11804 ) | ( ~n11798 & n11805 ) | ( n11804 & n11805 ) ;
  assign n11807 = n2476 & n4625 ;
  assign n11808 = x44 & n11807 ;
  assign n11809 = x94 & n4791 ;
  assign n11810 = x93 & n4621 ;
  assign n11811 = n11809 | n11810 ;
  assign n11812 = x92 & n4795 ;
  assign n11813 = n11811 | n11812 ;
  assign n11814 = ( ~x44 & n11807 ) | ( ~x44 & n11813 ) | ( n11807 & n11813 ) ;
  assign n11815 = x44 & ~n11813 ;
  assign n11816 = ( ~n11808 & n11814 ) | ( ~n11808 & n11815 ) | ( n11814 & n11815 ) ;
  assign n11817 = n1959 & n5223 ;
  assign n11818 = x47 & n11817 ;
  assign n11819 = x91 & n5230 ;
  assign n11820 = x90 & n5227 ;
  assign n11821 = n11819 | n11820 ;
  assign n11822 = x89 & n5434 ;
  assign n11823 = n11821 | n11822 ;
  assign n11824 = ( ~x47 & n11817 ) | ( ~x47 & n11823 ) | ( n11817 & n11823 ) ;
  assign n11825 = x47 & ~n11823 ;
  assign n11826 = ( ~n11818 & n11824 ) | ( ~n11818 & n11825 ) | ( n11824 & n11825 ) ;
  assign n11827 = n1602 & n5858 ;
  assign n11828 = x50 & n11827 ;
  assign n11829 = x88 & n5865 ;
  assign n11830 = x87 & n5862 ;
  assign n11831 = n11829 | n11830 ;
  assign n11832 = x86 & n6092 ;
  assign n11833 = n11831 | n11832 ;
  assign n11834 = ( ~x50 & n11827 ) | ( ~x50 & n11833 ) | ( n11827 & n11833 ) ;
  assign n11835 = x50 & ~n11833 ;
  assign n11836 = ( ~n11828 & n11834 ) | ( ~n11828 & n11835 ) | ( n11834 & n11835 ) ;
  assign n11837 = n1368 & n6546 ;
  assign n11838 = x53 & n11837 ;
  assign n11839 = x85 & n6553 ;
  assign n11840 = x84 & n6550 ;
  assign n11841 = n11839 | n11840 ;
  assign n11842 = x83 & n6787 ;
  assign n11843 = n11841 | n11842 ;
  assign n11844 = ( ~x53 & n11837 ) | ( ~x53 & n11843 ) | ( n11837 & n11843 ) ;
  assign n11845 = x53 & ~n11843 ;
  assign n11846 = ( ~n11838 & n11844 ) | ( ~n11838 & n11845 ) | ( n11844 & n11845 ) ;
  assign n11847 = n823 & n8067 ;
  assign n11848 = x59 & n11847 ;
  assign n11849 = x79 & n8074 ;
  assign n11850 = x78 & n8071 ;
  assign n11851 = n11849 | n11850 ;
  assign n11852 = x77 & n8298 ;
  assign n11853 = n11851 | n11852 ;
  assign n11854 = ( ~x59 & n11847 ) | ( ~x59 & n11853 ) | ( n11847 & n11853 ) ;
  assign n11855 = x59 & ~n11853 ;
  assign n11856 = ( ~n11848 & n11854 ) | ( ~n11848 & n11855 ) | ( n11854 & n11855 ) ;
  assign n11857 = n565 & n8859 ;
  assign n11858 = x62 & n11857 ;
  assign n11859 = x76 & n8866 ;
  assign n11860 = x75 & n8863 ;
  assign n11861 = n11859 | n11860 ;
  assign n11862 = x74 & n9125 ;
  assign n11863 = n11861 | n11862 ;
  assign n11864 = ( ~x62 & n11857 ) | ( ~x62 & n11863 ) | ( n11857 & n11863 ) ;
  assign n11865 = x62 & ~n11863 ;
  assign n11866 = ( ~n11858 & n11864 ) | ( ~n11858 & n11865 ) | ( n11864 & n11865 ) ;
  assign n11867 = ( x62 & x63 ) | ( x62 & x73 ) | ( x63 & x73 ) ;
  assign n11868 = ( x62 & x72 ) | ( x62 & ~n9394 ) | ( x72 & ~n9394 ) ;
  assign n11869 = ( x72 & n11867 ) | ( x72 & ~n11868 ) | ( n11867 & ~n11868 ) ;
  assign n11870 = ( x8 & n11620 ) | ( x8 & n11869 ) | ( n11620 & n11869 ) ;
  assign n11871 = ( ~x8 & n11620 ) | ( ~x8 & n11869 ) | ( n11620 & n11869 ) ;
  assign n11872 = ( x8 & ~n11870 ) | ( x8 & n11871 ) | ( ~n11870 & n11871 ) ;
  assign n11873 = ( n11622 & ~n11866 ) | ( n11622 & n11872 ) | ( ~n11866 & n11872 ) ;
  assign n11874 = ( n11622 & n11866 ) | ( n11622 & n11872 ) | ( n11866 & n11872 ) ;
  assign n11875 = ( n11866 & n11873 ) | ( n11866 & ~n11874 ) | ( n11873 & ~n11874 ) ;
  assign n11876 = ( n11624 & n11856 ) | ( n11624 & n11875 ) | ( n11856 & n11875 ) ;
  assign n11877 = ( ~n11624 & n11856 ) | ( ~n11624 & n11875 ) | ( n11856 & n11875 ) ;
  assign n11878 = ( n11624 & ~n11876 ) | ( n11624 & n11877 ) | ( ~n11876 & n11877 ) ;
  assign n11879 = n1006 & n7277 ;
  assign n11880 = x56 & n11879 ;
  assign n11881 = x82 & n7545 ;
  assign n11882 = x81 & n7273 ;
  assign n11883 = n11881 | n11882 ;
  assign n11884 = x80 & n7552 ;
  assign n11885 = n11883 | n11884 ;
  assign n11886 = ( ~x56 & n11879 ) | ( ~x56 & n11885 ) | ( n11879 & n11885 ) ;
  assign n11887 = x56 & ~n11885 ;
  assign n11888 = ( ~n11880 & n11886 ) | ( ~n11880 & n11887 ) | ( n11886 & n11887 ) ;
  assign n11889 = ( n11637 & n11878 ) | ( n11637 & n11888 ) | ( n11878 & n11888 ) ;
  assign n11890 = ( n11637 & ~n11878 ) | ( n11637 & n11888 ) | ( ~n11878 & n11888 ) ;
  assign n11891 = ( n11878 & ~n11889 ) | ( n11878 & n11890 ) | ( ~n11889 & n11890 ) ;
  assign n11892 = ( n11641 & n11846 ) | ( n11641 & n11891 ) | ( n11846 & n11891 ) ;
  assign n11893 = ( n11641 & ~n11846 ) | ( n11641 & n11891 ) | ( ~n11846 & n11891 ) ;
  assign n11894 = ( n11846 & ~n11892 ) | ( n11846 & n11893 ) | ( ~n11892 & n11893 ) ;
  assign n11895 = ( n11643 & n11836 ) | ( n11643 & n11894 ) | ( n11836 & n11894 ) ;
  assign n11896 = ( ~n11643 & n11836 ) | ( ~n11643 & n11894 ) | ( n11836 & n11894 ) ;
  assign n11897 = ( n11643 & ~n11895 ) | ( n11643 & n11896 ) | ( ~n11895 & n11896 ) ;
  assign n11898 = ( n11646 & n11826 ) | ( n11646 & n11897 ) | ( n11826 & n11897 ) ;
  assign n11899 = ( n11646 & ~n11826 ) | ( n11646 & n11897 ) | ( ~n11826 & n11897 ) ;
  assign n11900 = ( n11826 & ~n11898 ) | ( n11826 & n11899 ) | ( ~n11898 & n11899 ) ;
  assign n11901 = ( n11649 & n11816 ) | ( n11649 & n11900 ) | ( n11816 & n11900 ) ;
  assign n11902 = ( ~n11649 & n11816 ) | ( ~n11649 & n11900 ) | ( n11816 & n11900 ) ;
  assign n11903 = ( n11649 & ~n11901 ) | ( n11649 & n11902 ) | ( ~n11901 & n11902 ) ;
  assign n11904 = ( n11652 & n11806 ) | ( n11652 & n11903 ) | ( n11806 & n11903 ) ;
  assign n11905 = ( ~n11652 & n11806 ) | ( ~n11652 & n11903 ) | ( n11806 & n11903 ) ;
  assign n11906 = ( n11652 & ~n11904 ) | ( n11652 & n11905 ) | ( ~n11904 & n11905 ) ;
  assign n11907 = ( n11655 & n11796 ) | ( n11655 & n11906 ) | ( n11796 & n11906 ) ;
  assign n11908 = ( ~n11655 & n11796 ) | ( ~n11655 & n11906 ) | ( n11796 & n11906 ) ;
  assign n11909 = ( n11655 & ~n11907 ) | ( n11655 & n11908 ) | ( ~n11907 & n11908 ) ;
  assign n11910 = ( n11658 & n11786 ) | ( n11658 & n11909 ) | ( n11786 & n11909 ) ;
  assign n11911 = ( n11658 & ~n11786 ) | ( n11658 & n11909 ) | ( ~n11786 & n11909 ) ;
  assign n11912 = ( n11786 & ~n11910 ) | ( n11786 & n11911 ) | ( ~n11910 & n11911 ) ;
  assign n11913 = ( n11661 & n11776 ) | ( n11661 & n11912 ) | ( n11776 & n11912 ) ;
  assign n11914 = ( ~n11661 & n11776 ) | ( ~n11661 & n11912 ) | ( n11776 & n11912 ) ;
  assign n11915 = ( n11661 & ~n11913 ) | ( n11661 & n11914 ) | ( ~n11913 & n11914 ) ;
  assign n11916 = ( n11664 & n11766 ) | ( n11664 & n11915 ) | ( n11766 & n11915 ) ;
  assign n11917 = ( ~n11664 & n11766 ) | ( ~n11664 & n11915 ) | ( n11766 & n11915 ) ;
  assign n11918 = ( n11664 & ~n11916 ) | ( n11664 & n11917 ) | ( ~n11916 & n11917 ) ;
  assign n11919 = ( n11667 & n11756 ) | ( n11667 & n11918 ) | ( n11756 & n11918 ) ;
  assign n11920 = ( n11667 & ~n11756 ) | ( n11667 & n11918 ) | ( ~n11756 & n11918 ) ;
  assign n11921 = ( n11756 & ~n11919 ) | ( n11756 & n11920 ) | ( ~n11919 & n11920 ) ;
  assign n11922 = ( n11670 & n11746 ) | ( n11670 & n11921 ) | ( n11746 & n11921 ) ;
  assign n11923 = ( ~n11670 & n11746 ) | ( ~n11670 & n11921 ) | ( n11746 & n11921 ) ;
  assign n11924 = ( n11670 & ~n11922 ) | ( n11670 & n11923 ) | ( ~n11922 & n11923 ) ;
  assign n11925 = ( n11673 & n11736 ) | ( n11673 & n11924 ) | ( n11736 & n11924 ) ;
  assign n11926 = ( ~n11673 & n11736 ) | ( ~n11673 & n11924 ) | ( n11736 & n11924 ) ;
  assign n11927 = ( n11673 & ~n11925 ) | ( n11673 & n11926 ) | ( ~n11925 & n11926 ) ;
  assign n11928 = ( n11676 & n11726 ) | ( n11676 & n11927 ) | ( n11726 & n11927 ) ;
  assign n11929 = ( n11676 & ~n11726 ) | ( n11676 & n11927 ) | ( ~n11726 & n11927 ) ;
  assign n11930 = ( n11726 & ~n11928 ) | ( n11726 & n11929 ) | ( ~n11928 & n11929 ) ;
  assign n11931 = ( n11679 & n11716 ) | ( n11679 & n11930 ) | ( n11716 & n11930 ) ;
  assign n11932 = ( ~n11679 & n11716 ) | ( ~n11679 & n11930 ) | ( n11716 & n11930 ) ;
  assign n11933 = ( n11679 & ~n11931 ) | ( n11679 & n11932 ) | ( ~n11931 & n11932 ) ;
  assign n11934 = ( n11682 & n11706 ) | ( n11682 & n11933 ) | ( n11706 & n11933 ) ;
  assign n11935 = ( ~n11682 & n11706 ) | ( ~n11682 & n11933 ) | ( n11706 & n11933 ) ;
  assign n11936 = ( n11682 & ~n11934 ) | ( n11682 & n11935 ) | ( ~n11934 & n11935 ) ;
  assign n11937 = ( n11691 & n11695 ) | ( n11691 & n11936 ) | ( n11695 & n11936 ) ;
  assign n11938 = ( n11691 & ~n11695 ) | ( n11691 & n11936 ) | ( ~n11695 & n11936 ) ;
  assign n11939 = ( n11695 & ~n11937 ) | ( n11695 & n11938 ) | ( ~n11937 & n11938 ) ;
  assign n11940 = x127 & n453 ;
  assign n11941 = n449 | n11940 ;
  assign n11942 = ( n9867 & n11940 ) | ( n9867 & n11941 ) | ( n11940 & n11941 ) ;
  assign n11943 = x126 & n536 ;
  assign n11944 = ( ~x11 & n11942 ) | ( ~x11 & n11943 ) | ( n11942 & n11943 ) ;
  assign n11945 = ( x11 & ~n11942 ) | ( x11 & n11943 ) | ( ~n11942 & n11943 ) ;
  assign n11946 = ~n11943 & n11945 ;
  assign n11947 = n11944 | n11946 ;
  assign n11948 = n649 & n9009 ;
  assign n11949 = x14 & n11948 ;
  assign n11950 = x125 & n656 ;
  assign n11951 = x124 & n653 ;
  assign n11952 = n11950 | n11951 ;
  assign n11953 = x123 & n744 ;
  assign n11954 = n11952 | n11953 ;
  assign n11955 = ( ~x14 & n11948 ) | ( ~x14 & n11954 ) | ( n11948 & n11954 ) ;
  assign n11956 = x14 & ~n11954 ;
  assign n11957 = ( ~n11949 & n11955 ) | ( ~n11949 & n11956 ) | ( n11955 & n11956 ) ;
  assign n11958 = n874 & n8207 ;
  assign n11959 = x17 & n11958 ;
  assign n11960 = x122 & n881 ;
  assign n11961 = x121 & n878 ;
  assign n11962 = n11960 | n11961 ;
  assign n11963 = x120 & n959 ;
  assign n11964 = n11962 | n11963 ;
  assign n11965 = ( ~x17 & n11958 ) | ( ~x17 & n11964 ) | ( n11958 & n11964 ) ;
  assign n11966 = x17 & ~n11964 ;
  assign n11967 = ( ~n11959 & n11965 ) | ( ~n11959 & n11966 ) | ( n11965 & n11966 ) ;
  assign n11968 = n1146 & n7181 ;
  assign n11969 = x20 & n11968 ;
  assign n11970 = x119 & n1153 ;
  assign n11971 = x118 & n1150 ;
  assign n11972 = n11970 | n11971 ;
  assign n11973 = x117 & n1217 ;
  assign n11974 = n11972 | n11973 ;
  assign n11975 = ( ~x20 & n11968 ) | ( ~x20 & n11974 ) | ( n11968 & n11974 ) ;
  assign n11976 = x20 & ~n11974 ;
  assign n11977 = ( ~n11969 & n11975 ) | ( ~n11969 & n11976 ) | ( n11975 & n11976 ) ;
  assign n11978 = n1427 & n6462 ;
  assign n11979 = x23 & n11978 ;
  assign n11980 = x116 & n1434 ;
  assign n11981 = x115 & n1431 ;
  assign n11982 = n11980 | n11981 ;
  assign n11983 = x114 & n1531 ;
  assign n11984 = n11982 | n11983 ;
  assign n11985 = ( ~x23 & n11978 ) | ( ~x23 & n11984 ) | ( n11978 & n11984 ) ;
  assign n11986 = x23 & ~n11984 ;
  assign n11987 = ( ~n11979 & n11985 ) | ( ~n11979 & n11986 ) | ( n11985 & n11986 ) ;
  assign n11988 = n1755 & n5774 ;
  assign n11989 = x26 & n11988 ;
  assign n11990 = x113 & n1762 ;
  assign n11991 = x112 & n1759 ;
  assign n11992 = n11990 | n11991 ;
  assign n11993 = x111 & n1895 ;
  assign n11994 = n11992 | n11993 ;
  assign n11995 = ( ~x26 & n11988 ) | ( ~x26 & n11994 ) | ( n11988 & n11994 ) ;
  assign n11996 = x26 & ~n11994 ;
  assign n11997 = ( ~n11989 & n11995 ) | ( ~n11989 & n11996 ) | ( n11995 & n11996 ) ;
  assign n11998 = n2137 & n5331 ;
  assign n11999 = x29 & n11998 ;
  assign n12000 = x110 & n2144 ;
  assign n12001 = x109 & n2141 ;
  assign n12002 = n12000 | n12001 ;
  assign n12003 = x108 & n2267 ;
  assign n12004 = n12002 | n12003 ;
  assign n12005 = ( ~x29 & n11998 ) | ( ~x29 & n12004 ) | ( n11998 & n12004 ) ;
  assign n12006 = x29 & ~n12004 ;
  assign n12007 = ( ~n11999 & n12005 ) | ( ~n11999 & n12006 ) | ( n12005 & n12006 ) ;
  assign n12008 = n2545 & n4523 ;
  assign n12009 = x32 & n12008 ;
  assign n12010 = x107 & n2552 ;
  assign n12011 = x106 & n2549 ;
  assign n12012 = n12010 | n12011 ;
  assign n12013 = x105 & n2696 ;
  assign n12014 = n12012 | n12013 ;
  assign n12015 = ( ~x32 & n12008 ) | ( ~x32 & n12014 ) | ( n12008 & n12014 ) ;
  assign n12016 = x32 & ~n12014 ;
  assign n12017 = ( ~n12009 & n12015 ) | ( ~n12009 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12018 = n2982 & n3957 ;
  assign n12019 = x35 & n12018 ;
  assign n12020 = x104 & n2989 ;
  assign n12021 = x103 & n2986 ;
  assign n12022 = n12020 | n12021 ;
  assign n12023 = x102 & n3159 ;
  assign n12024 = n12022 | n12023 ;
  assign n12025 = ( ~x35 & n12018 ) | ( ~x35 & n12024 ) | ( n12018 & n12024 ) ;
  assign n12026 = x35 & ~n12024 ;
  assign n12027 = ( ~n12019 & n12025 ) | ( ~n12019 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12028 = n3492 & n3591 ;
  assign n12029 = x38 & n12028 ;
  assign n12030 = x101 & n3499 ;
  assign n12031 = x100 & n3496 ;
  assign n12032 = n12030 | n12031 ;
  assign n12033 = x99 & n3662 ;
  assign n12034 = n12032 | n12033 ;
  assign n12035 = ( ~x38 & n12028 ) | ( ~x38 & n12034 ) | ( n12028 & n12034 ) ;
  assign n12036 = x38 & ~n12034 ;
  assign n12037 = ( ~n12029 & n12035 ) | ( ~n12029 & n12036 ) | ( n12035 & n12036 ) ;
  assign n12038 = n2939 & n4020 ;
  assign n12039 = x41 & n12038 ;
  assign n12040 = x98 & n4027 ;
  assign n12041 = x97 & n4024 ;
  assign n12042 = n12040 | n12041 ;
  assign n12043 = x96 & n4223 ;
  assign n12044 = n12042 | n12043 ;
  assign n12045 = ( ~x41 & n12038 ) | ( ~x41 & n12044 ) | ( n12038 & n12044 ) ;
  assign n12046 = x41 & ~n12044 ;
  assign n12047 = ( ~n12039 & n12045 ) | ( ~n12039 & n12046 ) | ( n12045 & n12046 ) ;
  assign n12048 = x94 & n4621 ;
  assign n12049 = x93 | n12048 ;
  assign n12050 = ( n4795 & n12048 ) | ( n4795 & n12049 ) | ( n12048 & n12049 ) ;
  assign n12051 = n2492 & n4625 ;
  assign n12052 = n12050 | n12051 ;
  assign n12053 = x95 & n4791 ;
  assign n12054 = ( ~x44 & n12052 ) | ( ~x44 & n12053 ) | ( n12052 & n12053 ) ;
  assign n12055 = ( x44 & ~n12052 ) | ( x44 & n12053 ) | ( ~n12052 & n12053 ) ;
  assign n12056 = ~n12053 & n12055 ;
  assign n12057 = n12054 | n12056 ;
  assign n12058 = n2083 & n5223 ;
  assign n12059 = x47 & n12058 ;
  assign n12060 = x92 & n5230 ;
  assign n12061 = x91 & n5227 ;
  assign n12062 = n12060 | n12061 ;
  assign n12063 = x90 & n5434 ;
  assign n12064 = n12062 | n12063 ;
  assign n12065 = ( ~x47 & n12058 ) | ( ~x47 & n12064 ) | ( n12058 & n12064 ) ;
  assign n12066 = x47 & ~n12064 ;
  assign n12067 = ( ~n12059 & n12065 ) | ( ~n12059 & n12066 ) | ( n12065 & n12066 ) ;
  assign n12068 = n1822 & n5858 ;
  assign n12069 = x50 & n12068 ;
  assign n12070 = x89 & n5865 ;
  assign n12071 = x88 & n5862 ;
  assign n12072 = n12070 | n12071 ;
  assign n12073 = x87 & n6092 ;
  assign n12074 = n12072 | n12073 ;
  assign n12075 = ( ~x50 & n12068 ) | ( ~x50 & n12074 ) | ( n12068 & n12074 ) ;
  assign n12076 = x50 & ~n12074 ;
  assign n12077 = ( ~n12069 & n12075 ) | ( ~n12069 & n12076 ) | ( n12075 & n12076 ) ;
  assign n12078 = n1384 & n6546 ;
  assign n12079 = x53 & n12078 ;
  assign n12080 = x86 & n6553 ;
  assign n12081 = x85 & n6550 ;
  assign n12082 = n12080 | n12081 ;
  assign n12083 = x84 & n6787 ;
  assign n12084 = n12082 | n12083 ;
  assign n12085 = ( ~x53 & n12078 ) | ( ~x53 & n12084 ) | ( n12078 & n12084 ) ;
  assign n12086 = x53 & ~n12084 ;
  assign n12087 = ( ~n12079 & n12085 ) | ( ~n12079 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12088 = n1093 & n7277 ;
  assign n12089 = x56 & n12088 ;
  assign n12090 = x83 & n7545 ;
  assign n12091 = x82 & n7273 ;
  assign n12092 = n12090 | n12091 ;
  assign n12093 = x81 & n7552 ;
  assign n12094 = n12092 | n12093 ;
  assign n12095 = ( ~x56 & n12088 ) | ( ~x56 & n12094 ) | ( n12088 & n12094 ) ;
  assign n12096 = x56 & ~n12094 ;
  assign n12097 = ( ~n12089 & n12095 ) | ( ~n12089 & n12096 ) | ( n12095 & n12096 ) ;
  assign n12098 = n840 & n8067 ;
  assign n12099 = x59 & n12098 ;
  assign n12100 = x80 & n8074 ;
  assign n12101 = x79 & n8071 ;
  assign n12102 = n12100 | n12101 ;
  assign n12103 = x78 & n8298 ;
  assign n12104 = n12102 | n12103 ;
  assign n12105 = ( ~x59 & n12098 ) | ( ~x59 & n12104 ) | ( n12098 & n12104 ) ;
  assign n12106 = x59 & ~n12104 ;
  assign n12107 = ( ~n12099 & n12105 ) | ( ~n12099 & n12106 ) | ( n12105 & n12106 ) ;
  assign n12108 = ( x62 & x63 ) | ( x62 & x74 ) | ( x63 & x74 ) ;
  assign n12109 = ( x62 & x73 ) | ( x62 & ~n9394 ) | ( x73 & ~n9394 ) ;
  assign n12110 = ( x73 & n12108 ) | ( x73 & ~n12109 ) | ( n12108 & ~n12109 ) ;
  assign n12111 = n626 & n8859 ;
  assign n12112 = x62 & n12111 ;
  assign n12113 = x77 & n8866 ;
  assign n12114 = x76 & n8863 ;
  assign n12115 = n12113 | n12114 ;
  assign n12116 = x75 & n9125 ;
  assign n12117 = n12115 | n12116 ;
  assign n12118 = ( ~x62 & n12111 ) | ( ~x62 & n12117 ) | ( n12111 & n12117 ) ;
  assign n12119 = x62 & ~n12117 ;
  assign n12120 = ( ~n12112 & n12118 ) | ( ~n12112 & n12119 ) | ( n12118 & n12119 ) ;
  assign n12121 = ( ~n11871 & n12110 ) | ( ~n11871 & n12120 ) | ( n12110 & n12120 ) ;
  assign n12122 = ( n11871 & n12110 ) | ( n11871 & ~n12120 ) | ( n12110 & ~n12120 ) ;
  assign n12123 = ( ~n12110 & n12121 ) | ( ~n12110 & n12122 ) | ( n12121 & n12122 ) ;
  assign n12124 = ( n11873 & ~n12107 ) | ( n11873 & n12123 ) | ( ~n12107 & n12123 ) ;
  assign n12125 = ( n11873 & n12107 ) | ( n11873 & n12123 ) | ( n12107 & n12123 ) ;
  assign n12126 = ( n12107 & n12124 ) | ( n12107 & ~n12125 ) | ( n12124 & ~n12125 ) ;
  assign n12127 = ( n11876 & n12097 ) | ( n11876 & n12126 ) | ( n12097 & n12126 ) ;
  assign n12128 = ( n11876 & ~n12097 ) | ( n11876 & n12126 ) | ( ~n12097 & n12126 ) ;
  assign n12129 = ( n12097 & ~n12127 ) | ( n12097 & n12128 ) | ( ~n12127 & n12128 ) ;
  assign n12130 = ( n11889 & n12087 ) | ( n11889 & n12129 ) | ( n12087 & n12129 ) ;
  assign n12131 = ( n11889 & ~n12087 ) | ( n11889 & n12129 ) | ( ~n12087 & n12129 ) ;
  assign n12132 = ( n12087 & ~n12130 ) | ( n12087 & n12131 ) | ( ~n12130 & n12131 ) ;
  assign n12133 = ( n11892 & n12077 ) | ( n11892 & n12132 ) | ( n12077 & n12132 ) ;
  assign n12134 = ( n11892 & ~n12077 ) | ( n11892 & n12132 ) | ( ~n12077 & n12132 ) ;
  assign n12135 = ( n12077 & ~n12133 ) | ( n12077 & n12134 ) | ( ~n12133 & n12134 ) ;
  assign n12136 = ( n11895 & n12067 ) | ( n11895 & n12135 ) | ( n12067 & n12135 ) ;
  assign n12137 = ( n11895 & ~n12067 ) | ( n11895 & n12135 ) | ( ~n12067 & n12135 ) ;
  assign n12138 = ( n12067 & ~n12136 ) | ( n12067 & n12137 ) | ( ~n12136 & n12137 ) ;
  assign n12139 = ( n11898 & n12057 ) | ( n11898 & n12138 ) | ( n12057 & n12138 ) ;
  assign n12140 = ( n11898 & ~n12057 ) | ( n11898 & n12138 ) | ( ~n12057 & n12138 ) ;
  assign n12141 = ( n12057 & ~n12139 ) | ( n12057 & n12140 ) | ( ~n12139 & n12140 ) ;
  assign n12142 = ( n11901 & n12047 ) | ( n11901 & n12141 ) | ( n12047 & n12141 ) ;
  assign n12143 = ( n11901 & ~n12047 ) | ( n11901 & n12141 ) | ( ~n12047 & n12141 ) ;
  assign n12144 = ( n12047 & ~n12142 ) | ( n12047 & n12143 ) | ( ~n12142 & n12143 ) ;
  assign n12145 = ( n11904 & n12037 ) | ( n11904 & n12144 ) | ( n12037 & n12144 ) ;
  assign n12146 = ( n11904 & ~n12037 ) | ( n11904 & n12144 ) | ( ~n12037 & n12144 ) ;
  assign n12147 = ( n12037 & ~n12145 ) | ( n12037 & n12146 ) | ( ~n12145 & n12146 ) ;
  assign n12148 = ( n11907 & n12027 ) | ( n11907 & n12147 ) | ( n12027 & n12147 ) ;
  assign n12149 = ( n11907 & ~n12027 ) | ( n11907 & n12147 ) | ( ~n12027 & n12147 ) ;
  assign n12150 = ( n12027 & ~n12148 ) | ( n12027 & n12149 ) | ( ~n12148 & n12149 ) ;
  assign n12151 = ( n11910 & n12017 ) | ( n11910 & n12150 ) | ( n12017 & n12150 ) ;
  assign n12152 = ( n11910 & ~n12017 ) | ( n11910 & n12150 ) | ( ~n12017 & n12150 ) ;
  assign n12153 = ( n12017 & ~n12151 ) | ( n12017 & n12152 ) | ( ~n12151 & n12152 ) ;
  assign n12154 = ( n11913 & n12007 ) | ( n11913 & n12153 ) | ( n12007 & n12153 ) ;
  assign n12155 = ( n11913 & ~n12007 ) | ( n11913 & n12153 ) | ( ~n12007 & n12153 ) ;
  assign n12156 = ( n12007 & ~n12154 ) | ( n12007 & n12155 ) | ( ~n12154 & n12155 ) ;
  assign n12157 = ( n11916 & n11997 ) | ( n11916 & n12156 ) | ( n11997 & n12156 ) ;
  assign n12158 = ( n11916 & ~n11997 ) | ( n11916 & n12156 ) | ( ~n11997 & n12156 ) ;
  assign n12159 = ( n11997 & ~n12157 ) | ( n11997 & n12158 ) | ( ~n12157 & n12158 ) ;
  assign n12160 = ( n11919 & n11987 ) | ( n11919 & n12159 ) | ( n11987 & n12159 ) ;
  assign n12161 = ( n11919 & ~n11987 ) | ( n11919 & n12159 ) | ( ~n11987 & n12159 ) ;
  assign n12162 = ( n11987 & ~n12160 ) | ( n11987 & n12161 ) | ( ~n12160 & n12161 ) ;
  assign n12163 = ( n11922 & n11977 ) | ( n11922 & n12162 ) | ( n11977 & n12162 ) ;
  assign n12164 = ( n11922 & ~n11977 ) | ( n11922 & n12162 ) | ( ~n11977 & n12162 ) ;
  assign n12165 = ( n11977 & ~n12163 ) | ( n11977 & n12164 ) | ( ~n12163 & n12164 ) ;
  assign n12166 = ( n11925 & n11967 ) | ( n11925 & n12165 ) | ( n11967 & n12165 ) ;
  assign n12167 = ( n11925 & ~n11967 ) | ( n11925 & n12165 ) | ( ~n11967 & n12165 ) ;
  assign n12168 = ( n11967 & ~n12166 ) | ( n11967 & n12167 ) | ( ~n12166 & n12167 ) ;
  assign n12169 = ( n11928 & n11957 ) | ( n11928 & n12168 ) | ( n11957 & n12168 ) ;
  assign n12170 = ( n11928 & ~n11957 ) | ( n11928 & n12168 ) | ( ~n11957 & n12168 ) ;
  assign n12171 = ( n11957 & ~n12169 ) | ( n11957 & n12170 ) | ( ~n12169 & n12170 ) ;
  assign n12172 = ( n11931 & n11947 ) | ( n11931 & n12171 ) | ( n11947 & n12171 ) ;
  assign n12173 = ( n11931 & ~n11947 ) | ( n11931 & n12171 ) | ( ~n11947 & n12171 ) ;
  assign n12174 = ( n11947 & ~n12172 ) | ( n11947 & n12173 ) | ( ~n12172 & n12173 ) ;
  assign n12175 = ( n11934 & ~n11937 ) | ( n11934 & n12174 ) | ( ~n11937 & n12174 ) ;
  assign n12176 = ( n11934 & n11937 ) | ( n11934 & n12174 ) | ( n11937 & n12174 ) ;
  assign n12177 = ( n11937 & n12175 ) | ( n11937 & ~n12176 ) | ( n12175 & ~n12176 ) ;
  assign n12178 = n649 & n9038 ;
  assign n12179 = x14 & n12178 ;
  assign n12180 = x126 & n656 ;
  assign n12181 = x125 & n653 ;
  assign n12182 = n12180 | n12181 ;
  assign n12183 = x124 & n744 ;
  assign n12184 = n12182 | n12183 ;
  assign n12185 = ( ~x14 & n12178 ) | ( ~x14 & n12184 ) | ( n12178 & n12184 ) ;
  assign n12186 = x14 & ~n12184 ;
  assign n12187 = ( ~n12179 & n12185 ) | ( ~n12179 & n12186 ) | ( n12185 & n12186 ) ;
  assign n12188 = n874 & n8461 ;
  assign n12189 = x17 & n12188 ;
  assign n12190 = x123 & n881 ;
  assign n12191 = x122 & n878 ;
  assign n12192 = n12190 | n12191 ;
  assign n12193 = x121 & n959 ;
  assign n12194 = n12192 | n12193 ;
  assign n12195 = ( ~x17 & n12188 ) | ( ~x17 & n12194 ) | ( n12188 & n12194 ) ;
  assign n12196 = x17 & ~n12194 ;
  assign n12197 = ( ~n12189 & n12195 ) | ( ~n12189 & n12196 ) | ( n12195 & n12196 ) ;
  assign n12198 = n1146 & n7444 ;
  assign n12199 = x20 & n12198 ;
  assign n12200 = x120 & n1153 ;
  assign n12201 = x119 & n1150 ;
  assign n12202 = n12200 | n12201 ;
  assign n12203 = x118 & n1217 ;
  assign n12204 = n12202 | n12203 ;
  assign n12205 = ( ~x20 & n12198 ) | ( ~x20 & n12204 ) | ( n12198 & n12204 ) ;
  assign n12206 = x20 & ~n12204 ;
  assign n12207 = ( ~n12199 & n12205 ) | ( ~n12199 & n12206 ) | ( n12205 & n12206 ) ;
  assign n12208 = n1427 & n6924 ;
  assign n12209 = x23 & n12208 ;
  assign n12210 = x117 & n1434 ;
  assign n12211 = x116 & n1431 ;
  assign n12212 = n12210 | n12211 ;
  assign n12213 = x115 & n1531 ;
  assign n12214 = n12212 | n12213 ;
  assign n12215 = ( ~x23 & n12208 ) | ( ~x23 & n12214 ) | ( n12208 & n12214 ) ;
  assign n12216 = x23 & ~n12214 ;
  assign n12217 = ( ~n12209 & n12215 ) | ( ~n12209 & n12216 ) | ( n12215 & n12216 ) ;
  assign n12218 = n1755 & n6002 ;
  assign n12219 = x26 & n12218 ;
  assign n12220 = x114 & n1762 ;
  assign n12221 = x113 & n1759 ;
  assign n12222 = n12220 | n12221 ;
  assign n12223 = x112 & n1895 ;
  assign n12224 = n12222 | n12223 ;
  assign n12225 = ( ~x26 & n12218 ) | ( ~x26 & n12224 ) | ( n12218 & n12224 ) ;
  assign n12226 = x26 & ~n12224 ;
  assign n12227 = ( ~n12219 & n12225 ) | ( ~n12219 & n12226 ) | ( n12225 & n12226 ) ;
  assign n12228 = n2137 & n5347 ;
  assign n12229 = x29 & n12228 ;
  assign n12230 = x111 & n2144 ;
  assign n12231 = x110 & n2141 ;
  assign n12232 = n12230 | n12231 ;
  assign n12233 = x109 & n2267 ;
  assign n12234 = n12232 | n12233 ;
  assign n12235 = ( ~x29 & n12228 ) | ( ~x29 & n12234 ) | ( n12228 & n12234 ) ;
  assign n12236 = x29 & ~n12234 ;
  assign n12237 = ( ~n12229 & n12235 ) | ( ~n12229 & n12236 ) | ( n12235 & n12236 ) ;
  assign n12238 = n2545 & n4914 ;
  assign n12239 = x32 & n12238 ;
  assign n12240 = x108 & n2552 ;
  assign n12241 = x107 & n2549 ;
  assign n12242 = n12240 | n12241 ;
  assign n12243 = x106 & n2696 ;
  assign n12244 = n12242 | n12243 ;
  assign n12245 = ( ~x32 & n12238 ) | ( ~x32 & n12244 ) | ( n12238 & n12244 ) ;
  assign n12246 = x32 & ~n12244 ;
  assign n12247 = ( ~n12239 & n12245 ) | ( ~n12239 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12248 = n2982 & n4145 ;
  assign n12249 = x35 & n12248 ;
  assign n12250 = x105 & n2989 ;
  assign n12251 = x104 & n2986 ;
  assign n12252 = n12250 | n12251 ;
  assign n12253 = x103 & n3159 ;
  assign n12254 = n12252 | n12253 ;
  assign n12255 = ( ~x35 & n12248 ) | ( ~x35 & n12254 ) | ( n12248 & n12254 ) ;
  assign n12256 = x35 & ~n12254 ;
  assign n12257 = ( ~n12249 & n12255 ) | ( ~n12249 & n12256 ) | ( n12255 & n12256 ) ;
  assign n12258 = n3492 & n3764 ;
  assign n12259 = x38 & n12258 ;
  assign n12260 = x102 & n3499 ;
  assign n12261 = x101 & n3496 ;
  assign n12262 = n12260 | n12261 ;
  assign n12263 = x100 & n3662 ;
  assign n12264 = n12262 | n12263 ;
  assign n12265 = ( ~x38 & n12258 ) | ( ~x38 & n12264 ) | ( n12258 & n12264 ) ;
  assign n12266 = x38 & ~n12264 ;
  assign n12267 = ( ~n12259 & n12265 ) | ( ~n12259 & n12266 ) | ( n12265 & n12266 ) ;
  assign n12268 = n3248 & n4020 ;
  assign n12269 = x41 & n12268 ;
  assign n12270 = x99 & n4027 ;
  assign n12271 = x98 & n4024 ;
  assign n12272 = n12270 | n12271 ;
  assign n12273 = x97 & n4223 ;
  assign n12274 = n12272 | n12273 ;
  assign n12275 = ( ~x41 & n12268 ) | ( ~x41 & n12274 ) | ( n12268 & n12274 ) ;
  assign n12276 = x41 & ~n12274 ;
  assign n12277 = ( ~n12269 & n12275 ) | ( ~n12269 & n12276 ) | ( n12275 & n12276 ) ;
  assign n12278 = n2772 & n4625 ;
  assign n12279 = x44 & n12278 ;
  assign n12280 = x96 & n4791 ;
  assign n12281 = x95 & n4621 ;
  assign n12282 = n12280 | n12281 ;
  assign n12283 = x94 & n4795 ;
  assign n12284 = n12282 | n12283 ;
  assign n12285 = ( ~x44 & n12278 ) | ( ~x44 & n12284 ) | ( n12278 & n12284 ) ;
  assign n12286 = x44 & ~n12284 ;
  assign n12287 = ( ~n12279 & n12285 ) | ( ~n12279 & n12286 ) | ( n12285 & n12286 ) ;
  assign n12288 = n2220 & n5223 ;
  assign n12289 = x47 & n12288 ;
  assign n12290 = x93 & n5230 ;
  assign n12291 = x92 & n5227 ;
  assign n12292 = n12290 | n12291 ;
  assign n12293 = x91 & n5434 ;
  assign n12294 = n12292 | n12293 ;
  assign n12295 = ( ~x47 & n12288 ) | ( ~x47 & n12294 ) | ( n12288 & n12294 ) ;
  assign n12296 = x47 & ~n12294 ;
  assign n12297 = ( ~n12289 & n12295 ) | ( ~n12289 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12298 = n1838 & n5858 ;
  assign n12299 = x50 & n12298 ;
  assign n12300 = x90 & n5865 ;
  assign n12301 = x89 & n5862 ;
  assign n12302 = n12300 | n12301 ;
  assign n12303 = x88 & n6092 ;
  assign n12304 = n12302 | n12303 ;
  assign n12305 = ( ~x50 & n12298 ) | ( ~x50 & n12304 ) | ( n12298 & n12304 ) ;
  assign n12306 = x50 & ~n12304 ;
  assign n12307 = ( ~n12299 & n12305 ) | ( ~n12299 & n12306 ) | ( n12305 & n12306 ) ;
  assign n12308 = n1494 & n6546 ;
  assign n12309 = x53 & n12308 ;
  assign n12310 = x87 & n6553 ;
  assign n12311 = x86 & n6550 ;
  assign n12312 = n12310 | n12311 ;
  assign n12313 = x85 & n6787 ;
  assign n12314 = n12312 | n12313 ;
  assign n12315 = ( ~x53 & n12308 ) | ( ~x53 & n12314 ) | ( n12308 & n12314 ) ;
  assign n12316 = x53 & ~n12314 ;
  assign n12317 = ( ~n12309 & n12315 ) | ( ~n12309 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12318 = n1190 & n7277 ;
  assign n12319 = x56 & n12318 ;
  assign n12320 = x84 & n7545 ;
  assign n12321 = x83 & n7273 ;
  assign n12322 = n12320 | n12321 ;
  assign n12323 = x82 & n7552 ;
  assign n12324 = n12322 | n12323 ;
  assign n12325 = ( ~x56 & n12318 ) | ( ~x56 & n12324 ) | ( n12318 & n12324 ) ;
  assign n12326 = x56 & ~n12324 ;
  assign n12327 = ( ~n12319 & n12325 ) | ( ~n12319 & n12326 ) | ( n12325 & n12326 ) ;
  assign n12328 = n990 & n8067 ;
  assign n12329 = x59 & n12328 ;
  assign n12330 = x81 & n8074 ;
  assign n12331 = x80 & n8071 ;
  assign n12332 = n12330 | n12331 ;
  assign n12333 = x79 & n8298 ;
  assign n12334 = n12332 | n12333 ;
  assign n12335 = ( ~x59 & n12328 ) | ( ~x59 & n12334 ) | ( n12328 & n12334 ) ;
  assign n12336 = x59 & ~n12334 ;
  assign n12337 = ( ~n12329 & n12335 ) | ( ~n12329 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12338 = n697 & n8859 ;
  assign n12339 = x62 & n12338 ;
  assign n12340 = x78 & n8866 ;
  assign n12341 = x77 & n8863 ;
  assign n12342 = n12340 | n12341 ;
  assign n12343 = x76 & n9125 ;
  assign n12344 = n12342 | n12343 ;
  assign n12345 = ( ~x62 & n12338 ) | ( ~x62 & n12344 ) | ( n12338 & n12344 ) ;
  assign n12346 = x62 & ~n12344 ;
  assign n12347 = ( ~n12339 & n12345 ) | ( ~n12339 & n12346 ) | ( n12345 & n12346 ) ;
  assign n12348 = ( x62 & x63 ) | ( x62 & x75 ) | ( x63 & x75 ) ;
  assign n12349 = ( x62 & x74 ) | ( x62 & ~n9394 ) | ( x74 & ~n9394 ) ;
  assign n12350 = ( x74 & n12348 ) | ( x74 & ~n12349 ) | ( n12348 & ~n12349 ) ;
  assign n12351 = ( ~n11871 & n12120 ) | ( ~n11871 & n12350 ) | ( n12120 & n12350 ) ;
  assign n12352 = ( n11871 & ~n12110 ) | ( n11871 & n12351 ) | ( ~n12110 & n12351 ) ;
  assign n12353 = ( n11871 & n12121 ) | ( n11871 & n12350 ) | ( n12121 & n12350 ) ;
  assign n12354 = ( n12110 & n12352 ) | ( n12110 & ~n12353 ) | ( n12352 & ~n12353 ) ;
  assign n12355 = ( n12337 & n12347 ) | ( n12337 & ~n12354 ) | ( n12347 & ~n12354 ) ;
  assign n12356 = ( n12337 & ~n12347 ) | ( n12337 & n12354 ) | ( ~n12347 & n12354 ) ;
  assign n12357 = ( ~n12337 & n12355 ) | ( ~n12337 & n12356 ) | ( n12355 & n12356 ) ;
  assign n12358 = ( n12124 & n12327 ) | ( n12124 & n12357 ) | ( n12327 & n12357 ) ;
  assign n12359 = ( n12124 & ~n12327 ) | ( n12124 & n12357 ) | ( ~n12327 & n12357 ) ;
  assign n12360 = ( n12327 & ~n12358 ) | ( n12327 & n12359 ) | ( ~n12358 & n12359 ) ;
  assign n12361 = ( n12127 & n12317 ) | ( n12127 & n12360 ) | ( n12317 & n12360 ) ;
  assign n12362 = ( n12127 & ~n12317 ) | ( n12127 & n12360 ) | ( ~n12317 & n12360 ) ;
  assign n12363 = ( n12317 & ~n12361 ) | ( n12317 & n12362 ) | ( ~n12361 & n12362 ) ;
  assign n12364 = ( n12130 & n12307 ) | ( n12130 & n12363 ) | ( n12307 & n12363 ) ;
  assign n12365 = ( n12130 & ~n12307 ) | ( n12130 & n12363 ) | ( ~n12307 & n12363 ) ;
  assign n12366 = ( n12307 & ~n12364 ) | ( n12307 & n12365 ) | ( ~n12364 & n12365 ) ;
  assign n12367 = ( n12133 & n12297 ) | ( n12133 & n12366 ) | ( n12297 & n12366 ) ;
  assign n12368 = ( n12133 & ~n12297 ) | ( n12133 & n12366 ) | ( ~n12297 & n12366 ) ;
  assign n12369 = ( n12297 & ~n12367 ) | ( n12297 & n12368 ) | ( ~n12367 & n12368 ) ;
  assign n12370 = ( n12136 & n12287 ) | ( n12136 & n12369 ) | ( n12287 & n12369 ) ;
  assign n12371 = ( n12136 & ~n12287 ) | ( n12136 & n12369 ) | ( ~n12287 & n12369 ) ;
  assign n12372 = ( n12287 & ~n12370 ) | ( n12287 & n12371 ) | ( ~n12370 & n12371 ) ;
  assign n12373 = ( n12139 & n12277 ) | ( n12139 & n12372 ) | ( n12277 & n12372 ) ;
  assign n12374 = ( n12139 & ~n12277 ) | ( n12139 & n12372 ) | ( ~n12277 & n12372 ) ;
  assign n12375 = ( n12277 & ~n12373 ) | ( n12277 & n12374 ) | ( ~n12373 & n12374 ) ;
  assign n12376 = ( n12142 & n12267 ) | ( n12142 & n12375 ) | ( n12267 & n12375 ) ;
  assign n12377 = ( n12142 & ~n12267 ) | ( n12142 & n12375 ) | ( ~n12267 & n12375 ) ;
  assign n12378 = ( n12267 & ~n12376 ) | ( n12267 & n12377 ) | ( ~n12376 & n12377 ) ;
  assign n12379 = ( n12145 & n12257 ) | ( n12145 & n12378 ) | ( n12257 & n12378 ) ;
  assign n12380 = ( n12145 & ~n12257 ) | ( n12145 & n12378 ) | ( ~n12257 & n12378 ) ;
  assign n12381 = ( n12257 & ~n12379 ) | ( n12257 & n12380 ) | ( ~n12379 & n12380 ) ;
  assign n12382 = ( n12148 & n12247 ) | ( n12148 & n12381 ) | ( n12247 & n12381 ) ;
  assign n12383 = ( n12148 & ~n12247 ) | ( n12148 & n12381 ) | ( ~n12247 & n12381 ) ;
  assign n12384 = ( n12247 & ~n12382 ) | ( n12247 & n12383 ) | ( ~n12382 & n12383 ) ;
  assign n12385 = ( n12151 & n12237 ) | ( n12151 & n12384 ) | ( n12237 & n12384 ) ;
  assign n12386 = ( n12151 & ~n12237 ) | ( n12151 & n12384 ) | ( ~n12237 & n12384 ) ;
  assign n12387 = ( n12237 & ~n12385 ) | ( n12237 & n12386 ) | ( ~n12385 & n12386 ) ;
  assign n12388 = ( n12154 & n12227 ) | ( n12154 & n12387 ) | ( n12227 & n12387 ) ;
  assign n12389 = ( n12154 & ~n12227 ) | ( n12154 & n12387 ) | ( ~n12227 & n12387 ) ;
  assign n12390 = ( n12227 & ~n12388 ) | ( n12227 & n12389 ) | ( ~n12388 & n12389 ) ;
  assign n12391 = ( n12157 & n12217 ) | ( n12157 & n12390 ) | ( n12217 & n12390 ) ;
  assign n12392 = ( n12157 & ~n12217 ) | ( n12157 & n12390 ) | ( ~n12217 & n12390 ) ;
  assign n12393 = ( n12217 & ~n12391 ) | ( n12217 & n12392 ) | ( ~n12391 & n12392 ) ;
  assign n12394 = ( n12160 & n12207 ) | ( n12160 & n12393 ) | ( n12207 & n12393 ) ;
  assign n12395 = ( n12160 & ~n12207 ) | ( n12160 & n12393 ) | ( ~n12207 & n12393 ) ;
  assign n12396 = ( n12207 & ~n12394 ) | ( n12207 & n12395 ) | ( ~n12394 & n12395 ) ;
  assign n12397 = ( n12163 & n12197 ) | ( n12163 & n12396 ) | ( n12197 & n12396 ) ;
  assign n12398 = ( ~n12163 & n12197 ) | ( ~n12163 & n12396 ) | ( n12197 & n12396 ) ;
  assign n12399 = ( n12163 & ~n12397 ) | ( n12163 & n12398 ) | ( ~n12397 & n12398 ) ;
  assign n12400 = ( n12166 & n12187 ) | ( n12166 & n12399 ) | ( n12187 & n12399 ) ;
  assign n12401 = ( n12166 & ~n12187 ) | ( n12166 & n12399 ) | ( ~n12187 & n12399 ) ;
  assign n12402 = ( n12187 & ~n12400 ) | ( n12187 & n12401 ) | ( ~n12400 & n12401 ) ;
  assign n12403 = x127 & n536 ;
  assign n12404 = n449 | n12403 ;
  assign n12405 = ( n9865 & n12403 ) | ( n9865 & n12404 ) | ( n12403 & n12404 ) ;
  assign n12406 = x11 & ~n12405 ;
  assign n12407 = ~x11 & n12405 ;
  assign n12408 = n12406 | n12407 ;
  assign n12409 = ( n12169 & n12402 ) | ( n12169 & n12408 ) | ( n12402 & n12408 ) ;
  assign n12410 = ( n12169 & ~n12402 ) | ( n12169 & n12408 ) | ( ~n12402 & n12408 ) ;
  assign n12411 = ( n12402 & ~n12409 ) | ( n12402 & n12410 ) | ( ~n12409 & n12410 ) ;
  assign n12412 = ( n12172 & ~n12176 ) | ( n12172 & n12411 ) | ( ~n12176 & n12411 ) ;
  assign n12413 = ( n12172 & n12176 ) | ( n12172 & n12411 ) | ( n12176 & n12411 ) ;
  assign n12414 = ( n12176 & n12412 ) | ( n12176 & ~n12413 ) | ( n12412 & ~n12413 ) ;
  assign n12415 = n649 & n9576 ;
  assign n12416 = x14 & n12415 ;
  assign n12417 = x127 & n656 ;
  assign n12418 = x126 & n653 ;
  assign n12419 = n12417 | n12418 ;
  assign n12420 = x125 & n744 ;
  assign n12421 = n12419 | n12420 ;
  assign n12422 = ( ~x14 & n12415 ) | ( ~x14 & n12421 ) | ( n12415 & n12421 ) ;
  assign n12423 = x14 & ~n12421 ;
  assign n12424 = ( ~n12416 & n12422 ) | ( ~n12416 & n12423 ) | ( n12422 & n12423 ) ;
  assign n12425 = n874 & n8729 ;
  assign n12426 = x17 & n12425 ;
  assign n12427 = x124 & n881 ;
  assign n12428 = x123 & n878 ;
  assign n12429 = n12427 | n12428 ;
  assign n12430 = x122 & n959 ;
  assign n12431 = n12429 | n12430 ;
  assign n12432 = ( ~x17 & n12425 ) | ( ~x17 & n12431 ) | ( n12425 & n12431 ) ;
  assign n12433 = x17 & ~n12431 ;
  assign n12434 = ( ~n12426 & n12432 ) | ( ~n12426 & n12433 ) | ( n12432 & n12433 ) ;
  assign n12435 = n1146 & n7696 ;
  assign n12436 = x20 & n12435 ;
  assign n12437 = x121 & n1153 ;
  assign n12438 = x120 & n1150 ;
  assign n12439 = n12437 | n12438 ;
  assign n12440 = x119 & n1217 ;
  assign n12441 = n12439 | n12440 ;
  assign n12442 = ( ~x20 & n12435 ) | ( ~x20 & n12441 ) | ( n12435 & n12441 ) ;
  assign n12443 = x20 & ~n12441 ;
  assign n12444 = ( ~n12436 & n12442 ) | ( ~n12436 & n12443 ) | ( n12442 & n12443 ) ;
  assign n12445 = n1427 & n6940 ;
  assign n12446 = x23 & n12445 ;
  assign n12447 = x118 & n1434 ;
  assign n12448 = x117 & n1431 ;
  assign n12449 = n12447 | n12448 ;
  assign n12450 = x116 & n1531 ;
  assign n12451 = n12449 | n12450 ;
  assign n12452 = ( ~x23 & n12445 ) | ( ~x23 & n12451 ) | ( n12445 & n12451 ) ;
  assign n12453 = x23 & ~n12451 ;
  assign n12454 = ( ~n12446 & n12452 ) | ( ~n12446 & n12453 ) | ( n12452 & n12453 ) ;
  assign n12455 = n1755 & n6446 ;
  assign n12456 = x26 & n12455 ;
  assign n12457 = x115 & n1762 ;
  assign n12458 = x114 & n1759 ;
  assign n12459 = n12457 | n12458 ;
  assign n12460 = x113 & n1895 ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = ( ~x26 & n12455 ) | ( ~x26 & n12461 ) | ( n12455 & n12461 ) ;
  assign n12463 = x26 & ~n12461 ;
  assign n12464 = ( ~n12456 & n12462 ) | ( ~n12456 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = n2137 & n5558 ;
  assign n12466 = x29 & n12465 ;
  assign n12467 = x112 & n2144 ;
  assign n12468 = x111 & n2141 ;
  assign n12469 = n12467 | n12468 ;
  assign n12470 = x110 & n2267 ;
  assign n12471 = n12469 | n12470 ;
  assign n12472 = ( ~x29 & n12465 ) | ( ~x29 & n12471 ) | ( n12465 & n12471 ) ;
  assign n12473 = x29 & ~n12471 ;
  assign n12474 = ( ~n12466 & n12472 ) | ( ~n12466 & n12473 ) | ( n12472 & n12473 ) ;
  assign n12475 = n2545 & n4930 ;
  assign n12476 = x32 & n12475 ;
  assign n12477 = x109 & n2552 ;
  assign n12478 = x108 & n2549 ;
  assign n12479 = n12477 | n12478 ;
  assign n12480 = x107 & n2696 ;
  assign n12481 = n12479 | n12480 ;
  assign n12482 = ( ~x32 & n12475 ) | ( ~x32 & n12481 ) | ( n12475 & n12481 ) ;
  assign n12483 = x32 & ~n12481 ;
  assign n12484 = ( ~n12476 & n12482 ) | ( ~n12476 & n12483 ) | ( n12482 & n12483 ) ;
  assign n12485 = n2982 & n4331 ;
  assign n12486 = x35 & n12485 ;
  assign n12487 = x106 & n2989 ;
  assign n12488 = x105 & n2986 ;
  assign n12489 = n12487 | n12488 ;
  assign n12490 = x104 & n3159 ;
  assign n12491 = n12489 | n12490 ;
  assign n12492 = ( ~x35 & n12485 ) | ( ~x35 & n12491 ) | ( n12485 & n12491 ) ;
  assign n12493 = x35 & ~n12491 ;
  assign n12494 = ( ~n12486 & n12492 ) | ( ~n12486 & n12493 ) | ( n12492 & n12493 ) ;
  assign n12495 = n3492 & n3941 ;
  assign n12496 = x38 & n12495 ;
  assign n12497 = x102 & n3496 ;
  assign n12498 = x101 & n3662 ;
  assign n12499 = n12497 | n12498 ;
  assign n12500 = x103 & n3499 ;
  assign n12501 = n12499 | n12500 ;
  assign n12502 = ( ~x38 & n12495 ) | ( ~x38 & n12501 ) | ( n12495 & n12501 ) ;
  assign n12503 = x38 & ~n12501 ;
  assign n12504 = ( ~n12496 & n12502 ) | ( ~n12496 & n12503 ) | ( n12502 & n12503 ) ;
  assign n12505 = n3264 & n4020 ;
  assign n12506 = x41 & n12505 ;
  assign n12507 = x100 & n4027 ;
  assign n12508 = x99 & n4024 ;
  assign n12509 = n12507 | n12508 ;
  assign n12510 = x98 & n4223 ;
  assign n12511 = n12509 | n12510 ;
  assign n12512 = ( ~x41 & n12505 ) | ( ~x41 & n12511 ) | ( n12505 & n12511 ) ;
  assign n12513 = x41 & ~n12511 ;
  assign n12514 = ( ~n12506 & n12512 ) | ( ~n12506 & n12513 ) | ( n12512 & n12513 ) ;
  assign n12515 = n2788 & n4625 ;
  assign n12516 = x44 & n12515 ;
  assign n12517 = x97 & n4791 ;
  assign n12518 = x96 & n4621 ;
  assign n12519 = n12517 | n12518 ;
  assign n12520 = x95 & n4795 ;
  assign n12521 = n12519 | n12520 ;
  assign n12522 = ( ~x44 & n12515 ) | ( ~x44 & n12521 ) | ( n12515 & n12521 ) ;
  assign n12523 = x44 & ~n12521 ;
  assign n12524 = ( ~n12516 & n12522 ) | ( ~n12516 & n12523 ) | ( n12522 & n12523 ) ;
  assign n12525 = n2476 & n5223 ;
  assign n12526 = x47 & n12525 ;
  assign n12527 = x94 & n5230 ;
  assign n12528 = x93 & n5227 ;
  assign n12529 = n12527 | n12528 ;
  assign n12530 = x92 & n5434 ;
  assign n12531 = n12529 | n12530 ;
  assign n12532 = ( ~x47 & n12525 ) | ( ~x47 & n12531 ) | ( n12525 & n12531 ) ;
  assign n12533 = x47 & ~n12531 ;
  assign n12534 = ( ~n12526 & n12532 ) | ( ~n12526 & n12533 ) | ( n12532 & n12533 ) ;
  assign n12535 = n1959 & n5858 ;
  assign n12536 = x50 & n12535 ;
  assign n12537 = x91 & n5865 ;
  assign n12538 = x90 & n5862 ;
  assign n12539 = n12537 | n12538 ;
  assign n12540 = x89 & n6092 ;
  assign n12541 = n12539 | n12540 ;
  assign n12542 = ( ~x50 & n12535 ) | ( ~x50 & n12541 ) | ( n12535 & n12541 ) ;
  assign n12543 = x50 & ~n12541 ;
  assign n12544 = ( ~n12536 & n12542 ) | ( ~n12536 & n12543 ) | ( n12542 & n12543 ) ;
  assign n12545 = n1602 & n6546 ;
  assign n12546 = x53 & n12545 ;
  assign n12547 = x88 & n6553 ;
  assign n12548 = x87 & n6550 ;
  assign n12549 = n12547 | n12548 ;
  assign n12550 = x86 & n6787 ;
  assign n12551 = n12549 | n12550 ;
  assign n12552 = ( ~x53 & n12545 ) | ( ~x53 & n12551 ) | ( n12545 & n12551 ) ;
  assign n12553 = x53 & ~n12551 ;
  assign n12554 = ( ~n12546 & n12552 ) | ( ~n12546 & n12553 ) | ( n12552 & n12553 ) ;
  assign n12555 = n1368 & n7277 ;
  assign n12556 = x56 & n12555 ;
  assign n12557 = x85 & n7545 ;
  assign n12558 = x84 & n7273 ;
  assign n12559 = n12557 | n12558 ;
  assign n12560 = x83 & n7552 ;
  assign n12561 = n12559 | n12560 ;
  assign n12562 = ( ~x56 & n12555 ) | ( ~x56 & n12561 ) | ( n12555 & n12561 ) ;
  assign n12563 = x56 & ~n12561 ;
  assign n12564 = ( ~n12556 & n12562 ) | ( ~n12556 & n12563 ) | ( n12562 & n12563 ) ;
  assign n12565 = n1006 & n8067 ;
  assign n12566 = x59 & n12565 ;
  assign n12567 = x82 & n8074 ;
  assign n12568 = x81 & n8071 ;
  assign n12569 = n12567 | n12568 ;
  assign n12570 = x80 & n8298 ;
  assign n12571 = n12569 | n12570 ;
  assign n12572 = ( ~x59 & n12565 ) | ( ~x59 & n12571 ) | ( n12565 & n12571 ) ;
  assign n12573 = x59 & ~n12571 ;
  assign n12574 = ( ~n12566 & n12572 ) | ( ~n12566 & n12573 ) | ( n12572 & n12573 ) ;
  assign n12575 = n823 & n8859 ;
  assign n12576 = x62 & n12575 ;
  assign n12577 = x79 & n8866 ;
  assign n12578 = x78 & n8863 ;
  assign n12579 = n12577 | n12578 ;
  assign n12580 = x77 & n9125 ;
  assign n12581 = n12579 | n12580 ;
  assign n12582 = ( ~x62 & n12575 ) | ( ~x62 & n12581 ) | ( n12575 & n12581 ) ;
  assign n12583 = x62 & ~n12581 ;
  assign n12584 = ( ~n12576 & n12582 ) | ( ~n12576 & n12583 ) | ( n12582 & n12583 ) ;
  assign n12585 = ( x62 & x63 ) | ( x62 & x76 ) | ( x63 & x76 ) ;
  assign n12586 = ( x62 & x75 ) | ( x62 & ~n9394 ) | ( x75 & ~n9394 ) ;
  assign n12587 = ( x75 & n12585 ) | ( x75 & ~n12586 ) | ( n12585 & ~n12586 ) ;
  assign n12588 = ( x11 & n12110 ) | ( x11 & n12587 ) | ( n12110 & n12587 ) ;
  assign n12589 = ( ~x11 & n12110 ) | ( ~x11 & n12587 ) | ( n12110 & n12587 ) ;
  assign n12590 = ( x11 & ~n12588 ) | ( x11 & n12589 ) | ( ~n12588 & n12589 ) ;
  assign n12591 = ( n12352 & n12584 ) | ( n12352 & ~n12590 ) | ( n12584 & ~n12590 ) ;
  assign n12592 = ( n12352 & ~n12584 ) | ( n12352 & n12590 ) | ( ~n12584 & n12590 ) ;
  assign n12593 = ( ~n12352 & n12591 ) | ( ~n12352 & n12592 ) | ( n12591 & n12592 ) ;
  assign n12594 = ( n12355 & n12574 ) | ( n12355 & ~n12593 ) | ( n12574 & ~n12593 ) ;
  assign n12595 = ( n12355 & ~n12574 ) | ( n12355 & n12593 ) | ( ~n12574 & n12593 ) ;
  assign n12596 = ( ~n12355 & n12594 ) | ( ~n12355 & n12595 ) | ( n12594 & n12595 ) ;
  assign n12597 = ( n12359 & ~n12564 ) | ( n12359 & n12596 ) | ( ~n12564 & n12596 ) ;
  assign n12598 = ( n12359 & n12564 ) | ( n12359 & ~n12596 ) | ( n12564 & ~n12596 ) ;
  assign n12599 = ( ~n12359 & n12597 ) | ( ~n12359 & n12598 ) | ( n12597 & n12598 ) ;
  assign n12600 = ( n12361 & n12554 ) | ( n12361 & n12599 ) | ( n12554 & n12599 ) ;
  assign n12601 = ( ~n12361 & n12554 ) | ( ~n12361 & n12599 ) | ( n12554 & n12599 ) ;
  assign n12602 = ( n12361 & ~n12600 ) | ( n12361 & n12601 ) | ( ~n12600 & n12601 ) ;
  assign n12603 = ( n12364 & n12544 ) | ( n12364 & n12602 ) | ( n12544 & n12602 ) ;
  assign n12604 = ( ~n12364 & n12544 ) | ( ~n12364 & n12602 ) | ( n12544 & n12602 ) ;
  assign n12605 = ( n12364 & ~n12603 ) | ( n12364 & n12604 ) | ( ~n12603 & n12604 ) ;
  assign n12606 = ( n12367 & n12534 ) | ( n12367 & n12605 ) | ( n12534 & n12605 ) ;
  assign n12607 = ( n12367 & ~n12534 ) | ( n12367 & n12605 ) | ( ~n12534 & n12605 ) ;
  assign n12608 = ( n12534 & ~n12606 ) | ( n12534 & n12607 ) | ( ~n12606 & n12607 ) ;
  assign n12609 = ( n12370 & n12524 ) | ( n12370 & n12608 ) | ( n12524 & n12608 ) ;
  assign n12610 = ( ~n12370 & n12524 ) | ( ~n12370 & n12608 ) | ( n12524 & n12608 ) ;
  assign n12611 = ( n12370 & ~n12609 ) | ( n12370 & n12610 ) | ( ~n12609 & n12610 ) ;
  assign n12612 = ( n12373 & n12514 ) | ( n12373 & n12611 ) | ( n12514 & n12611 ) ;
  assign n12613 = ( ~n12373 & n12514 ) | ( ~n12373 & n12611 ) | ( n12514 & n12611 ) ;
  assign n12614 = ( n12373 & ~n12612 ) | ( n12373 & n12613 ) | ( ~n12612 & n12613 ) ;
  assign n12615 = ( n12376 & n12504 ) | ( n12376 & n12614 ) | ( n12504 & n12614 ) ;
  assign n12616 = ( n12376 & ~n12504 ) | ( n12376 & n12614 ) | ( ~n12504 & n12614 ) ;
  assign n12617 = ( n12504 & ~n12615 ) | ( n12504 & n12616 ) | ( ~n12615 & n12616 ) ;
  assign n12618 = ( n12379 & n12494 ) | ( n12379 & n12617 ) | ( n12494 & n12617 ) ;
  assign n12619 = ( ~n12379 & n12494 ) | ( ~n12379 & n12617 ) | ( n12494 & n12617 ) ;
  assign n12620 = ( n12379 & ~n12618 ) | ( n12379 & n12619 ) | ( ~n12618 & n12619 ) ;
  assign n12621 = ( n12382 & n12484 ) | ( n12382 & n12620 ) | ( n12484 & n12620 ) ;
  assign n12622 = ( ~n12382 & n12484 ) | ( ~n12382 & n12620 ) | ( n12484 & n12620 ) ;
  assign n12623 = ( n12382 & ~n12621 ) | ( n12382 & n12622 ) | ( ~n12621 & n12622 ) ;
  assign n12624 = ( n12385 & n12474 ) | ( n12385 & n12623 ) | ( n12474 & n12623 ) ;
  assign n12625 = ( ~n12385 & n12474 ) | ( ~n12385 & n12623 ) | ( n12474 & n12623 ) ;
  assign n12626 = ( n12385 & ~n12624 ) | ( n12385 & n12625 ) | ( ~n12624 & n12625 ) ;
  assign n12627 = ( n12388 & n12464 ) | ( n12388 & n12626 ) | ( n12464 & n12626 ) ;
  assign n12628 = ( ~n12388 & n12464 ) | ( ~n12388 & n12626 ) | ( n12464 & n12626 ) ;
  assign n12629 = ( n12388 & ~n12627 ) | ( n12388 & n12628 ) | ( ~n12627 & n12628 ) ;
  assign n12630 = ( n12391 & n12454 ) | ( n12391 & n12629 ) | ( n12454 & n12629 ) ;
  assign n12631 = ( ~n12391 & n12454 ) | ( ~n12391 & n12629 ) | ( n12454 & n12629 ) ;
  assign n12632 = ( n12391 & ~n12630 ) | ( n12391 & n12631 ) | ( ~n12630 & n12631 ) ;
  assign n12633 = ( n12394 & n12444 ) | ( n12394 & n12632 ) | ( n12444 & n12632 ) ;
  assign n12634 = ( ~n12394 & n12444 ) | ( ~n12394 & n12632 ) | ( n12444 & n12632 ) ;
  assign n12635 = ( n12394 & ~n12633 ) | ( n12394 & n12634 ) | ( ~n12633 & n12634 ) ;
  assign n12636 = ( n12397 & n12434 ) | ( n12397 & n12635 ) | ( n12434 & n12635 ) ;
  assign n12637 = ( ~n12397 & n12434 ) | ( ~n12397 & n12635 ) | ( n12434 & n12635 ) ;
  assign n12638 = ( n12397 & ~n12636 ) | ( n12397 & n12637 ) | ( ~n12636 & n12637 ) ;
  assign n12639 = ( n12400 & n12424 ) | ( n12400 & n12638 ) | ( n12424 & n12638 ) ;
  assign n12640 = ( ~n12400 & n12424 ) | ( ~n12400 & n12638 ) | ( n12424 & n12638 ) ;
  assign n12641 = ( n12400 & ~n12639 ) | ( n12400 & n12640 ) | ( ~n12639 & n12640 ) ;
  assign n12642 = ( n12409 & n12413 ) | ( n12409 & n12641 ) | ( n12413 & n12641 ) ;
  assign n12643 = ( n12409 & ~n12413 ) | ( n12409 & n12641 ) | ( ~n12413 & n12641 ) ;
  assign n12644 = ( n12413 & ~n12642 ) | ( n12413 & n12643 ) | ( ~n12642 & n12643 ) ;
  assign n12645 = x126 & n744 ;
  assign n12646 = x14 & n12645 ;
  assign n12647 = x127 & n653 ;
  assign n12648 = n649 | n12647 ;
  assign n12649 = ( n9867 & n12647 ) | ( n9867 & n12648 ) | ( n12647 & n12648 ) ;
  assign n12650 = ( ~x14 & n12645 ) | ( ~x14 & n12649 ) | ( n12645 & n12649 ) ;
  assign n12651 = x14 & ~n12649 ;
  assign n12652 = ( ~n12646 & n12650 ) | ( ~n12646 & n12651 ) | ( n12650 & n12651 ) ;
  assign n12653 = n874 & n9009 ;
  assign n12654 = x17 & n12653 ;
  assign n12655 = x125 & n881 ;
  assign n12656 = x124 & n878 ;
  assign n12657 = n12655 | n12656 ;
  assign n12658 = x123 & n959 ;
  assign n12659 = n12657 | n12658 ;
  assign n12660 = ( ~x17 & n12653 ) | ( ~x17 & n12659 ) | ( n12653 & n12659 ) ;
  assign n12661 = x17 & ~n12659 ;
  assign n12662 = ( ~n12654 & n12660 ) | ( ~n12654 & n12661 ) | ( n12660 & n12661 ) ;
  assign n12663 = n1146 & n8207 ;
  assign n12664 = x20 & n12663 ;
  assign n12665 = x122 & n1153 ;
  assign n12666 = x121 & n1150 ;
  assign n12667 = n12665 | n12666 ;
  assign n12668 = x120 & n1217 ;
  assign n12669 = n12667 | n12668 ;
  assign n12670 = ( ~x20 & n12663 ) | ( ~x20 & n12669 ) | ( n12663 & n12669 ) ;
  assign n12671 = x20 & ~n12669 ;
  assign n12672 = ( ~n12664 & n12670 ) | ( ~n12664 & n12671 ) | ( n12670 & n12671 ) ;
  assign n12673 = n1427 & n7181 ;
  assign n12674 = x23 & n12673 ;
  assign n12675 = x119 & n1434 ;
  assign n12676 = x118 & n1431 ;
  assign n12677 = n12675 | n12676 ;
  assign n12678 = x117 & n1531 ;
  assign n12679 = n12677 | n12678 ;
  assign n12680 = ( ~x23 & n12673 ) | ( ~x23 & n12679 ) | ( n12673 & n12679 ) ;
  assign n12681 = x23 & ~n12679 ;
  assign n12682 = ( ~n12674 & n12680 ) | ( ~n12674 & n12681 ) | ( n12680 & n12681 ) ;
  assign n12683 = n1755 & n6462 ;
  assign n12684 = x26 & n12683 ;
  assign n12685 = x116 & n1762 ;
  assign n12686 = x115 & n1759 ;
  assign n12687 = n12685 | n12686 ;
  assign n12688 = x114 & n1895 ;
  assign n12689 = n12687 | n12688 ;
  assign n12690 = ( ~x26 & n12683 ) | ( ~x26 & n12689 ) | ( n12683 & n12689 ) ;
  assign n12691 = x26 & ~n12689 ;
  assign n12692 = ( ~n12684 & n12690 ) | ( ~n12684 & n12691 ) | ( n12690 & n12691 ) ;
  assign n12693 = n2137 & n5774 ;
  assign n12694 = x29 & n12693 ;
  assign n12695 = x113 & n2144 ;
  assign n12696 = x112 & n2141 ;
  assign n12697 = n12695 | n12696 ;
  assign n12698 = x111 & n2267 ;
  assign n12699 = n12697 | n12698 ;
  assign n12700 = ( ~x29 & n12693 ) | ( ~x29 & n12699 ) | ( n12693 & n12699 ) ;
  assign n12701 = x29 & ~n12699 ;
  assign n12702 = ( ~n12694 & n12700 ) | ( ~n12694 & n12701 ) | ( n12700 & n12701 ) ;
  assign n12703 = n2545 & n5331 ;
  assign n12704 = x32 & n12703 ;
  assign n12705 = x110 & n2552 ;
  assign n12706 = x109 & n2549 ;
  assign n12707 = n12705 | n12706 ;
  assign n12708 = x108 & n2696 ;
  assign n12709 = n12707 | n12708 ;
  assign n12710 = ( ~x32 & n12703 ) | ( ~x32 & n12709 ) | ( n12703 & n12709 ) ;
  assign n12711 = x32 & ~n12709 ;
  assign n12712 = ( ~n12704 & n12710 ) | ( ~n12704 & n12711 ) | ( n12710 & n12711 ) ;
  assign n12713 = n2982 & n4523 ;
  assign n12714 = x35 & n12713 ;
  assign n12715 = x107 & n2989 ;
  assign n12716 = x106 & n2986 ;
  assign n12717 = n12715 | n12716 ;
  assign n12718 = x105 & n3159 ;
  assign n12719 = n12717 | n12718 ;
  assign n12720 = ( ~x35 & n12713 ) | ( ~x35 & n12719 ) | ( n12713 & n12719 ) ;
  assign n12721 = x35 & ~n12719 ;
  assign n12722 = ( ~n12714 & n12720 ) | ( ~n12714 & n12721 ) | ( n12720 & n12721 ) ;
  assign n12723 = n3492 & n3957 ;
  assign n12724 = x38 & n12723 ;
  assign n12725 = x104 & n3499 ;
  assign n12726 = x103 & n3496 ;
  assign n12727 = n12725 | n12726 ;
  assign n12728 = x102 & n3662 ;
  assign n12729 = n12727 | n12728 ;
  assign n12730 = ( ~x38 & n12723 ) | ( ~x38 & n12729 ) | ( n12723 & n12729 ) ;
  assign n12731 = x38 & ~n12729 ;
  assign n12732 = ( ~n12724 & n12730 ) | ( ~n12724 & n12731 ) | ( n12730 & n12731 ) ;
  assign n12733 = n3591 & n4020 ;
  assign n12734 = x41 & n12733 ;
  assign n12735 = x101 & n4027 ;
  assign n12736 = x100 & n4024 ;
  assign n12737 = n12735 | n12736 ;
  assign n12738 = x99 & n4223 ;
  assign n12739 = n12737 | n12738 ;
  assign n12740 = ( ~x41 & n12733 ) | ( ~x41 & n12739 ) | ( n12733 & n12739 ) ;
  assign n12741 = x41 & ~n12739 ;
  assign n12742 = ( ~n12734 & n12740 ) | ( ~n12734 & n12741 ) | ( n12740 & n12741 ) ;
  assign n12743 = n2939 & n4625 ;
  assign n12744 = x44 & n12743 ;
  assign n12745 = x98 & n4791 ;
  assign n12746 = x97 & n4621 ;
  assign n12747 = n12745 | n12746 ;
  assign n12748 = x96 & n4795 ;
  assign n12749 = n12747 | n12748 ;
  assign n12750 = ( ~x44 & n12743 ) | ( ~x44 & n12749 ) | ( n12743 & n12749 ) ;
  assign n12751 = x44 & ~n12749 ;
  assign n12752 = ( ~n12744 & n12750 ) | ( ~n12744 & n12751 ) | ( n12750 & n12751 ) ;
  assign n12753 = n2492 & n5223 ;
  assign n12754 = x47 & n12753 ;
  assign n12755 = x95 & n5230 ;
  assign n12756 = x94 & n5227 ;
  assign n12757 = n12755 | n12756 ;
  assign n12758 = x93 & n5434 ;
  assign n12759 = n12757 | n12758 ;
  assign n12760 = ( ~x47 & n12753 ) | ( ~x47 & n12759 ) | ( n12753 & n12759 ) ;
  assign n12761 = x47 & ~n12759 ;
  assign n12762 = ( ~n12754 & n12760 ) | ( ~n12754 & n12761 ) | ( n12760 & n12761 ) ;
  assign n12763 = n2083 & n5858 ;
  assign n12764 = x50 & n12763 ;
  assign n12765 = x92 & n5865 ;
  assign n12766 = x91 & n5862 ;
  assign n12767 = n12765 | n12766 ;
  assign n12768 = x90 & n6092 ;
  assign n12769 = n12767 | n12768 ;
  assign n12770 = ( ~x50 & n12763 ) | ( ~x50 & n12769 ) | ( n12763 & n12769 ) ;
  assign n12771 = x50 & ~n12769 ;
  assign n12772 = ( ~n12764 & n12770 ) | ( ~n12764 & n12771 ) | ( n12770 & n12771 ) ;
  assign n12773 = n1822 & n6546 ;
  assign n12774 = x53 & n12773 ;
  assign n12775 = x89 & n6553 ;
  assign n12776 = x88 & n6550 ;
  assign n12777 = n12775 | n12776 ;
  assign n12778 = x87 & n6787 ;
  assign n12779 = n12777 | n12778 ;
  assign n12780 = ( ~x53 & n12773 ) | ( ~x53 & n12779 ) | ( n12773 & n12779 ) ;
  assign n12781 = x53 & ~n12779 ;
  assign n12782 = ( ~n12774 & n12780 ) | ( ~n12774 & n12781 ) | ( n12780 & n12781 ) ;
  assign n12783 = n1384 & n7277 ;
  assign n12784 = x56 & n12783 ;
  assign n12785 = x86 & n7545 ;
  assign n12786 = x85 & n7273 ;
  assign n12787 = n12785 | n12786 ;
  assign n12788 = x84 & n7552 ;
  assign n12789 = n12787 | n12788 ;
  assign n12790 = ( ~x56 & n12783 ) | ( ~x56 & n12789 ) | ( n12783 & n12789 ) ;
  assign n12791 = x56 & ~n12789 ;
  assign n12792 = ( ~n12784 & n12790 ) | ( ~n12784 & n12791 ) | ( n12790 & n12791 ) ;
  assign n12793 = n1093 & n8067 ;
  assign n12794 = x59 & n12793 ;
  assign n12795 = x83 & n8074 ;
  assign n12796 = x82 & n8071 ;
  assign n12797 = n12795 | n12796 ;
  assign n12798 = x81 & n8298 ;
  assign n12799 = n12797 | n12798 ;
  assign n12800 = ( ~x59 & n12793 ) | ( ~x59 & n12799 ) | ( n12793 & n12799 ) ;
  assign n12801 = x59 & ~n12799 ;
  assign n12802 = ( ~n12794 & n12800 ) | ( ~n12794 & n12801 ) | ( n12800 & n12801 ) ;
  assign n12803 = n840 & n8859 ;
  assign n12804 = x62 & n12803 ;
  assign n12805 = x80 & n8866 ;
  assign n12806 = x79 & n8863 ;
  assign n12807 = n12805 | n12806 ;
  assign n12808 = x78 & n9125 ;
  assign n12809 = n12807 | n12808 ;
  assign n12810 = ( ~x62 & n12803 ) | ( ~x62 & n12809 ) | ( n12803 & n12809 ) ;
  assign n12811 = x62 & ~n12809 ;
  assign n12812 = ( ~n12804 & n12810 ) | ( ~n12804 & n12811 ) | ( n12810 & n12811 ) ;
  assign n12813 = ( x62 & x63 ) | ( x62 & x77 ) | ( x63 & x77 ) ;
  assign n12814 = ( x62 & x76 ) | ( x62 & ~n9394 ) | ( x76 & ~n9394 ) ;
  assign n12815 = ( x76 & n12813 ) | ( x76 & ~n12814 ) | ( n12813 & ~n12814 ) ;
  assign n12816 = ( n12589 & n12812 ) | ( n12589 & ~n12815 ) | ( n12812 & ~n12815 ) ;
  assign n12817 = ( ~n12589 & n12812 ) | ( ~n12589 & n12815 ) | ( n12812 & n12815 ) ;
  assign n12818 = ( ~n12812 & n12816 ) | ( ~n12812 & n12817 ) | ( n12816 & n12817 ) ;
  assign n12819 = ( n12591 & n12802 ) | ( n12591 & ~n12818 ) | ( n12802 & ~n12818 ) ;
  assign n12820 = ( ~n12591 & n12802 ) | ( ~n12591 & n12818 ) | ( n12802 & n12818 ) ;
  assign n12821 = ( ~n12802 & n12819 ) | ( ~n12802 & n12820 ) | ( n12819 & n12820 ) ;
  assign n12822 = ( n12594 & n12792 ) | ( n12594 & ~n12821 ) | ( n12792 & ~n12821 ) ;
  assign n12823 = ( ~n12594 & n12792 ) | ( ~n12594 & n12821 ) | ( n12792 & n12821 ) ;
  assign n12824 = ( ~n12792 & n12822 ) | ( ~n12792 & n12823 ) | ( n12822 & n12823 ) ;
  assign n12825 = ( n12597 & n12782 ) | ( n12597 & n12824 ) | ( n12782 & n12824 ) ;
  assign n12826 = ( n12597 & ~n12782 ) | ( n12597 & n12824 ) | ( ~n12782 & n12824 ) ;
  assign n12827 = ( n12782 & ~n12825 ) | ( n12782 & n12826 ) | ( ~n12825 & n12826 ) ;
  assign n12828 = ( n12600 & ~n12772 ) | ( n12600 & n12827 ) | ( ~n12772 & n12827 ) ;
  assign n12829 = ( n12600 & n12772 ) | ( n12600 & n12827 ) | ( n12772 & n12827 ) ;
  assign n12830 = ( n12772 & n12828 ) | ( n12772 & ~n12829 ) | ( n12828 & ~n12829 ) ;
  assign n12831 = ( n12603 & ~n12762 ) | ( n12603 & n12830 ) | ( ~n12762 & n12830 ) ;
  assign n12832 = ( n12603 & n12762 ) | ( n12603 & n12830 ) | ( n12762 & n12830 ) ;
  assign n12833 = ( n12762 & n12831 ) | ( n12762 & ~n12832 ) | ( n12831 & ~n12832 ) ;
  assign n12834 = ( n12606 & ~n12752 ) | ( n12606 & n12833 ) | ( ~n12752 & n12833 ) ;
  assign n12835 = ( n12606 & n12752 ) | ( n12606 & n12833 ) | ( n12752 & n12833 ) ;
  assign n12836 = ( n12752 & n12834 ) | ( n12752 & ~n12835 ) | ( n12834 & ~n12835 ) ;
  assign n12837 = ( n12609 & n12742 ) | ( n12609 & n12836 ) | ( n12742 & n12836 ) ;
  assign n12838 = ( n12609 & ~n12742 ) | ( n12609 & n12836 ) | ( ~n12742 & n12836 ) ;
  assign n12839 = ( n12742 & ~n12837 ) | ( n12742 & n12838 ) | ( ~n12837 & n12838 ) ;
  assign n12840 = ( n12612 & n12732 ) | ( n12612 & n12839 ) | ( n12732 & n12839 ) ;
  assign n12841 = ( n12612 & ~n12732 ) | ( n12612 & n12839 ) | ( ~n12732 & n12839 ) ;
  assign n12842 = ( n12732 & ~n12840 ) | ( n12732 & n12841 ) | ( ~n12840 & n12841 ) ;
  assign n12843 = ( n12615 & n12722 ) | ( n12615 & n12842 ) | ( n12722 & n12842 ) ;
  assign n12844 = ( n12615 & ~n12722 ) | ( n12615 & n12842 ) | ( ~n12722 & n12842 ) ;
  assign n12845 = ( n12722 & ~n12843 ) | ( n12722 & n12844 ) | ( ~n12843 & n12844 ) ;
  assign n12846 = ( n12618 & ~n12712 ) | ( n12618 & n12845 ) | ( ~n12712 & n12845 ) ;
  assign n12847 = ( n12618 & n12712 ) | ( n12618 & n12845 ) | ( n12712 & n12845 ) ;
  assign n12848 = ( n12712 & n12846 ) | ( n12712 & ~n12847 ) | ( n12846 & ~n12847 ) ;
  assign n12849 = ( n12621 & n12702 ) | ( n12621 & n12848 ) | ( n12702 & n12848 ) ;
  assign n12850 = ( n12621 & ~n12702 ) | ( n12621 & n12848 ) | ( ~n12702 & n12848 ) ;
  assign n12851 = ( n12702 & ~n12849 ) | ( n12702 & n12850 ) | ( ~n12849 & n12850 ) ;
  assign n12852 = ( n12624 & n12692 ) | ( n12624 & n12851 ) | ( n12692 & n12851 ) ;
  assign n12853 = ( n12624 & ~n12692 ) | ( n12624 & n12851 ) | ( ~n12692 & n12851 ) ;
  assign n12854 = ( n12692 & ~n12852 ) | ( n12692 & n12853 ) | ( ~n12852 & n12853 ) ;
  assign n12855 = ( n12627 & n12682 ) | ( n12627 & n12854 ) | ( n12682 & n12854 ) ;
  assign n12856 = ( n12627 & ~n12682 ) | ( n12627 & n12854 ) | ( ~n12682 & n12854 ) ;
  assign n12857 = ( n12682 & ~n12855 ) | ( n12682 & n12856 ) | ( ~n12855 & n12856 ) ;
  assign n12858 = ( n12630 & n12672 ) | ( n12630 & n12857 ) | ( n12672 & n12857 ) ;
  assign n12859 = ( n12630 & ~n12672 ) | ( n12630 & n12857 ) | ( ~n12672 & n12857 ) ;
  assign n12860 = ( n12672 & ~n12858 ) | ( n12672 & n12859 ) | ( ~n12858 & n12859 ) ;
  assign n12861 = ( n12633 & n12662 ) | ( n12633 & n12860 ) | ( n12662 & n12860 ) ;
  assign n12862 = ( n12633 & ~n12662 ) | ( n12633 & n12860 ) | ( ~n12662 & n12860 ) ;
  assign n12863 = ( n12662 & ~n12861 ) | ( n12662 & n12862 ) | ( ~n12861 & n12862 ) ;
  assign n12864 = ( n12636 & ~n12652 ) | ( n12636 & n12863 ) | ( ~n12652 & n12863 ) ;
  assign n12865 = ( n12636 & n12652 ) | ( n12636 & n12863 ) | ( n12652 & n12863 ) ;
  assign n12866 = ( n12652 & n12864 ) | ( n12652 & ~n12865 ) | ( n12864 & ~n12865 ) ;
  assign n12867 = ( n12639 & n12642 ) | ( n12639 & n12866 ) | ( n12642 & n12866 ) ;
  assign n12868 = ( n12639 & ~n12642 ) | ( n12639 & n12866 ) | ( ~n12642 & n12866 ) ;
  assign n12869 = ( n12642 & ~n12867 ) | ( n12642 & n12868 ) | ( ~n12867 & n12868 ) ;
  assign n12870 = n874 & n9038 ;
  assign n12871 = x17 & n12870 ;
  assign n12872 = x126 & n881 ;
  assign n12873 = x125 & n878 ;
  assign n12874 = n12872 | n12873 ;
  assign n12875 = x124 & n959 ;
  assign n12876 = n12874 | n12875 ;
  assign n12877 = ( ~x17 & n12870 ) | ( ~x17 & n12876 ) | ( n12870 & n12876 ) ;
  assign n12878 = x17 & ~n12876 ;
  assign n12879 = ( ~n12871 & n12877 ) | ( ~n12871 & n12878 ) | ( n12877 & n12878 ) ;
  assign n12880 = n1146 & n8461 ;
  assign n12881 = x20 & n12880 ;
  assign n12882 = x123 & n1153 ;
  assign n12883 = x122 & n1150 ;
  assign n12884 = n12882 | n12883 ;
  assign n12885 = x121 & n1217 ;
  assign n12886 = n12884 | n12885 ;
  assign n12887 = ( ~x20 & n12880 ) | ( ~x20 & n12886 ) | ( n12880 & n12886 ) ;
  assign n12888 = x20 & ~n12886 ;
  assign n12889 = ( ~n12881 & n12887 ) | ( ~n12881 & n12888 ) | ( n12887 & n12888 ) ;
  assign n12890 = n1427 & n7444 ;
  assign n12891 = x23 & n12890 ;
  assign n12892 = x120 & n1434 ;
  assign n12893 = x119 & n1431 ;
  assign n12894 = n12892 | n12893 ;
  assign n12895 = x118 & n1531 ;
  assign n12896 = n12894 | n12895 ;
  assign n12897 = ( ~x23 & n12890 ) | ( ~x23 & n12896 ) | ( n12890 & n12896 ) ;
  assign n12898 = x23 & ~n12896 ;
  assign n12899 = ( ~n12891 & n12897 ) | ( ~n12891 & n12898 ) | ( n12897 & n12898 ) ;
  assign n12900 = n1755 & n6924 ;
  assign n12901 = x26 & n12900 ;
  assign n12902 = x117 & n1762 ;
  assign n12903 = x116 & n1759 ;
  assign n12904 = n12902 | n12903 ;
  assign n12905 = x115 & n1895 ;
  assign n12906 = n12904 | n12905 ;
  assign n12907 = ( ~x26 & n12900 ) | ( ~x26 & n12906 ) | ( n12900 & n12906 ) ;
  assign n12908 = x26 & ~n12906 ;
  assign n12909 = ( ~n12901 & n12907 ) | ( ~n12901 & n12908 ) | ( n12907 & n12908 ) ;
  assign n12910 = n2137 & n6002 ;
  assign n12911 = x29 & n12910 ;
  assign n12912 = x114 & n2144 ;
  assign n12913 = x113 & n2141 ;
  assign n12914 = n12912 | n12913 ;
  assign n12915 = x112 & n2267 ;
  assign n12916 = n12914 | n12915 ;
  assign n12917 = ( ~x29 & n12910 ) | ( ~x29 & n12916 ) | ( n12910 & n12916 ) ;
  assign n12918 = x29 & ~n12916 ;
  assign n12919 = ( ~n12911 & n12917 ) | ( ~n12911 & n12918 ) | ( n12917 & n12918 ) ;
  assign n12920 = n2545 & n5347 ;
  assign n12921 = x32 & n12920 ;
  assign n12922 = x111 & n2552 ;
  assign n12923 = x110 & n2549 ;
  assign n12924 = n12922 | n12923 ;
  assign n12925 = x109 & n2696 ;
  assign n12926 = n12924 | n12925 ;
  assign n12927 = ( ~x32 & n12920 ) | ( ~x32 & n12926 ) | ( n12920 & n12926 ) ;
  assign n12928 = x32 & ~n12926 ;
  assign n12929 = ( ~n12921 & n12927 ) | ( ~n12921 & n12928 ) | ( n12927 & n12928 ) ;
  assign n12930 = n2982 & n4914 ;
  assign n12931 = x35 & n12930 ;
  assign n12932 = x108 & n2989 ;
  assign n12933 = x107 & n2986 ;
  assign n12934 = n12932 | n12933 ;
  assign n12935 = x106 & n3159 ;
  assign n12936 = n12934 | n12935 ;
  assign n12937 = ( ~x35 & n12930 ) | ( ~x35 & n12936 ) | ( n12930 & n12936 ) ;
  assign n12938 = x35 & ~n12936 ;
  assign n12939 = ( ~n12931 & n12937 ) | ( ~n12931 & n12938 ) | ( n12937 & n12938 ) ;
  assign n12940 = n3492 & n4145 ;
  assign n12941 = x38 & n12940 ;
  assign n12942 = x105 & n3499 ;
  assign n12943 = x104 & n3496 ;
  assign n12944 = n12942 | n12943 ;
  assign n12945 = x103 & n3662 ;
  assign n12946 = n12944 | n12945 ;
  assign n12947 = ( ~x38 & n12940 ) | ( ~x38 & n12946 ) | ( n12940 & n12946 ) ;
  assign n12948 = x38 & ~n12946 ;
  assign n12949 = ( ~n12941 & n12947 ) | ( ~n12941 & n12948 ) | ( n12947 & n12948 ) ;
  assign n12950 = n3764 & n4020 ;
  assign n12951 = x41 & n12950 ;
  assign n12952 = x102 & n4027 ;
  assign n12953 = x101 & n4024 ;
  assign n12954 = n12952 | n12953 ;
  assign n12955 = x100 & n4223 ;
  assign n12956 = n12954 | n12955 ;
  assign n12957 = ( ~x41 & n12950 ) | ( ~x41 & n12956 ) | ( n12950 & n12956 ) ;
  assign n12958 = x41 & ~n12956 ;
  assign n12959 = ( ~n12951 & n12957 ) | ( ~n12951 & n12958 ) | ( n12957 & n12958 ) ;
  assign n12960 = n3248 & n4625 ;
  assign n12961 = x44 & n12960 ;
  assign n12962 = x99 & n4791 ;
  assign n12963 = x98 & n4621 ;
  assign n12964 = n12962 | n12963 ;
  assign n12965 = x97 & n4795 ;
  assign n12966 = n12964 | n12965 ;
  assign n12967 = ( ~x44 & n12960 ) | ( ~x44 & n12966 ) | ( n12960 & n12966 ) ;
  assign n12968 = x44 & ~n12966 ;
  assign n12969 = ( ~n12961 & n12967 ) | ( ~n12961 & n12968 ) | ( n12967 & n12968 ) ;
  assign n12970 = n2772 & n5223 ;
  assign n12971 = x47 & n12970 ;
  assign n12972 = x96 & n5230 ;
  assign n12973 = x95 & n5227 ;
  assign n12974 = n12972 | n12973 ;
  assign n12975 = x94 & n5434 ;
  assign n12976 = n12974 | n12975 ;
  assign n12977 = ( ~x47 & n12970 ) | ( ~x47 & n12976 ) | ( n12970 & n12976 ) ;
  assign n12978 = x47 & ~n12976 ;
  assign n12979 = ( ~n12971 & n12977 ) | ( ~n12971 & n12978 ) | ( n12977 & n12978 ) ;
  assign n12980 = n2220 & n5858 ;
  assign n12981 = x50 & n12980 ;
  assign n12982 = x93 & n5865 ;
  assign n12983 = x92 & n5862 ;
  assign n12984 = n12982 | n12983 ;
  assign n12985 = x91 & n6092 ;
  assign n12986 = n12984 | n12985 ;
  assign n12987 = ( ~x50 & n12980 ) | ( ~x50 & n12986 ) | ( n12980 & n12986 ) ;
  assign n12988 = x50 & ~n12986 ;
  assign n12989 = ( ~n12981 & n12987 ) | ( ~n12981 & n12988 ) | ( n12987 & n12988 ) ;
  assign n12990 = n1838 & n6546 ;
  assign n12991 = x53 & n12990 ;
  assign n12992 = x90 & n6553 ;
  assign n12993 = x89 & n6550 ;
  assign n12994 = n12992 | n12993 ;
  assign n12995 = x88 & n6787 ;
  assign n12996 = n12994 | n12995 ;
  assign n12997 = ( ~x53 & n12990 ) | ( ~x53 & n12996 ) | ( n12990 & n12996 ) ;
  assign n12998 = x53 & ~n12996 ;
  assign n12999 = ( ~n12991 & n12997 ) | ( ~n12991 & n12998 ) | ( n12997 & n12998 ) ;
  assign n13000 = n1494 & n7277 ;
  assign n13001 = x56 & n13000 ;
  assign n13002 = x87 & n7545 ;
  assign n13003 = x86 & n7273 ;
  assign n13004 = n13002 | n13003 ;
  assign n13005 = x85 & n7552 ;
  assign n13006 = n13004 | n13005 ;
  assign n13007 = ( ~x56 & n13000 ) | ( ~x56 & n13006 ) | ( n13000 & n13006 ) ;
  assign n13008 = x56 & ~n13006 ;
  assign n13009 = ( ~n13001 & n13007 ) | ( ~n13001 & n13008 ) | ( n13007 & n13008 ) ;
  assign n13010 = n1190 & n8067 ;
  assign n13011 = x59 & n13010 ;
  assign n13012 = x84 & n8074 ;
  assign n13013 = x83 & n8071 ;
  assign n13014 = n13012 | n13013 ;
  assign n13015 = x82 & n8298 ;
  assign n13016 = n13014 | n13015 ;
  assign n13017 = ( ~x59 & n13010 ) | ( ~x59 & n13016 ) | ( n13010 & n13016 ) ;
  assign n13018 = x59 & ~n13016 ;
  assign n13019 = ( ~n13011 & n13017 ) | ( ~n13011 & n13018 ) | ( n13017 & n13018 ) ;
  assign n13020 = n990 & n8859 ;
  assign n13021 = x62 & n13020 ;
  assign n13022 = x81 & n8866 ;
  assign n13023 = x80 & n8863 ;
  assign n13024 = n13022 | n13023 ;
  assign n13025 = x79 & n9125 ;
  assign n13026 = n13024 | n13025 ;
  assign n13027 = ( ~x62 & n13020 ) | ( ~x62 & n13026 ) | ( n13020 & n13026 ) ;
  assign n13028 = x62 & ~n13026 ;
  assign n13029 = ( ~n13021 & n13027 ) | ( ~n13021 & n13028 ) | ( n13027 & n13028 ) ;
  assign n13030 = ( x62 & x63 ) | ( x62 & x78 ) | ( x63 & x78 ) ;
  assign n13031 = ( x62 & x77 ) | ( x62 & ~n9394 ) | ( x77 & ~n9394 ) ;
  assign n13032 = ( x77 & n13030 ) | ( x77 & ~n13031 ) | ( n13030 & ~n13031 ) ;
  assign n13033 = ( ~n12815 & n13029 ) | ( ~n12815 & n13032 ) | ( n13029 & n13032 ) ;
  assign n13034 = ( n12815 & n13029 ) | ( n12815 & n13032 ) | ( n13029 & n13032 ) ;
  assign n13035 = ( n12815 & n13033 ) | ( n12815 & ~n13034 ) | ( n13033 & ~n13034 ) ;
  assign n13036 = ( n12816 & ~n13019 ) | ( n12816 & n13035 ) | ( ~n13019 & n13035 ) ;
  assign n13037 = ( n12816 & n13019 ) | ( n12816 & ~n13035 ) | ( n13019 & ~n13035 ) ;
  assign n13038 = ( ~n12816 & n13036 ) | ( ~n12816 & n13037 ) | ( n13036 & n13037 ) ;
  assign n13039 = ( n12819 & n13009 ) | ( n12819 & ~n13038 ) | ( n13009 & ~n13038 ) ;
  assign n13040 = ( ~n12819 & n13009 ) | ( ~n12819 & n13038 ) | ( n13009 & n13038 ) ;
  assign n13041 = ( ~n13009 & n13039 ) | ( ~n13009 & n13040 ) | ( n13039 & n13040 ) ;
  assign n13042 = ( n12822 & n12999 ) | ( n12822 & ~n13041 ) | ( n12999 & ~n13041 ) ;
  assign n13043 = ( ~n12822 & n12999 ) | ( ~n12822 & n13041 ) | ( n12999 & n13041 ) ;
  assign n13044 = ( ~n12999 & n13042 ) | ( ~n12999 & n13043 ) | ( n13042 & n13043 ) ;
  assign n13045 = ( n12826 & ~n12989 ) | ( n12826 & n13044 ) | ( ~n12989 & n13044 ) ;
  assign n13046 = ( n12826 & n12989 ) | ( n12826 & n13044 ) | ( n12989 & n13044 ) ;
  assign n13047 = ( n12989 & n13045 ) | ( n12989 & ~n13046 ) | ( n13045 & ~n13046 ) ;
  assign n13048 = ( n12829 & n12979 ) | ( n12829 & n13047 ) | ( n12979 & n13047 ) ;
  assign n13049 = ( n12829 & ~n12979 ) | ( n12829 & n13047 ) | ( ~n12979 & n13047 ) ;
  assign n13050 = ( n12979 & ~n13048 ) | ( n12979 & n13049 ) | ( ~n13048 & n13049 ) ;
  assign n13051 = ( n12832 & n12969 ) | ( n12832 & n13050 ) | ( n12969 & n13050 ) ;
  assign n13052 = ( n12832 & ~n12969 ) | ( n12832 & n13050 ) | ( ~n12969 & n13050 ) ;
  assign n13053 = ( n12969 & ~n13051 ) | ( n12969 & n13052 ) | ( ~n13051 & n13052 ) ;
  assign n13054 = ( n12835 & n12959 ) | ( n12835 & n13053 ) | ( n12959 & n13053 ) ;
  assign n13055 = ( n12835 & ~n12959 ) | ( n12835 & n13053 ) | ( ~n12959 & n13053 ) ;
  assign n13056 = ( n12959 & ~n13054 ) | ( n12959 & n13055 ) | ( ~n13054 & n13055 ) ;
  assign n13057 = ( n12837 & n12949 ) | ( n12837 & n13056 ) | ( n12949 & n13056 ) ;
  assign n13058 = ( n12837 & ~n12949 ) | ( n12837 & n13056 ) | ( ~n12949 & n13056 ) ;
  assign n13059 = ( n12949 & ~n13057 ) | ( n12949 & n13058 ) | ( ~n13057 & n13058 ) ;
  assign n13060 = ( n12840 & n12939 ) | ( n12840 & n13059 ) | ( n12939 & n13059 ) ;
  assign n13061 = ( n12840 & ~n12939 ) | ( n12840 & n13059 ) | ( ~n12939 & n13059 ) ;
  assign n13062 = ( n12939 & ~n13060 ) | ( n12939 & n13061 ) | ( ~n13060 & n13061 ) ;
  assign n13063 = ( n12843 & n12929 ) | ( n12843 & n13062 ) | ( n12929 & n13062 ) ;
  assign n13064 = ( n12843 & ~n12929 ) | ( n12843 & n13062 ) | ( ~n12929 & n13062 ) ;
  assign n13065 = ( n12929 & ~n13063 ) | ( n12929 & n13064 ) | ( ~n13063 & n13064 ) ;
  assign n13066 = ( n12847 & n12919 ) | ( n12847 & n13065 ) | ( n12919 & n13065 ) ;
  assign n13067 = ( n12847 & ~n12919 ) | ( n12847 & n13065 ) | ( ~n12919 & n13065 ) ;
  assign n13068 = ( n12919 & ~n13066 ) | ( n12919 & n13067 ) | ( ~n13066 & n13067 ) ;
  assign n13069 = ( n12849 & n12909 ) | ( n12849 & n13068 ) | ( n12909 & n13068 ) ;
  assign n13070 = ( n12849 & ~n12909 ) | ( n12849 & n13068 ) | ( ~n12909 & n13068 ) ;
  assign n13071 = ( n12909 & ~n13069 ) | ( n12909 & n13070 ) | ( ~n13069 & n13070 ) ;
  assign n13072 = ( n12852 & n12899 ) | ( n12852 & n13071 ) | ( n12899 & n13071 ) ;
  assign n13073 = ( n12852 & ~n12899 ) | ( n12852 & n13071 ) | ( ~n12899 & n13071 ) ;
  assign n13074 = ( n12899 & ~n13072 ) | ( n12899 & n13073 ) | ( ~n13072 & n13073 ) ;
  assign n13075 = ( n12855 & ~n12889 ) | ( n12855 & n13074 ) | ( ~n12889 & n13074 ) ;
  assign n13076 = ( n12855 & n12889 ) | ( n12855 & n13074 ) | ( n12889 & n13074 ) ;
  assign n13077 = ( n12889 & n13075 ) | ( n12889 & ~n13076 ) | ( n13075 & ~n13076 ) ;
  assign n13078 = ( n12858 & ~n12879 ) | ( n12858 & n13077 ) | ( ~n12879 & n13077 ) ;
  assign n13079 = ( n12858 & n12879 ) | ( n12858 & n13077 ) | ( n12879 & n13077 ) ;
  assign n13080 = ( n12879 & n13078 ) | ( n12879 & ~n13079 ) | ( n13078 & ~n13079 ) ;
  assign n13081 = x127 & n744 ;
  assign n13082 = n649 | n13081 ;
  assign n13083 = ( n9865 & n13081 ) | ( n9865 & n13082 ) | ( n13081 & n13082 ) ;
  assign n13084 = x14 & ~n13083 ;
  assign n13085 = ~x14 & n13083 ;
  assign n13086 = n13084 | n13085 ;
  assign n13087 = ( n12861 & n13080 ) | ( n12861 & n13086 ) | ( n13080 & n13086 ) ;
  assign n13088 = ( n12861 & ~n13080 ) | ( n12861 & n13086 ) | ( ~n13080 & n13086 ) ;
  assign n13089 = ( n13080 & ~n13087 ) | ( n13080 & n13088 ) | ( ~n13087 & n13088 ) ;
  assign n13090 = ( n12865 & n12867 ) | ( n12865 & n13089 ) | ( n12867 & n13089 ) ;
  assign n13091 = ( n12865 & ~n12867 ) | ( n12865 & n13089 ) | ( ~n12867 & n13089 ) ;
  assign n13092 = ( n12867 & ~n13090 ) | ( n12867 & n13091 ) | ( ~n13090 & n13091 ) ;
  assign n13093 = n874 & n9576 ;
  assign n13094 = x17 & n13093 ;
  assign n13095 = x127 & n881 ;
  assign n13096 = x126 & n878 ;
  assign n13097 = n13095 | n13096 ;
  assign n13098 = x125 & n959 ;
  assign n13099 = n13097 | n13098 ;
  assign n13100 = ( ~x17 & n13093 ) | ( ~x17 & n13099 ) | ( n13093 & n13099 ) ;
  assign n13101 = x17 & ~n13099 ;
  assign n13102 = ( ~n13094 & n13100 ) | ( ~n13094 & n13101 ) | ( n13100 & n13101 ) ;
  assign n13103 = n1146 & n8729 ;
  assign n13104 = x20 & n13103 ;
  assign n13105 = x124 & n1153 ;
  assign n13106 = x123 & n1150 ;
  assign n13107 = n13105 | n13106 ;
  assign n13108 = x122 & n1217 ;
  assign n13109 = n13107 | n13108 ;
  assign n13110 = ( ~x20 & n13103 ) | ( ~x20 & n13109 ) | ( n13103 & n13109 ) ;
  assign n13111 = x20 & ~n13109 ;
  assign n13112 = ( ~n13104 & n13110 ) | ( ~n13104 & n13111 ) | ( n13110 & n13111 ) ;
  assign n13113 = n1427 & n7696 ;
  assign n13114 = x23 & n13113 ;
  assign n13115 = x121 & n1434 ;
  assign n13116 = x120 & n1431 ;
  assign n13117 = n13115 | n13116 ;
  assign n13118 = x119 & n1531 ;
  assign n13119 = n13117 | n13118 ;
  assign n13120 = ( ~x23 & n13113 ) | ( ~x23 & n13119 ) | ( n13113 & n13119 ) ;
  assign n13121 = x23 & ~n13119 ;
  assign n13122 = ( ~n13114 & n13120 ) | ( ~n13114 & n13121 ) | ( n13120 & n13121 ) ;
  assign n13123 = n1755 & n6940 ;
  assign n13124 = x26 & n13123 ;
  assign n13125 = x118 & n1762 ;
  assign n13126 = x117 & n1759 ;
  assign n13127 = n13125 | n13126 ;
  assign n13128 = x116 & n1895 ;
  assign n13129 = n13127 | n13128 ;
  assign n13130 = ( ~x26 & n13123 ) | ( ~x26 & n13129 ) | ( n13123 & n13129 ) ;
  assign n13131 = x26 & ~n13129 ;
  assign n13132 = ( ~n13124 & n13130 ) | ( ~n13124 & n13131 ) | ( n13130 & n13131 ) ;
  assign n13133 = n2137 & n6446 ;
  assign n13134 = x29 & n13133 ;
  assign n13135 = x115 & n2144 ;
  assign n13136 = x114 & n2141 ;
  assign n13137 = n13135 | n13136 ;
  assign n13138 = x113 & n2267 ;
  assign n13139 = n13137 | n13138 ;
  assign n13140 = ( ~x29 & n13133 ) | ( ~x29 & n13139 ) | ( n13133 & n13139 ) ;
  assign n13141 = x29 & ~n13139 ;
  assign n13142 = ( ~n13134 & n13140 ) | ( ~n13134 & n13141 ) | ( n13140 & n13141 ) ;
  assign n13143 = n2545 & n5558 ;
  assign n13144 = x32 & n13143 ;
  assign n13145 = x112 & n2552 ;
  assign n13146 = x111 & n2549 ;
  assign n13147 = n13145 | n13146 ;
  assign n13148 = x110 & n2696 ;
  assign n13149 = n13147 | n13148 ;
  assign n13150 = ( ~x32 & n13143 ) | ( ~x32 & n13149 ) | ( n13143 & n13149 ) ;
  assign n13151 = x32 & ~n13149 ;
  assign n13152 = ( ~n13144 & n13150 ) | ( ~n13144 & n13151 ) | ( n13150 & n13151 ) ;
  assign n13153 = n2982 & n4930 ;
  assign n13154 = x35 & n13153 ;
  assign n13155 = x109 & n2989 ;
  assign n13156 = x108 & n2986 ;
  assign n13157 = n13155 | n13156 ;
  assign n13158 = x107 & n3159 ;
  assign n13159 = n13157 | n13158 ;
  assign n13160 = ( ~x35 & n13153 ) | ( ~x35 & n13159 ) | ( n13153 & n13159 ) ;
  assign n13161 = x35 & ~n13159 ;
  assign n13162 = ( ~n13154 & n13160 ) | ( ~n13154 & n13161 ) | ( n13160 & n13161 ) ;
  assign n13163 = n3492 & n4331 ;
  assign n13164 = x38 & n13163 ;
  assign n13165 = x106 & n3499 ;
  assign n13166 = x105 & n3496 ;
  assign n13167 = n13165 | n13166 ;
  assign n13168 = x104 & n3662 ;
  assign n13169 = n13167 | n13168 ;
  assign n13170 = ( ~x38 & n13163 ) | ( ~x38 & n13169 ) | ( n13163 & n13169 ) ;
  assign n13171 = x38 & ~n13169 ;
  assign n13172 = ( ~n13164 & n13170 ) | ( ~n13164 & n13171 ) | ( n13170 & n13171 ) ;
  assign n13173 = n3941 & n4020 ;
  assign n13174 = x41 & n13173 ;
  assign n13175 = x103 & n4027 ;
  assign n13176 = x102 & n4024 ;
  assign n13177 = n13175 | n13176 ;
  assign n13178 = x101 & n4223 ;
  assign n13179 = n13177 | n13178 ;
  assign n13180 = ( ~x41 & n13173 ) | ( ~x41 & n13179 ) | ( n13173 & n13179 ) ;
  assign n13181 = x41 & ~n13179 ;
  assign n13182 = ( ~n13174 & n13180 ) | ( ~n13174 & n13181 ) | ( n13180 & n13181 ) ;
  assign n13183 = n3264 & n4625 ;
  assign n13184 = x44 & n13183 ;
  assign n13185 = x100 & n4791 ;
  assign n13186 = x99 & n4621 ;
  assign n13187 = n13185 | n13186 ;
  assign n13188 = x98 & n4795 ;
  assign n13189 = n13187 | n13188 ;
  assign n13190 = ( ~x44 & n13183 ) | ( ~x44 & n13189 ) | ( n13183 & n13189 ) ;
  assign n13191 = x44 & ~n13189 ;
  assign n13192 = ( ~n13184 & n13190 ) | ( ~n13184 & n13191 ) | ( n13190 & n13191 ) ;
  assign n13193 = n2788 & n5223 ;
  assign n13194 = x47 & n13193 ;
  assign n13195 = x97 & n5230 ;
  assign n13196 = x96 & n5227 ;
  assign n13197 = n13195 | n13196 ;
  assign n13198 = x95 & n5434 ;
  assign n13199 = n13197 | n13198 ;
  assign n13200 = ( ~x47 & n13193 ) | ( ~x47 & n13199 ) | ( n13193 & n13199 ) ;
  assign n13201 = x47 & ~n13199 ;
  assign n13202 = ( ~n13194 & n13200 ) | ( ~n13194 & n13201 ) | ( n13200 & n13201 ) ;
  assign n13203 = n2476 & n5858 ;
  assign n13204 = x50 & n13203 ;
  assign n13205 = x94 & n5865 ;
  assign n13206 = x93 & n5862 ;
  assign n13207 = n13205 | n13206 ;
  assign n13208 = x92 & n6092 ;
  assign n13209 = n13207 | n13208 ;
  assign n13210 = ( ~x50 & n13203 ) | ( ~x50 & n13209 ) | ( n13203 & n13209 ) ;
  assign n13211 = x50 & ~n13209 ;
  assign n13212 = ( ~n13204 & n13210 ) | ( ~n13204 & n13211 ) | ( n13210 & n13211 ) ;
  assign n13213 = n1959 & n6546 ;
  assign n13214 = x53 & n13213 ;
  assign n13215 = x91 & n6553 ;
  assign n13216 = x90 & n6550 ;
  assign n13217 = n13215 | n13216 ;
  assign n13218 = x89 & n6787 ;
  assign n13219 = n13217 | n13218 ;
  assign n13220 = ( ~x53 & n13213 ) | ( ~x53 & n13219 ) | ( n13213 & n13219 ) ;
  assign n13221 = x53 & ~n13219 ;
  assign n13222 = ( ~n13214 & n13220 ) | ( ~n13214 & n13221 ) | ( n13220 & n13221 ) ;
  assign n13223 = n1602 & n7277 ;
  assign n13224 = x56 & n13223 ;
  assign n13225 = x88 & n7545 ;
  assign n13226 = x87 & n7273 ;
  assign n13227 = n13225 | n13226 ;
  assign n13228 = x86 & n7552 ;
  assign n13229 = n13227 | n13228 ;
  assign n13230 = ( ~x56 & n13223 ) | ( ~x56 & n13229 ) | ( n13223 & n13229 ) ;
  assign n13231 = x56 & ~n13229 ;
  assign n13232 = ( ~n13224 & n13230 ) | ( ~n13224 & n13231 ) | ( n13230 & n13231 ) ;
  assign n13233 = n1368 & n8067 ;
  assign n13234 = x59 & n13233 ;
  assign n13235 = x85 & n8074 ;
  assign n13236 = x84 & n8071 ;
  assign n13237 = n13235 | n13236 ;
  assign n13238 = x83 & n8298 ;
  assign n13239 = n13237 | n13238 ;
  assign n13240 = ( ~x59 & n13233 ) | ( ~x59 & n13239 ) | ( n13233 & n13239 ) ;
  assign n13241 = x59 & ~n13239 ;
  assign n13242 = ( ~n13234 & n13240 ) | ( ~n13234 & n13241 ) | ( n13240 & n13241 ) ;
  assign n13243 = n1006 & n8859 ;
  assign n13244 = x62 & n13243 ;
  assign n13245 = x82 & n8866 ;
  assign n13246 = x81 & n8863 ;
  assign n13247 = n13245 | n13246 ;
  assign n13248 = x80 & n9125 ;
  assign n13249 = n13247 | n13248 ;
  assign n13250 = ( ~x62 & n13243 ) | ( ~x62 & n13249 ) | ( n13243 & n13249 ) ;
  assign n13251 = x62 & ~n13249 ;
  assign n13252 = ( ~n13244 & n13250 ) | ( ~n13244 & n13251 ) | ( n13250 & n13251 ) ;
  assign n13253 = ( x62 & x63 ) | ( x62 & x79 ) | ( x63 & x79 ) ;
  assign n13254 = ( x62 & x78 ) | ( x62 & ~n9394 ) | ( x78 & ~n9394 ) ;
  assign n13255 = ( x78 & n13253 ) | ( x78 & ~n13254 ) | ( n13253 & ~n13254 ) ;
  assign n13256 = ( x14 & n12815 ) | ( x14 & n13255 ) | ( n12815 & n13255 ) ;
  assign n13257 = ( ~x14 & n12815 ) | ( ~x14 & n13255 ) | ( n12815 & n13255 ) ;
  assign n13258 = ( x14 & ~n13256 ) | ( x14 & n13257 ) | ( ~n13256 & n13257 ) ;
  assign n13259 = ( n13033 & n13252 ) | ( n13033 & ~n13258 ) | ( n13252 & ~n13258 ) ;
  assign n13260 = ( n13033 & ~n13252 ) | ( n13033 & n13258 ) | ( ~n13252 & n13258 ) ;
  assign n13261 = ( ~n13033 & n13259 ) | ( ~n13033 & n13260 ) | ( n13259 & n13260 ) ;
  assign n13262 = ( n13037 & n13242 ) | ( n13037 & ~n13261 ) | ( n13242 & ~n13261 ) ;
  assign n13263 = ( n13037 & ~n13242 ) | ( n13037 & n13261 ) | ( ~n13242 & n13261 ) ;
  assign n13264 = ( ~n13037 & n13262 ) | ( ~n13037 & n13263 ) | ( n13262 & n13263 ) ;
  assign n13265 = ( n13039 & n13232 ) | ( n13039 & ~n13264 ) | ( n13232 & ~n13264 ) ;
  assign n13266 = ( n13039 & ~n13232 ) | ( n13039 & n13264 ) | ( ~n13232 & n13264 ) ;
  assign n13267 = ( ~n13039 & n13265 ) | ( ~n13039 & n13266 ) | ( n13265 & n13266 ) ;
  assign n13268 = ( n13042 & n13222 ) | ( n13042 & ~n13267 ) | ( n13222 & ~n13267 ) ;
  assign n13269 = ( n13042 & ~n13222 ) | ( n13042 & n13267 ) | ( ~n13222 & n13267 ) ;
  assign n13270 = ( ~n13042 & n13268 ) | ( ~n13042 & n13269 ) | ( n13268 & n13269 ) ;
  assign n13271 = ( n13045 & ~n13212 ) | ( n13045 & n13270 ) | ( ~n13212 & n13270 ) ;
  assign n13272 = ( n13045 & n13212 ) | ( n13045 & n13270 ) | ( n13212 & n13270 ) ;
  assign n13273 = ( n13212 & n13271 ) | ( n13212 & ~n13272 ) | ( n13271 & ~n13272 ) ;
  assign n13274 = ( n13048 & n13202 ) | ( n13048 & n13273 ) | ( n13202 & n13273 ) ;
  assign n13275 = ( n13048 & ~n13202 ) | ( n13048 & n13273 ) | ( ~n13202 & n13273 ) ;
  assign n13276 = ( n13202 & ~n13274 ) | ( n13202 & n13275 ) | ( ~n13274 & n13275 ) ;
  assign n13277 = ( n13051 & n13192 ) | ( n13051 & n13276 ) | ( n13192 & n13276 ) ;
  assign n13278 = ( ~n13051 & n13192 ) | ( ~n13051 & n13276 ) | ( n13192 & n13276 ) ;
  assign n13279 = ( n13051 & ~n13277 ) | ( n13051 & n13278 ) | ( ~n13277 & n13278 ) ;
  assign n13280 = ( n13054 & n13182 ) | ( n13054 & n13279 ) | ( n13182 & n13279 ) ;
  assign n13281 = ( n13054 & ~n13182 ) | ( n13054 & n13279 ) | ( ~n13182 & n13279 ) ;
  assign n13282 = ( n13182 & ~n13280 ) | ( n13182 & n13281 ) | ( ~n13280 & n13281 ) ;
  assign n13283 = ( n13057 & n13172 ) | ( n13057 & n13282 ) | ( n13172 & n13282 ) ;
  assign n13284 = ( ~n13057 & n13172 ) | ( ~n13057 & n13282 ) | ( n13172 & n13282 ) ;
  assign n13285 = ( n13057 & ~n13283 ) | ( n13057 & n13284 ) | ( ~n13283 & n13284 ) ;
  assign n13286 = ( n13060 & n13162 ) | ( n13060 & n13285 ) | ( n13162 & n13285 ) ;
  assign n13287 = ( ~n13060 & n13162 ) | ( ~n13060 & n13285 ) | ( n13162 & n13285 ) ;
  assign n13288 = ( n13060 & ~n13286 ) | ( n13060 & n13287 ) | ( ~n13286 & n13287 ) ;
  assign n13289 = ( n13063 & n13152 ) | ( n13063 & n13288 ) | ( n13152 & n13288 ) ;
  assign n13290 = ( n13063 & ~n13152 ) | ( n13063 & n13288 ) | ( ~n13152 & n13288 ) ;
  assign n13291 = ( n13152 & ~n13289 ) | ( n13152 & n13290 ) | ( ~n13289 & n13290 ) ;
  assign n13292 = ( n13066 & ~n13142 ) | ( n13066 & n13291 ) | ( ~n13142 & n13291 ) ;
  assign n13293 = ( n13066 & n13142 ) | ( n13066 & n13291 ) | ( n13142 & n13291 ) ;
  assign n13294 = ( n13142 & n13292 ) | ( n13142 & ~n13293 ) | ( n13292 & ~n13293 ) ;
  assign n13295 = ( n13069 & n13132 ) | ( n13069 & n13294 ) | ( n13132 & n13294 ) ;
  assign n13296 = ( ~n13069 & n13132 ) | ( ~n13069 & n13294 ) | ( n13132 & n13294 ) ;
  assign n13297 = ( n13069 & ~n13295 ) | ( n13069 & n13296 ) | ( ~n13295 & n13296 ) ;
  assign n13298 = ( n13072 & n13122 ) | ( n13072 & n13297 ) | ( n13122 & n13297 ) ;
  assign n13299 = ( ~n13072 & n13122 ) | ( ~n13072 & n13297 ) | ( n13122 & n13297 ) ;
  assign n13300 = ( n13072 & ~n13298 ) | ( n13072 & n13299 ) | ( ~n13298 & n13299 ) ;
  assign n13301 = ( n13076 & n13112 ) | ( n13076 & n13300 ) | ( n13112 & n13300 ) ;
  assign n13302 = ( ~n13076 & n13112 ) | ( ~n13076 & n13300 ) | ( n13112 & n13300 ) ;
  assign n13303 = ( n13076 & ~n13301 ) | ( n13076 & n13302 ) | ( ~n13301 & n13302 ) ;
  assign n13304 = ( n13079 & n13102 ) | ( n13079 & n13303 ) | ( n13102 & n13303 ) ;
  assign n13305 = ( ~n13079 & n13102 ) | ( ~n13079 & n13303 ) | ( n13102 & n13303 ) ;
  assign n13306 = ( n13079 & ~n13304 ) | ( n13079 & n13305 ) | ( ~n13304 & n13305 ) ;
  assign n13307 = ( n13087 & n13090 ) | ( n13087 & n13306 ) | ( n13090 & n13306 ) ;
  assign n13308 = ( n13087 & ~n13090 ) | ( n13087 & n13306 ) | ( ~n13090 & n13306 ) ;
  assign n13309 = ( n13090 & ~n13307 ) | ( n13090 & n13308 ) | ( ~n13307 & n13308 ) ;
  assign n13310 = x127 & n878 ;
  assign n13311 = n874 | n13310 ;
  assign n13312 = ( n9867 & n13310 ) | ( n9867 & n13311 ) | ( n13310 & n13311 ) ;
  assign n13313 = x126 & n959 ;
  assign n13314 = ( ~x17 & n13312 ) | ( ~x17 & n13313 ) | ( n13312 & n13313 ) ;
  assign n13315 = ( x17 & ~n13312 ) | ( x17 & n13313 ) | ( ~n13312 & n13313 ) ;
  assign n13316 = ~n13313 & n13315 ;
  assign n13317 = n13314 | n13316 ;
  assign n13318 = n1146 & n9009 ;
  assign n13319 = x20 & n13318 ;
  assign n13320 = x125 & n1153 ;
  assign n13321 = x124 & n1150 ;
  assign n13322 = n13320 | n13321 ;
  assign n13323 = x123 & n1217 ;
  assign n13324 = n13322 | n13323 ;
  assign n13325 = ( ~x20 & n13318 ) | ( ~x20 & n13324 ) | ( n13318 & n13324 ) ;
  assign n13326 = x20 & ~n13324 ;
  assign n13327 = ( ~n13319 & n13325 ) | ( ~n13319 & n13326 ) | ( n13325 & n13326 ) ;
  assign n13328 = n1427 & n8207 ;
  assign n13329 = x23 & n13328 ;
  assign n13330 = x122 & n1434 ;
  assign n13331 = x121 & n1431 ;
  assign n13332 = n13330 | n13331 ;
  assign n13333 = x120 & n1531 ;
  assign n13334 = n13332 | n13333 ;
  assign n13335 = ( ~x23 & n13328 ) | ( ~x23 & n13334 ) | ( n13328 & n13334 ) ;
  assign n13336 = x23 & ~n13334 ;
  assign n13337 = ( ~n13329 & n13335 ) | ( ~n13329 & n13336 ) | ( n13335 & n13336 ) ;
  assign n13338 = n1755 & n7181 ;
  assign n13339 = x26 & n13338 ;
  assign n13340 = x119 & n1762 ;
  assign n13341 = x118 & n1759 ;
  assign n13342 = n13340 | n13341 ;
  assign n13343 = x117 & n1895 ;
  assign n13344 = n13342 | n13343 ;
  assign n13345 = ( ~x26 & n13338 ) | ( ~x26 & n13344 ) | ( n13338 & n13344 ) ;
  assign n13346 = x26 & ~n13344 ;
  assign n13347 = ( ~n13339 & n13345 ) | ( ~n13339 & n13346 ) | ( n13345 & n13346 ) ;
  assign n13348 = n2137 & n6462 ;
  assign n13349 = x29 & n13348 ;
  assign n13350 = x116 & n2144 ;
  assign n13351 = x115 & n2141 ;
  assign n13352 = n13350 | n13351 ;
  assign n13353 = x114 & n2267 ;
  assign n13354 = n13352 | n13353 ;
  assign n13355 = ( ~x29 & n13348 ) | ( ~x29 & n13354 ) | ( n13348 & n13354 ) ;
  assign n13356 = x29 & ~n13354 ;
  assign n13357 = ( ~n13349 & n13355 ) | ( ~n13349 & n13356 ) | ( n13355 & n13356 ) ;
  assign n13358 = n2545 & n5774 ;
  assign n13359 = x32 & n13358 ;
  assign n13360 = x113 & n2552 ;
  assign n13361 = x112 & n2549 ;
  assign n13362 = n13360 | n13361 ;
  assign n13363 = x111 & n2696 ;
  assign n13364 = n13362 | n13363 ;
  assign n13365 = ( ~x32 & n13358 ) | ( ~x32 & n13364 ) | ( n13358 & n13364 ) ;
  assign n13366 = x32 & ~n13364 ;
  assign n13367 = ( ~n13359 & n13365 ) | ( ~n13359 & n13366 ) | ( n13365 & n13366 ) ;
  assign n13368 = n2982 & n5331 ;
  assign n13369 = x35 & n13368 ;
  assign n13370 = x110 & n2989 ;
  assign n13371 = x109 & n2986 ;
  assign n13372 = n13370 | n13371 ;
  assign n13373 = x108 & n3159 ;
  assign n13374 = n13372 | n13373 ;
  assign n13375 = ( ~x35 & n13368 ) | ( ~x35 & n13374 ) | ( n13368 & n13374 ) ;
  assign n13376 = x35 & ~n13374 ;
  assign n13377 = ( ~n13369 & n13375 ) | ( ~n13369 & n13376 ) | ( n13375 & n13376 ) ;
  assign n13378 = n3492 & n4523 ;
  assign n13379 = x38 & n13378 ;
  assign n13380 = x107 & n3499 ;
  assign n13381 = x106 & n3496 ;
  assign n13382 = n13380 | n13381 ;
  assign n13383 = x105 & n3662 ;
  assign n13384 = n13382 | n13383 ;
  assign n13385 = ( ~x38 & n13378 ) | ( ~x38 & n13384 ) | ( n13378 & n13384 ) ;
  assign n13386 = x38 & ~n13384 ;
  assign n13387 = ( ~n13379 & n13385 ) | ( ~n13379 & n13386 ) | ( n13385 & n13386 ) ;
  assign n13388 = n3957 & n4020 ;
  assign n13389 = x41 & n13388 ;
  assign n13390 = x104 & n4027 ;
  assign n13391 = x103 & n4024 ;
  assign n13392 = n13390 | n13391 ;
  assign n13393 = x102 & n4223 ;
  assign n13394 = n13392 | n13393 ;
  assign n13395 = ( ~x41 & n13388 ) | ( ~x41 & n13394 ) | ( n13388 & n13394 ) ;
  assign n13396 = x41 & ~n13394 ;
  assign n13397 = ( ~n13389 & n13395 ) | ( ~n13389 & n13396 ) | ( n13395 & n13396 ) ;
  assign n13398 = n3591 & n4625 ;
  assign n13399 = x44 & n13398 ;
  assign n13400 = x101 & n4791 ;
  assign n13401 = x100 & n4621 ;
  assign n13402 = n13400 | n13401 ;
  assign n13403 = x99 & n4795 ;
  assign n13404 = n13402 | n13403 ;
  assign n13405 = ( ~x44 & n13398 ) | ( ~x44 & n13404 ) | ( n13398 & n13404 ) ;
  assign n13406 = x44 & ~n13404 ;
  assign n13407 = ( ~n13399 & n13405 ) | ( ~n13399 & n13406 ) | ( n13405 & n13406 ) ;
  assign n13408 = n2939 & n5223 ;
  assign n13409 = x47 & n13408 ;
  assign n13410 = x98 & n5230 ;
  assign n13411 = x97 & n5227 ;
  assign n13412 = n13410 | n13411 ;
  assign n13413 = x96 & n5434 ;
  assign n13414 = n13412 | n13413 ;
  assign n13415 = ( ~x47 & n13408 ) | ( ~x47 & n13414 ) | ( n13408 & n13414 ) ;
  assign n13416 = x47 & ~n13414 ;
  assign n13417 = ( ~n13409 & n13415 ) | ( ~n13409 & n13416 ) | ( n13415 & n13416 ) ;
  assign n13418 = n2492 & n5858 ;
  assign n13419 = x50 & n13418 ;
  assign n13420 = x95 & n5865 ;
  assign n13421 = x94 & n5862 ;
  assign n13422 = n13420 | n13421 ;
  assign n13423 = x93 & n6092 ;
  assign n13424 = n13422 | n13423 ;
  assign n13425 = ( ~x50 & n13418 ) | ( ~x50 & n13424 ) | ( n13418 & n13424 ) ;
  assign n13426 = x50 & ~n13424 ;
  assign n13427 = ( ~n13419 & n13425 ) | ( ~n13419 & n13426 ) | ( n13425 & n13426 ) ;
  assign n13428 = n2083 & n6546 ;
  assign n13429 = x53 & n13428 ;
  assign n13430 = x92 & n6553 ;
  assign n13431 = x91 & n6550 ;
  assign n13432 = n13430 | n13431 ;
  assign n13433 = x90 & n6787 ;
  assign n13434 = n13432 | n13433 ;
  assign n13435 = ( ~x53 & n13428 ) | ( ~x53 & n13434 ) | ( n13428 & n13434 ) ;
  assign n13436 = x53 & ~n13434 ;
  assign n13437 = ( ~n13429 & n13435 ) | ( ~n13429 & n13436 ) | ( n13435 & n13436 ) ;
  assign n13438 = n1822 & n7277 ;
  assign n13439 = x56 & n13438 ;
  assign n13440 = x89 & n7545 ;
  assign n13441 = x88 & n7273 ;
  assign n13442 = n13440 | n13441 ;
  assign n13443 = x87 & n7552 ;
  assign n13444 = n13442 | n13443 ;
  assign n13445 = ( ~x56 & n13438 ) | ( ~x56 & n13444 ) | ( n13438 & n13444 ) ;
  assign n13446 = x56 & ~n13444 ;
  assign n13447 = ( ~n13439 & n13445 ) | ( ~n13439 & n13446 ) | ( n13445 & n13446 ) ;
  assign n13448 = n1384 & n8067 ;
  assign n13449 = x59 & n13448 ;
  assign n13450 = x86 & n8074 ;
  assign n13451 = x85 & n8071 ;
  assign n13452 = n13450 | n13451 ;
  assign n13453 = x84 & n8298 ;
  assign n13454 = n13452 | n13453 ;
  assign n13455 = ( ~x59 & n13448 ) | ( ~x59 & n13454 ) | ( n13448 & n13454 ) ;
  assign n13456 = x59 & ~n13454 ;
  assign n13457 = ( ~n13449 & n13455 ) | ( ~n13449 & n13456 ) | ( n13455 & n13456 ) ;
  assign n13458 = n1093 & n8859 ;
  assign n13459 = x62 & n13458 ;
  assign n13460 = x83 & n8866 ;
  assign n13461 = x82 & n8863 ;
  assign n13462 = n13460 | n13461 ;
  assign n13463 = x81 & n9125 ;
  assign n13464 = n13462 | n13463 ;
  assign n13465 = ( ~x62 & n13458 ) | ( ~x62 & n13464 ) | ( n13458 & n13464 ) ;
  assign n13466 = x62 & ~n13464 ;
  assign n13467 = ( ~n13459 & n13465 ) | ( ~n13459 & n13466 ) | ( n13465 & n13466 ) ;
  assign n13468 = ( x62 & x63 ) | ( x62 & x80 ) | ( x63 & x80 ) ;
  assign n13469 = ( x62 & x79 ) | ( x62 & ~n9394 ) | ( x79 & ~n9394 ) ;
  assign n13470 = ( x79 & n13468 ) | ( x79 & ~n13469 ) | ( n13468 & ~n13469 ) ;
  assign n13471 = ( n13257 & n13467 ) | ( n13257 & ~n13470 ) | ( n13467 & ~n13470 ) ;
  assign n13472 = ( ~n13257 & n13467 ) | ( ~n13257 & n13470 ) | ( n13467 & n13470 ) ;
  assign n13473 = ( ~n13467 & n13471 ) | ( ~n13467 & n13472 ) | ( n13471 & n13472 ) ;
  assign n13474 = ( n13259 & n13457 ) | ( n13259 & ~n13473 ) | ( n13457 & ~n13473 ) ;
  assign n13475 = ( ~n13259 & n13457 ) | ( ~n13259 & n13473 ) | ( n13457 & n13473 ) ;
  assign n13476 = ( ~n13457 & n13474 ) | ( ~n13457 & n13475 ) | ( n13474 & n13475 ) ;
  assign n13477 = ( n13262 & n13447 ) | ( n13262 & ~n13476 ) | ( n13447 & ~n13476 ) ;
  assign n13478 = ( ~n13262 & n13447 ) | ( ~n13262 & n13476 ) | ( n13447 & n13476 ) ;
  assign n13479 = ( ~n13447 & n13477 ) | ( ~n13447 & n13478 ) | ( n13477 & n13478 ) ;
  assign n13480 = ( n13265 & n13437 ) | ( n13265 & ~n13479 ) | ( n13437 & ~n13479 ) ;
  assign n13481 = ( ~n13265 & n13437 ) | ( ~n13265 & n13479 ) | ( n13437 & n13479 ) ;
  assign n13482 = ( ~n13437 & n13480 ) | ( ~n13437 & n13481 ) | ( n13480 & n13481 ) ;
  assign n13483 = ( n13268 & n13427 ) | ( n13268 & ~n13482 ) | ( n13427 & ~n13482 ) ;
  assign n13484 = ( ~n13268 & n13427 ) | ( ~n13268 & n13482 ) | ( n13427 & n13482 ) ;
  assign n13485 = ( ~n13427 & n13483 ) | ( ~n13427 & n13484 ) | ( n13483 & n13484 ) ;
  assign n13486 = ( n13271 & n13417 ) | ( n13271 & n13485 ) | ( n13417 & n13485 ) ;
  assign n13487 = ( n13271 & ~n13417 ) | ( n13271 & n13485 ) | ( ~n13417 & n13485 ) ;
  assign n13488 = ( n13417 & ~n13486 ) | ( n13417 & n13487 ) | ( ~n13486 & n13487 ) ;
  assign n13489 = ( n13274 & n13407 ) | ( n13274 & n13488 ) | ( n13407 & n13488 ) ;
  assign n13490 = ( n13274 & ~n13407 ) | ( n13274 & n13488 ) | ( ~n13407 & n13488 ) ;
  assign n13491 = ( n13407 & ~n13489 ) | ( n13407 & n13490 ) | ( ~n13489 & n13490 ) ;
  assign n13492 = ( n13277 & n13397 ) | ( n13277 & n13491 ) | ( n13397 & n13491 ) ;
  assign n13493 = ( n13277 & ~n13397 ) | ( n13277 & n13491 ) | ( ~n13397 & n13491 ) ;
  assign n13494 = ( n13397 & ~n13492 ) | ( n13397 & n13493 ) | ( ~n13492 & n13493 ) ;
  assign n13495 = ( n13280 & n13387 ) | ( n13280 & n13494 ) | ( n13387 & n13494 ) ;
  assign n13496 = ( n13280 & ~n13387 ) | ( n13280 & n13494 ) | ( ~n13387 & n13494 ) ;
  assign n13497 = ( n13387 & ~n13495 ) | ( n13387 & n13496 ) | ( ~n13495 & n13496 ) ;
  assign n13498 = ( n13283 & n13377 ) | ( n13283 & n13497 ) | ( n13377 & n13497 ) ;
  assign n13499 = ( ~n13283 & n13377 ) | ( ~n13283 & n13497 ) | ( n13377 & n13497 ) ;
  assign n13500 = ( n13283 & ~n13498 ) | ( n13283 & n13499 ) | ( ~n13498 & n13499 ) ;
  assign n13501 = ( n13286 & n13367 ) | ( n13286 & n13500 ) | ( n13367 & n13500 ) ;
  assign n13502 = ( n13286 & ~n13367 ) | ( n13286 & n13500 ) | ( ~n13367 & n13500 ) ;
  assign n13503 = ( n13367 & ~n13501 ) | ( n13367 & n13502 ) | ( ~n13501 & n13502 ) ;
  assign n13504 = ( n13289 & n13357 ) | ( n13289 & n13503 ) | ( n13357 & n13503 ) ;
  assign n13505 = ( n13289 & ~n13357 ) | ( n13289 & n13503 ) | ( ~n13357 & n13503 ) ;
  assign n13506 = ( n13357 & ~n13504 ) | ( n13357 & n13505 ) | ( ~n13504 & n13505 ) ;
  assign n13507 = ( n13293 & n13347 ) | ( n13293 & n13506 ) | ( n13347 & n13506 ) ;
  assign n13508 = ( n13293 & ~n13347 ) | ( n13293 & n13506 ) | ( ~n13347 & n13506 ) ;
  assign n13509 = ( n13347 & ~n13507 ) | ( n13347 & n13508 ) | ( ~n13507 & n13508 ) ;
  assign n13510 = ( n13295 & n13337 ) | ( n13295 & n13509 ) | ( n13337 & n13509 ) ;
  assign n13511 = ( n13295 & ~n13337 ) | ( n13295 & n13509 ) | ( ~n13337 & n13509 ) ;
  assign n13512 = ( n13337 & ~n13510 ) | ( n13337 & n13511 ) | ( ~n13510 & n13511 ) ;
  assign n13513 = ( n13298 & n13327 ) | ( n13298 & n13512 ) | ( n13327 & n13512 ) ;
  assign n13514 = ( n13298 & ~n13327 ) | ( n13298 & n13512 ) | ( ~n13327 & n13512 ) ;
  assign n13515 = ( n13327 & ~n13513 ) | ( n13327 & n13514 ) | ( ~n13513 & n13514 ) ;
  assign n13516 = ( n13301 & ~n13317 ) | ( n13301 & n13515 ) | ( ~n13317 & n13515 ) ;
  assign n13517 = ( n13301 & n13317 ) | ( n13301 & n13515 ) | ( n13317 & n13515 ) ;
  assign n13518 = ( n13317 & n13516 ) | ( n13317 & ~n13517 ) | ( n13516 & ~n13517 ) ;
  assign n13519 = ( n13304 & n13307 ) | ( n13304 & n13518 ) | ( n13307 & n13518 ) ;
  assign n13520 = ( n13304 & ~n13307 ) | ( n13304 & n13518 ) | ( ~n13307 & n13518 ) ;
  assign n13521 = ( n13307 & ~n13519 ) | ( n13307 & n13520 ) | ( ~n13519 & n13520 ) ;
  assign n13522 = n958 | n9864 ;
  assign n13523 = x127 & ~n878 ;
  assign n13524 = n13522 & n13523 ;
  assign n13525 = x17 | n13524 ;
  assign n13526 = ~x16 & n13524 ;
  assign n13527 = n13525 & ~n13526 ;
  assign n13528 = n1146 & n9038 ;
  assign n13529 = x20 & n13528 ;
  assign n13530 = x126 & n1153 ;
  assign n13531 = x125 & n1150 ;
  assign n13532 = n13530 | n13531 ;
  assign n13533 = x124 & n1217 ;
  assign n13534 = n13532 | n13533 ;
  assign n13535 = ( ~x20 & n13528 ) | ( ~x20 & n13534 ) | ( n13528 & n13534 ) ;
  assign n13536 = x20 & ~n13534 ;
  assign n13537 = ( ~n13529 & n13535 ) | ( ~n13529 & n13536 ) | ( n13535 & n13536 ) ;
  assign n13538 = n1427 & n8461 ;
  assign n13539 = x23 & n13538 ;
  assign n13540 = x123 & n1434 ;
  assign n13541 = x122 & n1431 ;
  assign n13542 = n13540 | n13541 ;
  assign n13543 = x121 & n1531 ;
  assign n13544 = n13542 | n13543 ;
  assign n13545 = ( ~x23 & n13538 ) | ( ~x23 & n13544 ) | ( n13538 & n13544 ) ;
  assign n13546 = x23 & ~n13544 ;
  assign n13547 = ( ~n13539 & n13545 ) | ( ~n13539 & n13546 ) | ( n13545 & n13546 ) ;
  assign n13548 = n1755 & n7444 ;
  assign n13549 = x26 & n13548 ;
  assign n13550 = x120 & n1762 ;
  assign n13551 = x119 & n1759 ;
  assign n13552 = n13550 | n13551 ;
  assign n13553 = x118 & n1895 ;
  assign n13554 = n13552 | n13553 ;
  assign n13555 = ( ~x26 & n13548 ) | ( ~x26 & n13554 ) | ( n13548 & n13554 ) ;
  assign n13556 = x26 & ~n13554 ;
  assign n13557 = ( ~n13549 & n13555 ) | ( ~n13549 & n13556 ) | ( n13555 & n13556 ) ;
  assign n13558 = n2137 & n6924 ;
  assign n13559 = x29 & n13558 ;
  assign n13560 = x117 & n2144 ;
  assign n13561 = x116 & n2141 ;
  assign n13562 = n13560 | n13561 ;
  assign n13563 = x115 & n2267 ;
  assign n13564 = n13562 | n13563 ;
  assign n13565 = ( ~x29 & n13558 ) | ( ~x29 & n13564 ) | ( n13558 & n13564 ) ;
  assign n13566 = x29 & ~n13564 ;
  assign n13567 = ( ~n13559 & n13565 ) | ( ~n13559 & n13566 ) | ( n13565 & n13566 ) ;
  assign n13568 = n2545 & n6002 ;
  assign n13569 = x32 & n13568 ;
  assign n13570 = x114 & n2552 ;
  assign n13571 = x113 & n2549 ;
  assign n13572 = n13570 | n13571 ;
  assign n13573 = x112 & n2696 ;
  assign n13574 = n13572 | n13573 ;
  assign n13575 = ( ~x32 & n13568 ) | ( ~x32 & n13574 ) | ( n13568 & n13574 ) ;
  assign n13576 = x32 & ~n13574 ;
  assign n13577 = ( ~n13569 & n13575 ) | ( ~n13569 & n13576 ) | ( n13575 & n13576 ) ;
  assign n13578 = n2982 & n5347 ;
  assign n13579 = x35 & n13578 ;
  assign n13580 = x111 & n2989 ;
  assign n13581 = x110 & n2986 ;
  assign n13582 = n13580 | n13581 ;
  assign n13583 = x109 & n3159 ;
  assign n13584 = n13582 | n13583 ;
  assign n13585 = ( ~x35 & n13578 ) | ( ~x35 & n13584 ) | ( n13578 & n13584 ) ;
  assign n13586 = x35 & ~n13584 ;
  assign n13587 = ( ~n13579 & n13585 ) | ( ~n13579 & n13586 ) | ( n13585 & n13586 ) ;
  assign n13588 = n3492 & n4914 ;
  assign n13589 = x38 & n13588 ;
  assign n13590 = x108 & n3499 ;
  assign n13591 = x107 & n3496 ;
  assign n13592 = n13590 | n13591 ;
  assign n13593 = x106 & n3662 ;
  assign n13594 = n13592 | n13593 ;
  assign n13595 = ( ~x38 & n13588 ) | ( ~x38 & n13594 ) | ( n13588 & n13594 ) ;
  assign n13596 = x38 & ~n13594 ;
  assign n13597 = ( ~n13589 & n13595 ) | ( ~n13589 & n13596 ) | ( n13595 & n13596 ) ;
  assign n13598 = n4020 & n4145 ;
  assign n13599 = x41 & n13598 ;
  assign n13600 = x105 & n4027 ;
  assign n13601 = x104 & n4024 ;
  assign n13602 = n13600 | n13601 ;
  assign n13603 = x103 & n4223 ;
  assign n13604 = n13602 | n13603 ;
  assign n13605 = ( ~x41 & n13598 ) | ( ~x41 & n13604 ) | ( n13598 & n13604 ) ;
  assign n13606 = x41 & ~n13604 ;
  assign n13607 = ( ~n13599 & n13605 ) | ( ~n13599 & n13606 ) | ( n13605 & n13606 ) ;
  assign n13608 = n3764 & n4625 ;
  assign n13609 = x44 & n13608 ;
  assign n13610 = x102 & n4791 ;
  assign n13611 = x101 & n4621 ;
  assign n13612 = n13610 | n13611 ;
  assign n13613 = x100 & n4795 ;
  assign n13614 = n13612 | n13613 ;
  assign n13615 = ( ~x44 & n13608 ) | ( ~x44 & n13614 ) | ( n13608 & n13614 ) ;
  assign n13616 = x44 & ~n13614 ;
  assign n13617 = ( ~n13609 & n13615 ) | ( ~n13609 & n13616 ) | ( n13615 & n13616 ) ;
  assign n13618 = n3248 & n5223 ;
  assign n13619 = x47 & n13618 ;
  assign n13620 = x99 & n5230 ;
  assign n13621 = x98 & n5227 ;
  assign n13622 = n13620 | n13621 ;
  assign n13623 = x97 & n5434 ;
  assign n13624 = n13622 | n13623 ;
  assign n13625 = ( ~x47 & n13618 ) | ( ~x47 & n13624 ) | ( n13618 & n13624 ) ;
  assign n13626 = x47 & ~n13624 ;
  assign n13627 = ( ~n13619 & n13625 ) | ( ~n13619 & n13626 ) | ( n13625 & n13626 ) ;
  assign n13628 = n2772 & n5858 ;
  assign n13629 = x50 & n13628 ;
  assign n13630 = x96 & n5865 ;
  assign n13631 = x95 & n5862 ;
  assign n13632 = n13630 | n13631 ;
  assign n13633 = x94 & n6092 ;
  assign n13634 = n13632 | n13633 ;
  assign n13635 = ( ~x50 & n13628 ) | ( ~x50 & n13634 ) | ( n13628 & n13634 ) ;
  assign n13636 = x50 & ~n13634 ;
  assign n13637 = ( ~n13629 & n13635 ) | ( ~n13629 & n13636 ) | ( n13635 & n13636 ) ;
  assign n13638 = n2220 & n6546 ;
  assign n13639 = x53 & n13638 ;
  assign n13640 = x93 & n6553 ;
  assign n13641 = x92 & n6550 ;
  assign n13642 = n13640 | n13641 ;
  assign n13643 = x91 & n6787 ;
  assign n13644 = n13642 | n13643 ;
  assign n13645 = ( ~x53 & n13638 ) | ( ~x53 & n13644 ) | ( n13638 & n13644 ) ;
  assign n13646 = x53 & ~n13644 ;
  assign n13647 = ( ~n13639 & n13645 ) | ( ~n13639 & n13646 ) | ( n13645 & n13646 ) ;
  assign n13648 = n1838 & n7277 ;
  assign n13649 = x56 & n13648 ;
  assign n13650 = x90 & n7545 ;
  assign n13651 = x89 & n7273 ;
  assign n13652 = n13650 | n13651 ;
  assign n13653 = x88 & n7552 ;
  assign n13654 = n13652 | n13653 ;
  assign n13655 = ( ~x56 & n13648 ) | ( ~x56 & n13654 ) | ( n13648 & n13654 ) ;
  assign n13656 = x56 & ~n13654 ;
  assign n13657 = ( ~n13649 & n13655 ) | ( ~n13649 & n13656 ) | ( n13655 & n13656 ) ;
  assign n13658 = n1494 & n8067 ;
  assign n13659 = x59 & n13658 ;
  assign n13660 = x87 & n8074 ;
  assign n13661 = x86 & n8071 ;
  assign n13662 = n13660 | n13661 ;
  assign n13663 = x85 & n8298 ;
  assign n13664 = n13662 | n13663 ;
  assign n13665 = ( ~x59 & n13658 ) | ( ~x59 & n13664 ) | ( n13658 & n13664 ) ;
  assign n13666 = x59 & ~n13664 ;
  assign n13667 = ( ~n13659 & n13665 ) | ( ~n13659 & n13666 ) | ( n13665 & n13666 ) ;
  assign n13668 = ( x62 & x63 ) | ( x62 & x81 ) | ( x63 & x81 ) ;
  assign n13669 = ( x62 & x80 ) | ( x62 & ~n9394 ) | ( x80 & ~n9394 ) ;
  assign n13670 = ( x80 & n13668 ) | ( x80 & ~n13669 ) | ( n13668 & ~n13669 ) ;
  assign n13671 = n1190 & n8859 ;
  assign n13672 = x62 & n13671 ;
  assign n13673 = x84 & n8866 ;
  assign n13674 = x83 & n8863 ;
  assign n13675 = n13673 | n13674 ;
  assign n13676 = x82 & n9125 ;
  assign n13677 = n13675 | n13676 ;
  assign n13678 = ( ~x62 & n13671 ) | ( ~x62 & n13677 ) | ( n13671 & n13677 ) ;
  assign n13679 = x62 & ~n13677 ;
  assign n13680 = ( ~n13672 & n13678 ) | ( ~n13672 & n13679 ) | ( n13678 & n13679 ) ;
  assign n13681 = ( n13470 & n13670 ) | ( n13470 & n13680 ) | ( n13670 & n13680 ) ;
  assign n13682 = ( n13470 & ~n13670 ) | ( n13470 & n13680 ) | ( ~n13670 & n13680 ) ;
  assign n13683 = ( n13670 & ~n13681 ) | ( n13670 & n13682 ) | ( ~n13681 & n13682 ) ;
  assign n13684 = ( n13471 & ~n13667 ) | ( n13471 & n13683 ) | ( ~n13667 & n13683 ) ;
  assign n13685 = ( n13471 & n13667 ) | ( n13471 & ~n13683 ) | ( n13667 & ~n13683 ) ;
  assign n13686 = ( ~n13471 & n13684 ) | ( ~n13471 & n13685 ) | ( n13684 & n13685 ) ;
  assign n13687 = ( n13474 & n13657 ) | ( n13474 & ~n13686 ) | ( n13657 & ~n13686 ) ;
  assign n13688 = ( ~n13474 & n13657 ) | ( ~n13474 & n13686 ) | ( n13657 & n13686 ) ;
  assign n13689 = ( ~n13657 & n13687 ) | ( ~n13657 & n13688 ) | ( n13687 & n13688 ) ;
  assign n13690 = ( n13477 & n13647 ) | ( n13477 & ~n13689 ) | ( n13647 & ~n13689 ) ;
  assign n13691 = ( ~n13477 & n13647 ) | ( ~n13477 & n13689 ) | ( n13647 & n13689 ) ;
  assign n13692 = ( ~n13647 & n13690 ) | ( ~n13647 & n13691 ) | ( n13690 & n13691 ) ;
  assign n13693 = ( n13480 & n13637 ) | ( n13480 & ~n13692 ) | ( n13637 & ~n13692 ) ;
  assign n13694 = ( ~n13480 & n13637 ) | ( ~n13480 & n13692 ) | ( n13637 & n13692 ) ;
  assign n13695 = ( ~n13637 & n13693 ) | ( ~n13637 & n13694 ) | ( n13693 & n13694 ) ;
  assign n13696 = ( n13483 & n13627 ) | ( n13483 & ~n13695 ) | ( n13627 & ~n13695 ) ;
  assign n13697 = ( ~n13483 & n13627 ) | ( ~n13483 & n13695 ) | ( n13627 & n13695 ) ;
  assign n13698 = ( ~n13627 & n13696 ) | ( ~n13627 & n13697 ) | ( n13696 & n13697 ) ;
  assign n13699 = ( n13487 & n13617 ) | ( n13487 & n13698 ) | ( n13617 & n13698 ) ;
  assign n13700 = ( n13487 & ~n13617 ) | ( n13487 & n13698 ) | ( ~n13617 & n13698 ) ;
  assign n13701 = ( n13617 & ~n13699 ) | ( n13617 & n13700 ) | ( ~n13699 & n13700 ) ;
  assign n13702 = ( n13489 & n13607 ) | ( n13489 & n13701 ) | ( n13607 & n13701 ) ;
  assign n13703 = ( n13489 & ~n13607 ) | ( n13489 & n13701 ) | ( ~n13607 & n13701 ) ;
  assign n13704 = ( n13607 & ~n13702 ) | ( n13607 & n13703 ) | ( ~n13702 & n13703 ) ;
  assign n13705 = ( n13492 & n13597 ) | ( n13492 & n13704 ) | ( n13597 & n13704 ) ;
  assign n13706 = ( n13492 & ~n13597 ) | ( n13492 & n13704 ) | ( ~n13597 & n13704 ) ;
  assign n13707 = ( n13597 & ~n13705 ) | ( n13597 & n13706 ) | ( ~n13705 & n13706 ) ;
  assign n13708 = ( n13495 & n13587 ) | ( n13495 & n13707 ) | ( n13587 & n13707 ) ;
  assign n13709 = ( n13495 & ~n13587 ) | ( n13495 & n13707 ) | ( ~n13587 & n13707 ) ;
  assign n13710 = ( n13587 & ~n13708 ) | ( n13587 & n13709 ) | ( ~n13708 & n13709 ) ;
  assign n13711 = ( n13498 & n13577 ) | ( n13498 & n13710 ) | ( n13577 & n13710 ) ;
  assign n13712 = ( n13498 & ~n13577 ) | ( n13498 & n13710 ) | ( ~n13577 & n13710 ) ;
  assign n13713 = ( n13577 & ~n13711 ) | ( n13577 & n13712 ) | ( ~n13711 & n13712 ) ;
  assign n13714 = ( n13501 & n13567 ) | ( n13501 & n13713 ) | ( n13567 & n13713 ) ;
  assign n13715 = ( n13501 & ~n13567 ) | ( n13501 & n13713 ) | ( ~n13567 & n13713 ) ;
  assign n13716 = ( n13567 & ~n13714 ) | ( n13567 & n13715 ) | ( ~n13714 & n13715 ) ;
  assign n13717 = ( n13504 & n13557 ) | ( n13504 & n13716 ) | ( n13557 & n13716 ) ;
  assign n13718 = ( n13504 & ~n13557 ) | ( n13504 & n13716 ) | ( ~n13557 & n13716 ) ;
  assign n13719 = ( n13557 & ~n13717 ) | ( n13557 & n13718 ) | ( ~n13717 & n13718 ) ;
  assign n13720 = ( n13507 & n13547 ) | ( n13507 & n13719 ) | ( n13547 & n13719 ) ;
  assign n13721 = ( n13507 & ~n13547 ) | ( n13507 & n13719 ) | ( ~n13547 & n13719 ) ;
  assign n13722 = ( n13547 & ~n13720 ) | ( n13547 & n13721 ) | ( ~n13720 & n13721 ) ;
  assign n13723 = ( n13510 & n13537 ) | ( n13510 & n13722 ) | ( n13537 & n13722 ) ;
  assign n13724 = ( n13510 & ~n13537 ) | ( n13510 & n13722 ) | ( ~n13537 & n13722 ) ;
  assign n13725 = ( n13537 & ~n13723 ) | ( n13537 & n13724 ) | ( ~n13723 & n13724 ) ;
  assign n13726 = ( n13513 & ~n13527 ) | ( n13513 & n13725 ) | ( ~n13527 & n13725 ) ;
  assign n13727 = ( n13513 & n13527 ) | ( n13513 & n13725 ) | ( n13527 & n13725 ) ;
  assign n13728 = ( n13527 & n13726 ) | ( n13527 & ~n13727 ) | ( n13726 & ~n13727 ) ;
  assign n13729 = ( n13517 & n13519 ) | ( n13517 & n13728 ) | ( n13519 & n13728 ) ;
  assign n13730 = ( n13517 & ~n13519 ) | ( n13517 & n13728 ) | ( ~n13519 & n13728 ) ;
  assign n13731 = ( n13519 & ~n13729 ) | ( n13519 & n13730 ) | ( ~n13729 & n13730 ) ;
  assign n13732 = n1146 & n9576 ;
  assign n13733 = x20 & n13732 ;
  assign n13734 = x127 & n1153 ;
  assign n13735 = x126 & n1150 ;
  assign n13736 = n13734 | n13735 ;
  assign n13737 = x125 & n1217 ;
  assign n13738 = n13736 | n13737 ;
  assign n13739 = ( ~x20 & n13732 ) | ( ~x20 & n13738 ) | ( n13732 & n13738 ) ;
  assign n13740 = x20 & ~n13738 ;
  assign n13741 = ( ~n13733 & n13739 ) | ( ~n13733 & n13740 ) | ( n13739 & n13740 ) ;
  assign n13742 = n1427 & n8729 ;
  assign n13743 = x23 & n13742 ;
  assign n13744 = x124 & n1434 ;
  assign n13745 = x123 & n1431 ;
  assign n13746 = n13744 | n13745 ;
  assign n13747 = x122 & n1531 ;
  assign n13748 = n13746 | n13747 ;
  assign n13749 = ( ~x23 & n13742 ) | ( ~x23 & n13748 ) | ( n13742 & n13748 ) ;
  assign n13750 = x23 & ~n13748 ;
  assign n13751 = ( ~n13743 & n13749 ) | ( ~n13743 & n13750 ) | ( n13749 & n13750 ) ;
  assign n13752 = n1755 & n7696 ;
  assign n13753 = x26 & n13752 ;
  assign n13754 = x121 & n1762 ;
  assign n13755 = x120 & n1759 ;
  assign n13756 = n13754 | n13755 ;
  assign n13757 = x119 & n1895 ;
  assign n13758 = n13756 | n13757 ;
  assign n13759 = ( ~x26 & n13752 ) | ( ~x26 & n13758 ) | ( n13752 & n13758 ) ;
  assign n13760 = x26 & ~n13758 ;
  assign n13761 = ( ~n13753 & n13759 ) | ( ~n13753 & n13760 ) | ( n13759 & n13760 ) ;
  assign n13762 = n2137 & n6940 ;
  assign n13763 = x29 & n13762 ;
  assign n13764 = x118 & n2144 ;
  assign n13765 = x117 & n2141 ;
  assign n13766 = n13764 | n13765 ;
  assign n13767 = x116 & n2267 ;
  assign n13768 = n13766 | n13767 ;
  assign n13769 = ( ~x29 & n13762 ) | ( ~x29 & n13768 ) | ( n13762 & n13768 ) ;
  assign n13770 = x29 & ~n13768 ;
  assign n13771 = ( ~n13763 & n13769 ) | ( ~n13763 & n13770 ) | ( n13769 & n13770 ) ;
  assign n13772 = n2545 & n6446 ;
  assign n13773 = x32 & n13772 ;
  assign n13774 = x115 & n2552 ;
  assign n13775 = x114 & n2549 ;
  assign n13776 = n13774 | n13775 ;
  assign n13777 = x113 & n2696 ;
  assign n13778 = n13776 | n13777 ;
  assign n13779 = ( ~x32 & n13772 ) | ( ~x32 & n13778 ) | ( n13772 & n13778 ) ;
  assign n13780 = x32 & ~n13778 ;
  assign n13781 = ( ~n13773 & n13779 ) | ( ~n13773 & n13780 ) | ( n13779 & n13780 ) ;
  assign n13782 = n2982 & n5558 ;
  assign n13783 = x35 & n13782 ;
  assign n13784 = x112 & n2989 ;
  assign n13785 = x111 & n2986 ;
  assign n13786 = n13784 | n13785 ;
  assign n13787 = x110 & n3159 ;
  assign n13788 = n13786 | n13787 ;
  assign n13789 = ( ~x35 & n13782 ) | ( ~x35 & n13788 ) | ( n13782 & n13788 ) ;
  assign n13790 = x35 & ~n13788 ;
  assign n13791 = ( ~n13783 & n13789 ) | ( ~n13783 & n13790 ) | ( n13789 & n13790 ) ;
  assign n13792 = n3492 & n4930 ;
  assign n13793 = x38 & n13792 ;
  assign n13794 = x109 & n3499 ;
  assign n13795 = x108 & n3496 ;
  assign n13796 = n13794 | n13795 ;
  assign n13797 = x107 & n3662 ;
  assign n13798 = n13796 | n13797 ;
  assign n13799 = ( ~x38 & n13792 ) | ( ~x38 & n13798 ) | ( n13792 & n13798 ) ;
  assign n13800 = x38 & ~n13798 ;
  assign n13801 = ( ~n13793 & n13799 ) | ( ~n13793 & n13800 ) | ( n13799 & n13800 ) ;
  assign n13802 = n4020 & n4331 ;
  assign n13803 = x41 & n13802 ;
  assign n13804 = x106 & n4027 ;
  assign n13805 = x105 & n4024 ;
  assign n13806 = n13804 | n13805 ;
  assign n13807 = x104 & n4223 ;
  assign n13808 = n13806 | n13807 ;
  assign n13809 = ( ~x41 & n13802 ) | ( ~x41 & n13808 ) | ( n13802 & n13808 ) ;
  assign n13810 = x41 & ~n13808 ;
  assign n13811 = ( ~n13803 & n13809 ) | ( ~n13803 & n13810 ) | ( n13809 & n13810 ) ;
  assign n13812 = n3941 & n4625 ;
  assign n13813 = x44 & n13812 ;
  assign n13814 = x103 & n4791 ;
  assign n13815 = x102 & n4621 ;
  assign n13816 = n13814 | n13815 ;
  assign n13817 = x101 & n4795 ;
  assign n13818 = n13816 | n13817 ;
  assign n13819 = ( ~x44 & n13812 ) | ( ~x44 & n13818 ) | ( n13812 & n13818 ) ;
  assign n13820 = x44 & ~n13818 ;
  assign n13821 = ( ~n13813 & n13819 ) | ( ~n13813 & n13820 ) | ( n13819 & n13820 ) ;
  assign n13822 = n3264 & n5223 ;
  assign n13823 = x47 & n13822 ;
  assign n13824 = x100 & n5230 ;
  assign n13825 = x99 & n5227 ;
  assign n13826 = n13824 | n13825 ;
  assign n13827 = x98 & n5434 ;
  assign n13828 = n13826 | n13827 ;
  assign n13829 = ( ~x47 & n13822 ) | ( ~x47 & n13828 ) | ( n13822 & n13828 ) ;
  assign n13830 = x47 & ~n13828 ;
  assign n13831 = ( ~n13823 & n13829 ) | ( ~n13823 & n13830 ) | ( n13829 & n13830 ) ;
  assign n13832 = n2788 & n5858 ;
  assign n13833 = x50 & n13832 ;
  assign n13834 = x97 & n5865 ;
  assign n13835 = x96 & n5862 ;
  assign n13836 = n13834 | n13835 ;
  assign n13837 = x95 & n6092 ;
  assign n13838 = n13836 | n13837 ;
  assign n13839 = ( ~x50 & n13832 ) | ( ~x50 & n13838 ) | ( n13832 & n13838 ) ;
  assign n13840 = x50 & ~n13838 ;
  assign n13841 = ( ~n13833 & n13839 ) | ( ~n13833 & n13840 ) | ( n13839 & n13840 ) ;
  assign n13842 = n2476 & n6546 ;
  assign n13843 = x53 & n13842 ;
  assign n13844 = x94 & n6553 ;
  assign n13845 = x93 & n6550 ;
  assign n13846 = n13844 | n13845 ;
  assign n13847 = x92 & n6787 ;
  assign n13848 = n13846 | n13847 ;
  assign n13849 = ( ~x53 & n13842 ) | ( ~x53 & n13848 ) | ( n13842 & n13848 ) ;
  assign n13850 = x53 & ~n13848 ;
  assign n13851 = ( ~n13843 & n13849 ) | ( ~n13843 & n13850 ) | ( n13849 & n13850 ) ;
  assign n13852 = n1959 & n7277 ;
  assign n13853 = x56 & n13852 ;
  assign n13854 = x91 & n7545 ;
  assign n13855 = x90 & n7273 ;
  assign n13856 = n13854 | n13855 ;
  assign n13857 = x89 & n7552 ;
  assign n13858 = n13856 | n13857 ;
  assign n13859 = ( ~x56 & n13852 ) | ( ~x56 & n13858 ) | ( n13852 & n13858 ) ;
  assign n13860 = x56 & ~n13858 ;
  assign n13861 = ( ~n13853 & n13859 ) | ( ~n13853 & n13860 ) | ( n13859 & n13860 ) ;
  assign n13862 = n1602 & n8067 ;
  assign n13863 = x59 & n13862 ;
  assign n13864 = x88 & n8074 ;
  assign n13865 = x87 & n8071 ;
  assign n13866 = n13864 | n13865 ;
  assign n13867 = x86 & n8298 ;
  assign n13868 = n13866 | n13867 ;
  assign n13869 = ( ~x59 & n13862 ) | ( ~x59 & n13868 ) | ( n13862 & n13868 ) ;
  assign n13870 = x59 & ~n13868 ;
  assign n13871 = ( ~n13863 & n13869 ) | ( ~n13863 & n13870 ) | ( n13869 & n13870 ) ;
  assign n13872 = n1368 & n8859 ;
  assign n13873 = x62 & n13872 ;
  assign n13874 = x85 & n8866 ;
  assign n13875 = x84 & n8863 ;
  assign n13876 = n13874 | n13875 ;
  assign n13877 = x83 & n9125 ;
  assign n13878 = n13876 | n13877 ;
  assign n13879 = ( ~x62 & n13872 ) | ( ~x62 & n13878 ) | ( n13872 & n13878 ) ;
  assign n13880 = x62 & ~n13878 ;
  assign n13881 = ( ~n13873 & n13879 ) | ( ~n13873 & n13880 ) | ( n13879 & n13880 ) ;
  assign n13882 = ( x62 & x63 ) | ( x62 & x82 ) | ( x63 & x82 ) ;
  assign n13883 = ( x62 & x81 ) | ( x62 & ~n9394 ) | ( x81 & ~n9394 ) ;
  assign n13884 = ( x81 & n13882 ) | ( x81 & ~n13883 ) | ( n13882 & ~n13883 ) ;
  assign n13885 = ( x17 & n13670 ) | ( x17 & n13884 ) | ( n13670 & n13884 ) ;
  assign n13886 = ( ~x17 & n13670 ) | ( ~x17 & n13884 ) | ( n13670 & n13884 ) ;
  assign n13887 = ( x17 & ~n13885 ) | ( x17 & n13886 ) | ( ~n13885 & n13886 ) ;
  assign n13888 = ( n13682 & n13881 ) | ( n13682 & ~n13887 ) | ( n13881 & ~n13887 ) ;
  assign n13889 = ( ~n13682 & n13881 ) | ( ~n13682 & n13887 ) | ( n13881 & n13887 ) ;
  assign n13890 = ( ~n13881 & n13888 ) | ( ~n13881 & n13889 ) | ( n13888 & n13889 ) ;
  assign n13891 = ( n13685 & n13871 ) | ( n13685 & ~n13890 ) | ( n13871 & ~n13890 ) ;
  assign n13892 = ( n13685 & ~n13871 ) | ( n13685 & n13890 ) | ( ~n13871 & n13890 ) ;
  assign n13893 = ( ~n13685 & n13891 ) | ( ~n13685 & n13892 ) | ( n13891 & n13892 ) ;
  assign n13894 = ( n13687 & n13861 ) | ( n13687 & ~n13893 ) | ( n13861 & ~n13893 ) ;
  assign n13895 = ( n13687 & ~n13861 ) | ( n13687 & n13893 ) | ( ~n13861 & n13893 ) ;
  assign n13896 = ( ~n13687 & n13894 ) | ( ~n13687 & n13895 ) | ( n13894 & n13895 ) ;
  assign n13897 = ( n13690 & n13851 ) | ( n13690 & ~n13896 ) | ( n13851 & ~n13896 ) ;
  assign n13898 = ( n13690 & ~n13851 ) | ( n13690 & n13896 ) | ( ~n13851 & n13896 ) ;
  assign n13899 = ( ~n13690 & n13897 ) | ( ~n13690 & n13898 ) | ( n13897 & n13898 ) ;
  assign n13900 = ( n13693 & n13841 ) | ( n13693 & ~n13899 ) | ( n13841 & ~n13899 ) ;
  assign n13901 = ( n13693 & ~n13841 ) | ( n13693 & n13899 ) | ( ~n13841 & n13899 ) ;
  assign n13902 = ( ~n13693 & n13900 ) | ( ~n13693 & n13901 ) | ( n13900 & n13901 ) ;
  assign n13903 = ( n13696 & n13831 ) | ( n13696 & ~n13902 ) | ( n13831 & ~n13902 ) ;
  assign n13904 = ( n13696 & ~n13831 ) | ( n13696 & n13902 ) | ( ~n13831 & n13902 ) ;
  assign n13905 = ( ~n13696 & n13903 ) | ( ~n13696 & n13904 ) | ( n13903 & n13904 ) ;
  assign n13906 = ( n13700 & ~n13821 ) | ( n13700 & n13905 ) | ( ~n13821 & n13905 ) ;
  assign n13907 = ( n13700 & n13821 ) | ( n13700 & ~n13905 ) | ( n13821 & ~n13905 ) ;
  assign n13908 = ( ~n13700 & n13906 ) | ( ~n13700 & n13907 ) | ( n13906 & n13907 ) ;
  assign n13909 = ( n13702 & n13811 ) | ( n13702 & n13908 ) | ( n13811 & n13908 ) ;
  assign n13910 = ( ~n13702 & n13811 ) | ( ~n13702 & n13908 ) | ( n13811 & n13908 ) ;
  assign n13911 = ( n13702 & ~n13909 ) | ( n13702 & n13910 ) | ( ~n13909 & n13910 ) ;
  assign n13912 = ( n13705 & n13801 ) | ( n13705 & n13911 ) | ( n13801 & n13911 ) ;
  assign n13913 = ( ~n13705 & n13801 ) | ( ~n13705 & n13911 ) | ( n13801 & n13911 ) ;
  assign n13914 = ( n13705 & ~n13912 ) | ( n13705 & n13913 ) | ( ~n13912 & n13913 ) ;
  assign n13915 = ( n13708 & n13791 ) | ( n13708 & n13914 ) | ( n13791 & n13914 ) ;
  assign n13916 = ( ~n13708 & n13791 ) | ( ~n13708 & n13914 ) | ( n13791 & n13914 ) ;
  assign n13917 = ( n13708 & ~n13915 ) | ( n13708 & n13916 ) | ( ~n13915 & n13916 ) ;
  assign n13918 = ( n13711 & n13781 ) | ( n13711 & n13917 ) | ( n13781 & n13917 ) ;
  assign n13919 = ( ~n13711 & n13781 ) | ( ~n13711 & n13917 ) | ( n13781 & n13917 ) ;
  assign n13920 = ( n13711 & ~n13918 ) | ( n13711 & n13919 ) | ( ~n13918 & n13919 ) ;
  assign n13921 = ( n13714 & n13771 ) | ( n13714 & n13920 ) | ( n13771 & n13920 ) ;
  assign n13922 = ( ~n13714 & n13771 ) | ( ~n13714 & n13920 ) | ( n13771 & n13920 ) ;
  assign n13923 = ( n13714 & ~n13921 ) | ( n13714 & n13922 ) | ( ~n13921 & n13922 ) ;
  assign n13924 = ( n13717 & n13761 ) | ( n13717 & n13923 ) | ( n13761 & n13923 ) ;
  assign n13925 = ( n13717 & ~n13761 ) | ( n13717 & n13923 ) | ( ~n13761 & n13923 ) ;
  assign n13926 = ( n13761 & ~n13924 ) | ( n13761 & n13925 ) | ( ~n13924 & n13925 ) ;
  assign n13927 = ( n13720 & n13751 ) | ( n13720 & n13926 ) | ( n13751 & n13926 ) ;
  assign n13928 = ( ~n13720 & n13751 ) | ( ~n13720 & n13926 ) | ( n13751 & n13926 ) ;
  assign n13929 = ( n13720 & ~n13927 ) | ( n13720 & n13928 ) | ( ~n13927 & n13928 ) ;
  assign n13930 = ( ~n13723 & n13741 ) | ( ~n13723 & n13929 ) | ( n13741 & n13929 ) ;
  assign n13931 = ( n13723 & n13741 ) | ( n13723 & n13929 ) | ( n13741 & n13929 ) ;
  assign n13932 = ( n13723 & n13930 ) | ( n13723 & ~n13931 ) | ( n13930 & ~n13931 ) ;
  assign n13933 = ( n13727 & n13729 ) | ( n13727 & n13932 ) | ( n13729 & n13932 ) ;
  assign n13934 = ( n13727 & ~n13729 ) | ( n13727 & n13932 ) | ( ~n13729 & n13932 ) ;
  assign n13935 = ( n13729 & ~n13933 ) | ( n13729 & n13934 ) | ( ~n13933 & n13934 ) ;
  assign n13936 = x126 & n1217 ;
  assign n13937 = x20 & n13936 ;
  assign n13938 = x127 & n1150 ;
  assign n13939 = n1146 | n13938 ;
  assign n13940 = ( n9867 & n13938 ) | ( n9867 & n13939 ) | ( n13938 & n13939 ) ;
  assign n13941 = ( ~x20 & n13936 ) | ( ~x20 & n13940 ) | ( n13936 & n13940 ) ;
  assign n13942 = x20 & ~n13940 ;
  assign n13943 = ( ~n13937 & n13941 ) | ( ~n13937 & n13942 ) | ( n13941 & n13942 ) ;
  assign n13944 = n1427 & n9009 ;
  assign n13945 = x23 & n13944 ;
  assign n13946 = x125 & n1434 ;
  assign n13947 = x124 & n1431 ;
  assign n13948 = n13946 | n13947 ;
  assign n13949 = x123 & n1531 ;
  assign n13950 = n13948 | n13949 ;
  assign n13951 = ( ~x23 & n13944 ) | ( ~x23 & n13950 ) | ( n13944 & n13950 ) ;
  assign n13952 = x23 & ~n13950 ;
  assign n13953 = ( ~n13945 & n13951 ) | ( ~n13945 & n13952 ) | ( n13951 & n13952 ) ;
  assign n13954 = n1755 & n8207 ;
  assign n13955 = x26 & n13954 ;
  assign n13956 = x122 & n1762 ;
  assign n13957 = x121 & n1759 ;
  assign n13958 = n13956 | n13957 ;
  assign n13959 = x120 & n1895 ;
  assign n13960 = n13958 | n13959 ;
  assign n13961 = ( ~x26 & n13954 ) | ( ~x26 & n13960 ) | ( n13954 & n13960 ) ;
  assign n13962 = x26 & ~n13960 ;
  assign n13963 = ( ~n13955 & n13961 ) | ( ~n13955 & n13962 ) | ( n13961 & n13962 ) ;
  assign n13964 = n2137 & n7181 ;
  assign n13965 = x29 & n13964 ;
  assign n13966 = x119 & n2144 ;
  assign n13967 = x118 & n2141 ;
  assign n13968 = n13966 | n13967 ;
  assign n13969 = x117 & n2267 ;
  assign n13970 = n13968 | n13969 ;
  assign n13971 = ( ~x29 & n13964 ) | ( ~x29 & n13970 ) | ( n13964 & n13970 ) ;
  assign n13972 = x29 & ~n13970 ;
  assign n13973 = ( ~n13965 & n13971 ) | ( ~n13965 & n13972 ) | ( n13971 & n13972 ) ;
  assign n13974 = n2545 & n6462 ;
  assign n13975 = x32 & n13974 ;
  assign n13976 = x116 & n2552 ;
  assign n13977 = x115 & n2549 ;
  assign n13978 = n13976 | n13977 ;
  assign n13979 = x114 & n2696 ;
  assign n13980 = n13978 | n13979 ;
  assign n13981 = ( ~x32 & n13974 ) | ( ~x32 & n13980 ) | ( n13974 & n13980 ) ;
  assign n13982 = x32 & ~n13980 ;
  assign n13983 = ( ~n13975 & n13981 ) | ( ~n13975 & n13982 ) | ( n13981 & n13982 ) ;
  assign n13984 = n2982 & n5774 ;
  assign n13985 = x35 & n13984 ;
  assign n13986 = x113 & n2989 ;
  assign n13987 = x112 & n2986 ;
  assign n13988 = n13986 | n13987 ;
  assign n13989 = x111 & n3159 ;
  assign n13990 = n13988 | n13989 ;
  assign n13991 = ( ~x35 & n13984 ) | ( ~x35 & n13990 ) | ( n13984 & n13990 ) ;
  assign n13992 = x35 & ~n13990 ;
  assign n13993 = ( ~n13985 & n13991 ) | ( ~n13985 & n13992 ) | ( n13991 & n13992 ) ;
  assign n13994 = n3492 & n5331 ;
  assign n13995 = x38 & n13994 ;
  assign n13996 = x110 & n3499 ;
  assign n13997 = x109 & n3496 ;
  assign n13998 = n13996 | n13997 ;
  assign n13999 = x108 & n3662 ;
  assign n14000 = n13998 | n13999 ;
  assign n14001 = ( ~x38 & n13994 ) | ( ~x38 & n14000 ) | ( n13994 & n14000 ) ;
  assign n14002 = x38 & ~n14000 ;
  assign n14003 = ( ~n13995 & n14001 ) | ( ~n13995 & n14002 ) | ( n14001 & n14002 ) ;
  assign n14004 = n4020 & n4523 ;
  assign n14005 = x41 & n14004 ;
  assign n14006 = x107 & n4027 ;
  assign n14007 = x106 & n4024 ;
  assign n14008 = n14006 | n14007 ;
  assign n14009 = x105 & n4223 ;
  assign n14010 = n14008 | n14009 ;
  assign n14011 = ( ~x41 & n14004 ) | ( ~x41 & n14010 ) | ( n14004 & n14010 ) ;
  assign n14012 = x41 & ~n14010 ;
  assign n14013 = ( ~n14005 & n14011 ) | ( ~n14005 & n14012 ) | ( n14011 & n14012 ) ;
  assign n14014 = n3957 & n4625 ;
  assign n14015 = x44 & n14014 ;
  assign n14016 = x104 & n4791 ;
  assign n14017 = x103 & n4621 ;
  assign n14018 = n14016 | n14017 ;
  assign n14019 = x102 & n4795 ;
  assign n14020 = n14018 | n14019 ;
  assign n14021 = ( ~x44 & n14014 ) | ( ~x44 & n14020 ) | ( n14014 & n14020 ) ;
  assign n14022 = x44 & ~n14020 ;
  assign n14023 = ( ~n14015 & n14021 ) | ( ~n14015 & n14022 ) | ( n14021 & n14022 ) ;
  assign n14024 = n3591 & n5223 ;
  assign n14025 = x47 & n14024 ;
  assign n14026 = x101 & n5230 ;
  assign n14027 = x100 & n5227 ;
  assign n14028 = n14026 | n14027 ;
  assign n14029 = x99 & n5434 ;
  assign n14030 = n14028 | n14029 ;
  assign n14031 = ( ~x47 & n14024 ) | ( ~x47 & n14030 ) | ( n14024 & n14030 ) ;
  assign n14032 = x47 & ~n14030 ;
  assign n14033 = ( ~n14025 & n14031 ) | ( ~n14025 & n14032 ) | ( n14031 & n14032 ) ;
  assign n14034 = n2939 & n5858 ;
  assign n14035 = x50 & n14034 ;
  assign n14036 = x98 & n5865 ;
  assign n14037 = x97 & n5862 ;
  assign n14038 = n14036 | n14037 ;
  assign n14039 = x96 & n6092 ;
  assign n14040 = n14038 | n14039 ;
  assign n14041 = ( ~x50 & n14034 ) | ( ~x50 & n14040 ) | ( n14034 & n14040 ) ;
  assign n14042 = x50 & ~n14040 ;
  assign n14043 = ( ~n14035 & n14041 ) | ( ~n14035 & n14042 ) | ( n14041 & n14042 ) ;
  assign n14044 = n2492 & n6546 ;
  assign n14045 = x53 & n14044 ;
  assign n14046 = x95 & n6553 ;
  assign n14047 = x94 & n6550 ;
  assign n14048 = n14046 | n14047 ;
  assign n14049 = x93 & n6787 ;
  assign n14050 = n14048 | n14049 ;
  assign n14051 = ( ~x53 & n14044 ) | ( ~x53 & n14050 ) | ( n14044 & n14050 ) ;
  assign n14052 = x53 & ~n14050 ;
  assign n14053 = ( ~n14045 & n14051 ) | ( ~n14045 & n14052 ) | ( n14051 & n14052 ) ;
  assign n14054 = n2083 & n7277 ;
  assign n14055 = x56 & n14054 ;
  assign n14056 = x92 & n7545 ;
  assign n14057 = x91 & n7273 ;
  assign n14058 = n14056 | n14057 ;
  assign n14059 = x90 & n7552 ;
  assign n14060 = n14058 | n14059 ;
  assign n14061 = ( ~x56 & n14054 ) | ( ~x56 & n14060 ) | ( n14054 & n14060 ) ;
  assign n14062 = x56 & ~n14060 ;
  assign n14063 = ( ~n14055 & n14061 ) | ( ~n14055 & n14062 ) | ( n14061 & n14062 ) ;
  assign n14064 = n1822 & n8067 ;
  assign n14065 = x59 & n14064 ;
  assign n14066 = x89 & n8074 ;
  assign n14067 = x88 & n8071 ;
  assign n14068 = n14066 | n14067 ;
  assign n14069 = x87 & n8298 ;
  assign n14070 = n14068 | n14069 ;
  assign n14071 = ( ~x59 & n14064 ) | ( ~x59 & n14070 ) | ( n14064 & n14070 ) ;
  assign n14072 = x59 & ~n14070 ;
  assign n14073 = ( ~n14065 & n14071 ) | ( ~n14065 & n14072 ) | ( n14071 & n14072 ) ;
  assign n14074 = n1384 & n8859 ;
  assign n14075 = x62 & n14074 ;
  assign n14076 = x86 & n8866 ;
  assign n14077 = x85 & n8863 ;
  assign n14078 = n14076 | n14077 ;
  assign n14079 = x84 & n9125 ;
  assign n14080 = n14078 | n14079 ;
  assign n14081 = ( ~x62 & n14074 ) | ( ~x62 & n14080 ) | ( n14074 & n14080 ) ;
  assign n14082 = x62 & ~n14080 ;
  assign n14083 = ( ~n14075 & n14081 ) | ( ~n14075 & n14082 ) | ( n14081 & n14082 ) ;
  assign n14084 = ( x62 & x63 ) | ( x62 & x83 ) | ( x63 & x83 ) ;
  assign n14085 = ( x62 & x82 ) | ( x62 & ~n9394 ) | ( x82 & ~n9394 ) ;
  assign n14086 = ( x82 & n14084 ) | ( x82 & ~n14085 ) | ( n14084 & ~n14085 ) ;
  assign n14087 = ( n13886 & n14083 ) | ( n13886 & ~n14086 ) | ( n14083 & ~n14086 ) ;
  assign n14088 = ( ~n13886 & n14083 ) | ( ~n13886 & n14086 ) | ( n14083 & n14086 ) ;
  assign n14089 = ( ~n14083 & n14087 ) | ( ~n14083 & n14088 ) | ( n14087 & n14088 ) ;
  assign n14090 = ( ~n13888 & n14073 ) | ( ~n13888 & n14089 ) | ( n14073 & n14089 ) ;
  assign n14091 = ( n13888 & n14073 ) | ( n13888 & ~n14089 ) | ( n14073 & ~n14089 ) ;
  assign n14092 = ( ~n14073 & n14090 ) | ( ~n14073 & n14091 ) | ( n14090 & n14091 ) ;
  assign n14093 = ( n13891 & n14063 ) | ( n13891 & ~n14092 ) | ( n14063 & ~n14092 ) ;
  assign n14094 = ( ~n13891 & n14063 ) | ( ~n13891 & n14092 ) | ( n14063 & n14092 ) ;
  assign n14095 = ( ~n14063 & n14093 ) | ( ~n14063 & n14094 ) | ( n14093 & n14094 ) ;
  assign n14096 = ( n13894 & n14053 ) | ( n13894 & ~n14095 ) | ( n14053 & ~n14095 ) ;
  assign n14097 = ( ~n13894 & n14053 ) | ( ~n13894 & n14095 ) | ( n14053 & n14095 ) ;
  assign n14098 = ( ~n14053 & n14096 ) | ( ~n14053 & n14097 ) | ( n14096 & n14097 ) ;
  assign n14099 = ( n13897 & n14043 ) | ( n13897 & ~n14098 ) | ( n14043 & ~n14098 ) ;
  assign n14100 = ( ~n13897 & n14043 ) | ( ~n13897 & n14098 ) | ( n14043 & n14098 ) ;
  assign n14101 = ( ~n14043 & n14099 ) | ( ~n14043 & n14100 ) | ( n14099 & n14100 ) ;
  assign n14102 = ( ~n13900 & n14033 ) | ( ~n13900 & n14101 ) | ( n14033 & n14101 ) ;
  assign n14103 = ( n13900 & n14033 ) | ( n13900 & ~n14101 ) | ( n14033 & ~n14101 ) ;
  assign n14104 = ( ~n14033 & n14102 ) | ( ~n14033 & n14103 ) | ( n14102 & n14103 ) ;
  assign n14105 = ( n13903 & n14023 ) | ( n13903 & ~n14104 ) | ( n14023 & ~n14104 ) ;
  assign n14106 = ( ~n13903 & n14023 ) | ( ~n13903 & n14104 ) | ( n14023 & n14104 ) ;
  assign n14107 = ( ~n14023 & n14105 ) | ( ~n14023 & n14106 ) | ( n14105 & n14106 ) ;
  assign n14108 = ( n13906 & ~n14013 ) | ( n13906 & n14107 ) | ( ~n14013 & n14107 ) ;
  assign n14109 = ( n13906 & n14013 ) | ( n13906 & n14107 ) | ( n14013 & n14107 ) ;
  assign n14110 = ( n14013 & n14108 ) | ( n14013 & ~n14109 ) | ( n14108 & ~n14109 ) ;
  assign n14111 = ( n13909 & n14003 ) | ( n13909 & n14110 ) | ( n14003 & n14110 ) ;
  assign n14112 = ( n13909 & ~n14003 ) | ( n13909 & n14110 ) | ( ~n14003 & n14110 ) ;
  assign n14113 = ( n14003 & ~n14111 ) | ( n14003 & n14112 ) | ( ~n14111 & n14112 ) ;
  assign n14114 = ( n13912 & ~n13993 ) | ( n13912 & n14113 ) | ( ~n13993 & n14113 ) ;
  assign n14115 = ( n13912 & n13993 ) | ( n13912 & n14113 ) | ( n13993 & n14113 ) ;
  assign n14116 = ( n13993 & n14114 ) | ( n13993 & ~n14115 ) | ( n14114 & ~n14115 ) ;
  assign n14117 = ( n13915 & n13983 ) | ( n13915 & n14116 ) | ( n13983 & n14116 ) ;
  assign n14118 = ( n13915 & ~n13983 ) | ( n13915 & n14116 ) | ( ~n13983 & n14116 ) ;
  assign n14119 = ( n13983 & ~n14117 ) | ( n13983 & n14118 ) | ( ~n14117 & n14118 ) ;
  assign n14120 = ( n13918 & n13973 ) | ( n13918 & n14119 ) | ( n13973 & n14119 ) ;
  assign n14121 = ( n13918 & ~n13973 ) | ( n13918 & n14119 ) | ( ~n13973 & n14119 ) ;
  assign n14122 = ( n13973 & ~n14120 ) | ( n13973 & n14121 ) | ( ~n14120 & n14121 ) ;
  assign n14123 = ( n13921 & n13963 ) | ( n13921 & n14122 ) | ( n13963 & n14122 ) ;
  assign n14124 = ( n13921 & ~n13963 ) | ( n13921 & n14122 ) | ( ~n13963 & n14122 ) ;
  assign n14125 = ( n13963 & ~n14123 ) | ( n13963 & n14124 ) | ( ~n14123 & n14124 ) ;
  assign n14126 = ( n13924 & n13953 ) | ( n13924 & n14125 ) | ( n13953 & n14125 ) ;
  assign n14127 = ( n13924 & ~n13953 ) | ( n13924 & n14125 ) | ( ~n13953 & n14125 ) ;
  assign n14128 = ( n13953 & ~n14126 ) | ( n13953 & n14127 ) | ( ~n14126 & n14127 ) ;
  assign n14129 = ( n13927 & n13943 ) | ( n13927 & n14128 ) | ( n13943 & n14128 ) ;
  assign n14130 = ( n13927 & ~n13943 ) | ( n13927 & n14128 ) | ( ~n13943 & n14128 ) ;
  assign n14131 = ( n13943 & ~n14129 ) | ( n13943 & n14130 ) | ( ~n14129 & n14130 ) ;
  assign n14132 = ( n13931 & n13933 ) | ( n13931 & n14131 ) | ( n13933 & n14131 ) ;
  assign n14133 = ( n13931 & ~n13933 ) | ( n13931 & n14131 ) | ( ~n13933 & n14131 ) ;
  assign n14134 = ( n13933 & ~n14132 ) | ( n13933 & n14133 ) | ( ~n14132 & n14133 ) ;
  assign n14135 = x127 & n1217 ;
  assign n14136 = n1146 | n14135 ;
  assign n14137 = ( n9865 & n14135 ) | ( n9865 & n14136 ) | ( n14135 & n14136 ) ;
  assign n14138 = x20 & ~n14137 ;
  assign n14139 = ~x20 & n14137 ;
  assign n14140 = n14138 | n14139 ;
  assign n14141 = n1427 & n9038 ;
  assign n14142 = x23 & n14141 ;
  assign n14143 = x126 & n1434 ;
  assign n14144 = x125 & n1431 ;
  assign n14145 = n14143 | n14144 ;
  assign n14146 = x124 & n1531 ;
  assign n14147 = n14145 | n14146 ;
  assign n14148 = ( ~x23 & n14141 ) | ( ~x23 & n14147 ) | ( n14141 & n14147 ) ;
  assign n14149 = x23 & ~n14147 ;
  assign n14150 = ( ~n14142 & n14148 ) | ( ~n14142 & n14149 ) | ( n14148 & n14149 ) ;
  assign n14151 = n1755 & n8461 ;
  assign n14152 = x26 & n14151 ;
  assign n14153 = x123 & n1762 ;
  assign n14154 = x122 & n1759 ;
  assign n14155 = n14153 | n14154 ;
  assign n14156 = x121 & n1895 ;
  assign n14157 = n14155 | n14156 ;
  assign n14158 = ( ~x26 & n14151 ) | ( ~x26 & n14157 ) | ( n14151 & n14157 ) ;
  assign n14159 = x26 & ~n14157 ;
  assign n14160 = ( ~n14152 & n14158 ) | ( ~n14152 & n14159 ) | ( n14158 & n14159 ) ;
  assign n14161 = n2137 & n7444 ;
  assign n14162 = x29 & n14161 ;
  assign n14163 = x120 & n2144 ;
  assign n14164 = x119 & n2141 ;
  assign n14165 = n14163 | n14164 ;
  assign n14166 = x118 & n2267 ;
  assign n14167 = n14165 | n14166 ;
  assign n14168 = ( ~x29 & n14161 ) | ( ~x29 & n14167 ) | ( n14161 & n14167 ) ;
  assign n14169 = x29 & ~n14167 ;
  assign n14170 = ( ~n14162 & n14168 ) | ( ~n14162 & n14169 ) | ( n14168 & n14169 ) ;
  assign n14171 = n2545 & n6924 ;
  assign n14172 = x32 & n14171 ;
  assign n14173 = x117 & n2552 ;
  assign n14174 = x116 & n2549 ;
  assign n14175 = n14173 | n14174 ;
  assign n14176 = x115 & n2696 ;
  assign n14177 = n14175 | n14176 ;
  assign n14178 = ( ~x32 & n14171 ) | ( ~x32 & n14177 ) | ( n14171 & n14177 ) ;
  assign n14179 = x32 & ~n14177 ;
  assign n14180 = ( ~n14172 & n14178 ) | ( ~n14172 & n14179 ) | ( n14178 & n14179 ) ;
  assign n14181 = n2982 & n6002 ;
  assign n14182 = x35 & n14181 ;
  assign n14183 = x114 & n2989 ;
  assign n14184 = x113 & n2986 ;
  assign n14185 = n14183 | n14184 ;
  assign n14186 = x112 & n3159 ;
  assign n14187 = n14185 | n14186 ;
  assign n14188 = ( ~x35 & n14181 ) | ( ~x35 & n14187 ) | ( n14181 & n14187 ) ;
  assign n14189 = x35 & ~n14187 ;
  assign n14190 = ( ~n14182 & n14188 ) | ( ~n14182 & n14189 ) | ( n14188 & n14189 ) ;
  assign n14191 = n3492 & n5347 ;
  assign n14192 = x38 & n14191 ;
  assign n14193 = x111 & n3499 ;
  assign n14194 = x110 & n3496 ;
  assign n14195 = n14193 | n14194 ;
  assign n14196 = x109 & n3662 ;
  assign n14197 = n14195 | n14196 ;
  assign n14198 = ( ~x38 & n14191 ) | ( ~x38 & n14197 ) | ( n14191 & n14197 ) ;
  assign n14199 = x38 & ~n14197 ;
  assign n14200 = ( ~n14192 & n14198 ) | ( ~n14192 & n14199 ) | ( n14198 & n14199 ) ;
  assign n14201 = n4020 & n4914 ;
  assign n14202 = x41 & n14201 ;
  assign n14203 = x108 & n4027 ;
  assign n14204 = x107 & n4024 ;
  assign n14205 = n14203 | n14204 ;
  assign n14206 = x106 & n4223 ;
  assign n14207 = n14205 | n14206 ;
  assign n14208 = ( ~x41 & n14201 ) | ( ~x41 & n14207 ) | ( n14201 & n14207 ) ;
  assign n14209 = x41 & ~n14207 ;
  assign n14210 = ( ~n14202 & n14208 ) | ( ~n14202 & n14209 ) | ( n14208 & n14209 ) ;
  assign n14211 = n4145 & n4625 ;
  assign n14212 = x44 & n14211 ;
  assign n14213 = x105 & n4791 ;
  assign n14214 = x104 & n4621 ;
  assign n14215 = n14213 | n14214 ;
  assign n14216 = x103 & n4795 ;
  assign n14217 = n14215 | n14216 ;
  assign n14218 = ( ~x44 & n14211 ) | ( ~x44 & n14217 ) | ( n14211 & n14217 ) ;
  assign n14219 = x44 & ~n14217 ;
  assign n14220 = ( ~n14212 & n14218 ) | ( ~n14212 & n14219 ) | ( n14218 & n14219 ) ;
  assign n14221 = n3764 & n5223 ;
  assign n14222 = x47 & n14221 ;
  assign n14223 = x102 & n5230 ;
  assign n14224 = x101 & n5227 ;
  assign n14225 = n14223 | n14224 ;
  assign n14226 = x100 & n5434 ;
  assign n14227 = n14225 | n14226 ;
  assign n14228 = ( ~x47 & n14221 ) | ( ~x47 & n14227 ) | ( n14221 & n14227 ) ;
  assign n14229 = x47 & ~n14227 ;
  assign n14230 = ( ~n14222 & n14228 ) | ( ~n14222 & n14229 ) | ( n14228 & n14229 ) ;
  assign n14231 = n3248 & n5858 ;
  assign n14232 = x50 & n14231 ;
  assign n14233 = x99 & n5865 ;
  assign n14234 = x98 & n5862 ;
  assign n14235 = n14233 | n14234 ;
  assign n14236 = x97 & n6092 ;
  assign n14237 = n14235 | n14236 ;
  assign n14238 = ( ~x50 & n14231 ) | ( ~x50 & n14237 ) | ( n14231 & n14237 ) ;
  assign n14239 = x50 & ~n14237 ;
  assign n14240 = ( ~n14232 & n14238 ) | ( ~n14232 & n14239 ) | ( n14238 & n14239 ) ;
  assign n14241 = n2772 & n6546 ;
  assign n14242 = x53 & n14241 ;
  assign n14243 = x96 & n6553 ;
  assign n14244 = x95 & n6550 ;
  assign n14245 = n14243 | n14244 ;
  assign n14246 = x94 & n6787 ;
  assign n14247 = n14245 | n14246 ;
  assign n14248 = ( ~x53 & n14241 ) | ( ~x53 & n14247 ) | ( n14241 & n14247 ) ;
  assign n14249 = x53 & ~n14247 ;
  assign n14250 = ( ~n14242 & n14248 ) | ( ~n14242 & n14249 ) | ( n14248 & n14249 ) ;
  assign n14251 = n2220 & n7277 ;
  assign n14252 = x56 & n14251 ;
  assign n14253 = x93 & n7545 ;
  assign n14254 = x92 & n7273 ;
  assign n14255 = n14253 | n14254 ;
  assign n14256 = x91 & n7552 ;
  assign n14257 = n14255 | n14256 ;
  assign n14258 = ( ~x56 & n14251 ) | ( ~x56 & n14257 ) | ( n14251 & n14257 ) ;
  assign n14259 = x56 & ~n14257 ;
  assign n14260 = ( ~n14252 & n14258 ) | ( ~n14252 & n14259 ) | ( n14258 & n14259 ) ;
  assign n14261 = n1838 & n8067 ;
  assign n14262 = x59 & n14261 ;
  assign n14263 = x90 & n8074 ;
  assign n14264 = x89 & n8071 ;
  assign n14265 = n14263 | n14264 ;
  assign n14266 = x88 & n8298 ;
  assign n14267 = n14265 | n14266 ;
  assign n14268 = ( ~x59 & n14261 ) | ( ~x59 & n14267 ) | ( n14261 & n14267 ) ;
  assign n14269 = x59 & ~n14267 ;
  assign n14270 = ( ~n14262 & n14268 ) | ( ~n14262 & n14269 ) | ( n14268 & n14269 ) ;
  assign n14271 = ( x62 & x63 ) | ( x62 & x84 ) | ( x63 & x84 ) ;
  assign n14272 = ( x62 & x83 ) | ( x62 & ~n9394 ) | ( x83 & ~n9394 ) ;
  assign n14273 = ( x83 & n14271 ) | ( x83 & ~n14272 ) | ( n14271 & ~n14272 ) ;
  assign n14274 = n1494 & n8859 ;
  assign n14275 = x62 & n14274 ;
  assign n14276 = x87 & n8866 ;
  assign n14277 = x86 & n8863 ;
  assign n14278 = n14276 | n14277 ;
  assign n14279 = x85 & n9125 ;
  assign n14280 = n14278 | n14279 ;
  assign n14281 = ( ~x62 & n14274 ) | ( ~x62 & n14280 ) | ( n14274 & n14280 ) ;
  assign n14282 = x62 & ~n14280 ;
  assign n14283 = ( ~n14275 & n14281 ) | ( ~n14275 & n14282 ) | ( n14281 & n14282 ) ;
  assign n14284 = ( n14086 & n14273 ) | ( n14086 & n14283 ) | ( n14273 & n14283 ) ;
  assign n14285 = ( n14086 & ~n14273 ) | ( n14086 & n14283 ) | ( ~n14273 & n14283 ) ;
  assign n14286 = ( n14273 & ~n14284 ) | ( n14273 & n14285 ) | ( ~n14284 & n14285 ) ;
  assign n14287 = ( n14087 & n14270 ) | ( n14087 & ~n14286 ) | ( n14270 & ~n14286 ) ;
  assign n14288 = ( ~n14087 & n14270 ) | ( ~n14087 & n14286 ) | ( n14270 & n14286 ) ;
  assign n14289 = ( ~n14270 & n14287 ) | ( ~n14270 & n14288 ) | ( n14287 & n14288 ) ;
  assign n14290 = ( n14091 & n14260 ) | ( n14091 & ~n14289 ) | ( n14260 & ~n14289 ) ;
  assign n14291 = ( ~n14091 & n14260 ) | ( ~n14091 & n14289 ) | ( n14260 & n14289 ) ;
  assign n14292 = ( ~n14260 & n14290 ) | ( ~n14260 & n14291 ) | ( n14290 & n14291 ) ;
  assign n14293 = ( n14093 & n14250 ) | ( n14093 & ~n14292 ) | ( n14250 & ~n14292 ) ;
  assign n14294 = ( ~n14093 & n14250 ) | ( ~n14093 & n14292 ) | ( n14250 & n14292 ) ;
  assign n14295 = ( ~n14250 & n14293 ) | ( ~n14250 & n14294 ) | ( n14293 & n14294 ) ;
  assign n14296 = ( n14096 & n14240 ) | ( n14096 & ~n14295 ) | ( n14240 & ~n14295 ) ;
  assign n14297 = ( ~n14096 & n14240 ) | ( ~n14096 & n14295 ) | ( n14240 & n14295 ) ;
  assign n14298 = ( ~n14240 & n14296 ) | ( ~n14240 & n14297 ) | ( n14296 & n14297 ) ;
  assign n14299 = ( n14099 & n14230 ) | ( n14099 & ~n14298 ) | ( n14230 & ~n14298 ) ;
  assign n14300 = ( ~n14099 & n14230 ) | ( ~n14099 & n14298 ) | ( n14230 & n14298 ) ;
  assign n14301 = ( ~n14230 & n14299 ) | ( ~n14230 & n14300 ) | ( n14299 & n14300 ) ;
  assign n14302 = ( n14103 & n14220 ) | ( n14103 & ~n14301 ) | ( n14220 & ~n14301 ) ;
  assign n14303 = ( ~n14103 & n14220 ) | ( ~n14103 & n14301 ) | ( n14220 & n14301 ) ;
  assign n14304 = ( ~n14220 & n14302 ) | ( ~n14220 & n14303 ) | ( n14302 & n14303 ) ;
  assign n14305 = ( n14105 & n14210 ) | ( n14105 & ~n14304 ) | ( n14210 & ~n14304 ) ;
  assign n14306 = ( ~n14105 & n14210 ) | ( ~n14105 & n14304 ) | ( n14210 & n14304 ) ;
  assign n14307 = ( ~n14210 & n14305 ) | ( ~n14210 & n14306 ) | ( n14305 & n14306 ) ;
  assign n14308 = ( n14108 & ~n14200 ) | ( n14108 & n14307 ) | ( ~n14200 & n14307 ) ;
  assign n14309 = ( n14108 & n14200 ) | ( n14108 & n14307 ) | ( n14200 & n14307 ) ;
  assign n14310 = ( n14200 & n14308 ) | ( n14200 & ~n14309 ) | ( n14308 & ~n14309 ) ;
  assign n14311 = ( n14111 & n14190 ) | ( n14111 & n14310 ) | ( n14190 & n14310 ) ;
  assign n14312 = ( n14111 & ~n14190 ) | ( n14111 & n14310 ) | ( ~n14190 & n14310 ) ;
  assign n14313 = ( n14190 & ~n14311 ) | ( n14190 & n14312 ) | ( ~n14311 & n14312 ) ;
  assign n14314 = ( n14115 & n14180 ) | ( n14115 & n14313 ) | ( n14180 & n14313 ) ;
  assign n14315 = ( n14115 & ~n14180 ) | ( n14115 & n14313 ) | ( ~n14180 & n14313 ) ;
  assign n14316 = ( n14180 & ~n14314 ) | ( n14180 & n14315 ) | ( ~n14314 & n14315 ) ;
  assign n14317 = ( n14117 & ~n14170 ) | ( n14117 & n14316 ) | ( ~n14170 & n14316 ) ;
  assign n14318 = ( n14117 & n14170 ) | ( n14117 & n14316 ) | ( n14170 & n14316 ) ;
  assign n14319 = ( n14170 & n14317 ) | ( n14170 & ~n14318 ) | ( n14317 & ~n14318 ) ;
  assign n14320 = ( n14120 & n14160 ) | ( n14120 & n14319 ) | ( n14160 & n14319 ) ;
  assign n14321 = ( n14120 & ~n14160 ) | ( n14120 & n14319 ) | ( ~n14160 & n14319 ) ;
  assign n14322 = ( n14160 & ~n14320 ) | ( n14160 & n14321 ) | ( ~n14320 & n14321 ) ;
  assign n14323 = ( n14123 & n14150 ) | ( n14123 & n14322 ) | ( n14150 & n14322 ) ;
  assign n14324 = ( n14123 & ~n14150 ) | ( n14123 & n14322 ) | ( ~n14150 & n14322 ) ;
  assign n14325 = ( n14150 & ~n14323 ) | ( n14150 & n14324 ) | ( ~n14323 & n14324 ) ;
  assign n14326 = ( n14126 & ~n14140 ) | ( n14126 & n14325 ) | ( ~n14140 & n14325 ) ;
  assign n14327 = ( n14126 & n14140 ) | ( n14126 & n14325 ) | ( n14140 & n14325 ) ;
  assign n14328 = ( n14140 & n14326 ) | ( n14140 & ~n14327 ) | ( n14326 & ~n14327 ) ;
  assign n14329 = ( n14129 & n14132 ) | ( n14129 & n14328 ) | ( n14132 & n14328 ) ;
  assign n14330 = ( n14129 & ~n14132 ) | ( n14129 & n14328 ) | ( ~n14132 & n14328 ) ;
  assign n14331 = ( n14132 & ~n14329 ) | ( n14132 & n14330 ) | ( ~n14329 & n14330 ) ;
  assign n14332 = n1427 & n9576 ;
  assign n14333 = x23 & n14332 ;
  assign n14334 = x127 & n1434 ;
  assign n14335 = x126 & n1431 ;
  assign n14336 = n14334 | n14335 ;
  assign n14337 = x125 & n1531 ;
  assign n14338 = n14336 | n14337 ;
  assign n14339 = ( ~x23 & n14332 ) | ( ~x23 & n14338 ) | ( n14332 & n14338 ) ;
  assign n14340 = x23 & ~n14338 ;
  assign n14341 = ( ~n14333 & n14339 ) | ( ~n14333 & n14340 ) | ( n14339 & n14340 ) ;
  assign n14342 = n1755 & n8729 ;
  assign n14343 = x26 & n14342 ;
  assign n14344 = x124 & n1762 ;
  assign n14345 = x123 & n1759 ;
  assign n14346 = n14344 | n14345 ;
  assign n14347 = x122 & n1895 ;
  assign n14348 = n14346 | n14347 ;
  assign n14349 = ( ~x26 & n14342 ) | ( ~x26 & n14348 ) | ( n14342 & n14348 ) ;
  assign n14350 = x26 & ~n14348 ;
  assign n14351 = ( ~n14343 & n14349 ) | ( ~n14343 & n14350 ) | ( n14349 & n14350 ) ;
  assign n14352 = n2137 & n7696 ;
  assign n14353 = x29 & n14352 ;
  assign n14354 = x121 & n2144 ;
  assign n14355 = x120 & n2141 ;
  assign n14356 = n14354 | n14355 ;
  assign n14357 = x119 & n2267 ;
  assign n14358 = n14356 | n14357 ;
  assign n14359 = ( ~x29 & n14352 ) | ( ~x29 & n14358 ) | ( n14352 & n14358 ) ;
  assign n14360 = x29 & ~n14358 ;
  assign n14361 = ( ~n14353 & n14359 ) | ( ~n14353 & n14360 ) | ( n14359 & n14360 ) ;
  assign n14362 = n2545 & n6940 ;
  assign n14363 = x32 & n14362 ;
  assign n14364 = x118 & n2552 ;
  assign n14365 = x117 & n2549 ;
  assign n14366 = n14364 | n14365 ;
  assign n14367 = x116 & n2696 ;
  assign n14368 = n14366 | n14367 ;
  assign n14369 = ( ~x32 & n14362 ) | ( ~x32 & n14368 ) | ( n14362 & n14368 ) ;
  assign n14370 = x32 & ~n14368 ;
  assign n14371 = ( ~n14363 & n14369 ) | ( ~n14363 & n14370 ) | ( n14369 & n14370 ) ;
  assign n14372 = n2982 & n6446 ;
  assign n14373 = x35 & n14372 ;
  assign n14374 = x115 & n2989 ;
  assign n14375 = x114 & n2986 ;
  assign n14376 = n14374 | n14375 ;
  assign n14377 = x113 & n3159 ;
  assign n14378 = n14376 | n14377 ;
  assign n14379 = ( ~x35 & n14372 ) | ( ~x35 & n14378 ) | ( n14372 & n14378 ) ;
  assign n14380 = x35 & ~n14378 ;
  assign n14381 = ( ~n14373 & n14379 ) | ( ~n14373 & n14380 ) | ( n14379 & n14380 ) ;
  assign n14382 = n3492 & n5558 ;
  assign n14383 = x38 & n14382 ;
  assign n14384 = x112 & n3499 ;
  assign n14385 = x111 & n3496 ;
  assign n14386 = n14384 | n14385 ;
  assign n14387 = x110 & n3662 ;
  assign n14388 = n14386 | n14387 ;
  assign n14389 = ( ~x38 & n14382 ) | ( ~x38 & n14388 ) | ( n14382 & n14388 ) ;
  assign n14390 = x38 & ~n14388 ;
  assign n14391 = ( ~n14383 & n14389 ) | ( ~n14383 & n14390 ) | ( n14389 & n14390 ) ;
  assign n14392 = n4020 & n4930 ;
  assign n14393 = x41 & n14392 ;
  assign n14394 = x109 & n4027 ;
  assign n14395 = x108 & n4024 ;
  assign n14396 = n14394 | n14395 ;
  assign n14397 = x107 & n4223 ;
  assign n14398 = n14396 | n14397 ;
  assign n14399 = ( ~x41 & n14392 ) | ( ~x41 & n14398 ) | ( n14392 & n14398 ) ;
  assign n14400 = x41 & ~n14398 ;
  assign n14401 = ( ~n14393 & n14399 ) | ( ~n14393 & n14400 ) | ( n14399 & n14400 ) ;
  assign n14402 = n4331 & n4625 ;
  assign n14403 = x44 & n14402 ;
  assign n14404 = x106 & n4791 ;
  assign n14405 = x105 & n4621 ;
  assign n14406 = n14404 | n14405 ;
  assign n14407 = x104 & n4795 ;
  assign n14408 = n14406 | n14407 ;
  assign n14409 = ( ~x44 & n14402 ) | ( ~x44 & n14408 ) | ( n14402 & n14408 ) ;
  assign n14410 = x44 & ~n14408 ;
  assign n14411 = ( ~n14403 & n14409 ) | ( ~n14403 & n14410 ) | ( n14409 & n14410 ) ;
  assign n14412 = n3941 & n5223 ;
  assign n14413 = x47 & n14412 ;
  assign n14414 = x103 & n5230 ;
  assign n14415 = x102 & n5227 ;
  assign n14416 = n14414 | n14415 ;
  assign n14417 = x101 & n5434 ;
  assign n14418 = n14416 | n14417 ;
  assign n14419 = ( ~x47 & n14412 ) | ( ~x47 & n14418 ) | ( n14412 & n14418 ) ;
  assign n14420 = x47 & ~n14418 ;
  assign n14421 = ( ~n14413 & n14419 ) | ( ~n14413 & n14420 ) | ( n14419 & n14420 ) ;
  assign n14422 = n2788 & n6546 ;
  assign n14423 = x53 & n14422 ;
  assign n14424 = x97 & n6553 ;
  assign n14425 = x96 & n6550 ;
  assign n14426 = n14424 | n14425 ;
  assign n14427 = x95 & n6787 ;
  assign n14428 = n14426 | n14427 ;
  assign n14429 = ( ~x53 & n14422 ) | ( ~x53 & n14428 ) | ( n14422 & n14428 ) ;
  assign n14430 = x53 & ~n14428 ;
  assign n14431 = ( ~n14423 & n14429 ) | ( ~n14423 & n14430 ) | ( n14429 & n14430 ) ;
  assign n14432 = n2476 & n7277 ;
  assign n14433 = x56 & n14432 ;
  assign n14434 = x94 & n7545 ;
  assign n14435 = x93 & n7273 ;
  assign n14436 = n14434 | n14435 ;
  assign n14437 = x92 & n7552 ;
  assign n14438 = n14436 | n14437 ;
  assign n14439 = ( ~x56 & n14432 ) | ( ~x56 & n14438 ) | ( n14432 & n14438 ) ;
  assign n14440 = x56 & ~n14438 ;
  assign n14441 = ( ~n14433 & n14439 ) | ( ~n14433 & n14440 ) | ( n14439 & n14440 ) ;
  assign n14442 = n1959 & n8067 ;
  assign n14443 = x59 & n14442 ;
  assign n14444 = x91 & n8074 ;
  assign n14445 = x90 & n8071 ;
  assign n14446 = n14444 | n14445 ;
  assign n14447 = x89 & n8298 ;
  assign n14448 = n14446 | n14447 ;
  assign n14449 = ( ~x59 & n14442 ) | ( ~x59 & n14448 ) | ( n14442 & n14448 ) ;
  assign n14450 = x59 & ~n14448 ;
  assign n14451 = ( ~n14443 & n14449 ) | ( ~n14443 & n14450 ) | ( n14449 & n14450 ) ;
  assign n14452 = n1602 & n8859 ;
  assign n14453 = x62 & n14452 ;
  assign n14454 = x88 & n8866 ;
  assign n14455 = x87 & n8863 ;
  assign n14456 = n14454 | n14455 ;
  assign n14457 = x86 & n9125 ;
  assign n14458 = n14456 | n14457 ;
  assign n14459 = ( ~x62 & n14452 ) | ( ~x62 & n14458 ) | ( n14452 & n14458 ) ;
  assign n14460 = x62 & ~n14458 ;
  assign n14461 = ( ~n14453 & n14459 ) | ( ~n14453 & n14460 ) | ( n14459 & n14460 ) ;
  assign n14462 = ( x62 & x63 ) | ( x62 & x85 ) | ( x63 & x85 ) ;
  assign n14463 = ( x62 & x84 ) | ( x62 & ~n9394 ) | ( x84 & ~n9394 ) ;
  assign n14464 = ( x84 & n14462 ) | ( x84 & ~n14463 ) | ( n14462 & ~n14463 ) ;
  assign n14465 = ( x20 & n14273 ) | ( x20 & n14464 ) | ( n14273 & n14464 ) ;
  assign n14466 = ( ~x20 & n14273 ) | ( ~x20 & n14464 ) | ( n14273 & n14464 ) ;
  assign n14467 = ( x20 & ~n14465 ) | ( x20 & n14466 ) | ( ~n14465 & n14466 ) ;
  assign n14468 = ( n14285 & n14461 ) | ( n14285 & ~n14467 ) | ( n14461 & ~n14467 ) ;
  assign n14469 = ( ~n14285 & n14461 ) | ( ~n14285 & n14467 ) | ( n14461 & n14467 ) ;
  assign n14470 = ( ~n14461 & n14468 ) | ( ~n14461 & n14469 ) | ( n14468 & n14469 ) ;
  assign n14471 = ( n14287 & n14451 ) | ( n14287 & ~n14470 ) | ( n14451 & ~n14470 ) ;
  assign n14472 = ( ~n14287 & n14451 ) | ( ~n14287 & n14470 ) | ( n14451 & n14470 ) ;
  assign n14473 = ( ~n14451 & n14471 ) | ( ~n14451 & n14472 ) | ( n14471 & n14472 ) ;
  assign n14474 = ( n14290 & n14441 ) | ( n14290 & ~n14473 ) | ( n14441 & ~n14473 ) ;
  assign n14475 = ( n14290 & ~n14441 ) | ( n14290 & n14473 ) | ( ~n14441 & n14473 ) ;
  assign n14476 = ( ~n14290 & n14474 ) | ( ~n14290 & n14475 ) | ( n14474 & n14475 ) ;
  assign n14477 = ( n14293 & n14431 ) | ( n14293 & ~n14476 ) | ( n14431 & ~n14476 ) ;
  assign n14478 = ( ~n14293 & n14431 ) | ( ~n14293 & n14476 ) | ( n14431 & n14476 ) ;
  assign n14479 = ( ~n14431 & n14477 ) | ( ~n14431 & n14478 ) | ( n14477 & n14478 ) ;
  assign n14480 = n3264 & n5858 ;
  assign n14481 = x50 & n14480 ;
  assign n14482 = x100 & n5865 ;
  assign n14483 = x99 & n5862 ;
  assign n14484 = n14482 | n14483 ;
  assign n14485 = x98 & n6092 ;
  assign n14486 = n14484 | n14485 ;
  assign n14487 = ( ~x50 & n14480 ) | ( ~x50 & n14486 ) | ( n14480 & n14486 ) ;
  assign n14488 = x50 & ~n14486 ;
  assign n14489 = ( ~n14481 & n14487 ) | ( ~n14481 & n14488 ) | ( n14487 & n14488 ) ;
  assign n14490 = ( n14296 & ~n14479 ) | ( n14296 & n14489 ) | ( ~n14479 & n14489 ) ;
  assign n14491 = ( n14296 & n14479 ) | ( n14296 & n14489 ) | ( n14479 & n14489 ) ;
  assign n14492 = ( n14479 & n14490 ) | ( n14479 & ~n14491 ) | ( n14490 & ~n14491 ) ;
  assign n14493 = ( n14299 & n14421 ) | ( n14299 & ~n14492 ) | ( n14421 & ~n14492 ) ;
  assign n14494 = ( n14299 & ~n14421 ) | ( n14299 & n14492 ) | ( ~n14421 & n14492 ) ;
  assign n14495 = ( ~n14299 & n14493 ) | ( ~n14299 & n14494 ) | ( n14493 & n14494 ) ;
  assign n14496 = ( n14302 & n14411 ) | ( n14302 & ~n14495 ) | ( n14411 & ~n14495 ) ;
  assign n14497 = ( n14302 & ~n14411 ) | ( n14302 & n14495 ) | ( ~n14411 & n14495 ) ;
  assign n14498 = ( ~n14302 & n14496 ) | ( ~n14302 & n14497 ) | ( n14496 & n14497 ) ;
  assign n14499 = ( n14305 & n14401 ) | ( n14305 & ~n14498 ) | ( n14401 & ~n14498 ) ;
  assign n14500 = ( n14305 & ~n14401 ) | ( n14305 & n14498 ) | ( ~n14401 & n14498 ) ;
  assign n14501 = ( ~n14305 & n14499 ) | ( ~n14305 & n14500 ) | ( n14499 & n14500 ) ;
  assign n14502 = ( n14308 & n14391 ) | ( n14308 & n14501 ) | ( n14391 & n14501 ) ;
  assign n14503 = ( n14308 & ~n14391 ) | ( n14308 & n14501 ) | ( ~n14391 & n14501 ) ;
  assign n14504 = ( n14391 & ~n14502 ) | ( n14391 & n14503 ) | ( ~n14502 & n14503 ) ;
  assign n14505 = ( n14311 & n14381 ) | ( n14311 & n14504 ) | ( n14381 & n14504 ) ;
  assign n14506 = ( ~n14311 & n14381 ) | ( ~n14311 & n14504 ) | ( n14381 & n14504 ) ;
  assign n14507 = ( n14311 & ~n14505 ) | ( n14311 & n14506 ) | ( ~n14505 & n14506 ) ;
  assign n14508 = ( n14314 & n14371 ) | ( n14314 & n14507 ) | ( n14371 & n14507 ) ;
  assign n14509 = ( ~n14314 & n14371 ) | ( ~n14314 & n14507 ) | ( n14371 & n14507 ) ;
  assign n14510 = ( n14314 & ~n14508 ) | ( n14314 & n14509 ) | ( ~n14508 & n14509 ) ;
  assign n14511 = ( n14318 & n14361 ) | ( n14318 & n14510 ) | ( n14361 & n14510 ) ;
  assign n14512 = ( ~n14318 & n14361 ) | ( ~n14318 & n14510 ) | ( n14361 & n14510 ) ;
  assign n14513 = ( n14318 & ~n14511 ) | ( n14318 & n14512 ) | ( ~n14511 & n14512 ) ;
  assign n14514 = ( n14320 & n14351 ) | ( n14320 & n14513 ) | ( n14351 & n14513 ) ;
  assign n14515 = ( ~n14320 & n14351 ) | ( ~n14320 & n14513 ) | ( n14351 & n14513 ) ;
  assign n14516 = ( n14320 & ~n14514 ) | ( n14320 & n14515 ) | ( ~n14514 & n14515 ) ;
  assign n14517 = ( n14323 & n14341 ) | ( n14323 & n14516 ) | ( n14341 & n14516 ) ;
  assign n14518 = ( ~n14323 & n14341 ) | ( ~n14323 & n14516 ) | ( n14341 & n14516 ) ;
  assign n14519 = ( n14323 & ~n14517 ) | ( n14323 & n14518 ) | ( ~n14517 & n14518 ) ;
  assign n14520 = ( n14327 & ~n14329 ) | ( n14327 & n14519 ) | ( ~n14329 & n14519 ) ;
  assign n14521 = ( n14327 & n14329 ) | ( n14327 & n14519 ) | ( n14329 & n14519 ) ;
  assign n14522 = ( n14329 & n14520 ) | ( n14329 & ~n14521 ) | ( n14520 & ~n14521 ) ;
  assign n14523 = x127 & n1431 ;
  assign n14524 = n1427 | n14523 ;
  assign n14525 = ( n9867 & n14523 ) | ( n9867 & n14524 ) | ( n14523 & n14524 ) ;
  assign n14526 = x126 & n1531 ;
  assign n14527 = ( ~x23 & n14525 ) | ( ~x23 & n14526 ) | ( n14525 & n14526 ) ;
  assign n14528 = ( x23 & ~n14525 ) | ( x23 & n14526 ) | ( ~n14525 & n14526 ) ;
  assign n14529 = ~n14526 & n14528 ;
  assign n14530 = n14527 | n14529 ;
  assign n14531 = n1755 & n9009 ;
  assign n14532 = x26 & n14531 ;
  assign n14533 = x125 & n1762 ;
  assign n14534 = x124 & n1759 ;
  assign n14535 = n14533 | n14534 ;
  assign n14536 = x123 & n1895 ;
  assign n14537 = n14535 | n14536 ;
  assign n14538 = ( ~x26 & n14531 ) | ( ~x26 & n14537 ) | ( n14531 & n14537 ) ;
  assign n14539 = x26 & ~n14537 ;
  assign n14540 = ( ~n14532 & n14538 ) | ( ~n14532 & n14539 ) | ( n14538 & n14539 ) ;
  assign n14541 = n2137 & n8207 ;
  assign n14542 = x29 & n14541 ;
  assign n14543 = x122 & n2144 ;
  assign n14544 = x121 & n2141 ;
  assign n14545 = n14543 | n14544 ;
  assign n14546 = x120 & n2267 ;
  assign n14547 = n14545 | n14546 ;
  assign n14548 = ( ~x29 & n14541 ) | ( ~x29 & n14547 ) | ( n14541 & n14547 ) ;
  assign n14549 = x29 & ~n14547 ;
  assign n14550 = ( ~n14542 & n14548 ) | ( ~n14542 & n14549 ) | ( n14548 & n14549 ) ;
  assign n14551 = n2545 & n7181 ;
  assign n14552 = x32 & n14551 ;
  assign n14553 = x119 & n2552 ;
  assign n14554 = x118 & n2549 ;
  assign n14555 = n14553 | n14554 ;
  assign n14556 = x117 & n2696 ;
  assign n14557 = n14555 | n14556 ;
  assign n14558 = ( ~x32 & n14551 ) | ( ~x32 & n14557 ) | ( n14551 & n14557 ) ;
  assign n14559 = x32 & ~n14557 ;
  assign n14560 = ( ~n14552 & n14558 ) | ( ~n14552 & n14559 ) | ( n14558 & n14559 ) ;
  assign n14561 = n2982 & n6462 ;
  assign n14562 = x35 & n14561 ;
  assign n14563 = x116 & n2989 ;
  assign n14564 = x115 & n2986 ;
  assign n14565 = n14563 | n14564 ;
  assign n14566 = x114 & n3159 ;
  assign n14567 = n14565 | n14566 ;
  assign n14568 = ( ~x35 & n14561 ) | ( ~x35 & n14567 ) | ( n14561 & n14567 ) ;
  assign n14569 = x35 & ~n14567 ;
  assign n14570 = ( ~n14562 & n14568 ) | ( ~n14562 & n14569 ) | ( n14568 & n14569 ) ;
  assign n14571 = n3492 & n5774 ;
  assign n14572 = x38 & n14571 ;
  assign n14573 = x113 & n3499 ;
  assign n14574 = x112 & n3496 ;
  assign n14575 = n14573 | n14574 ;
  assign n14576 = x111 & n3662 ;
  assign n14577 = n14575 | n14576 ;
  assign n14578 = ( ~x38 & n14571 ) | ( ~x38 & n14577 ) | ( n14571 & n14577 ) ;
  assign n14579 = x38 & ~n14577 ;
  assign n14580 = ( ~n14572 & n14578 ) | ( ~n14572 & n14579 ) | ( n14578 & n14579 ) ;
  assign n14581 = n4020 & n5331 ;
  assign n14582 = x41 & n14581 ;
  assign n14583 = x110 & n4027 ;
  assign n14584 = x109 & n4024 ;
  assign n14585 = n14583 | n14584 ;
  assign n14586 = x108 & n4223 ;
  assign n14587 = n14585 | n14586 ;
  assign n14588 = ( ~x41 & n14581 ) | ( ~x41 & n14587 ) | ( n14581 & n14587 ) ;
  assign n14589 = x41 & ~n14587 ;
  assign n14590 = ( ~n14582 & n14588 ) | ( ~n14582 & n14589 ) | ( n14588 & n14589 ) ;
  assign n14591 = n4523 & n4625 ;
  assign n14592 = x44 & n14591 ;
  assign n14593 = x107 & n4791 ;
  assign n14594 = x106 & n4621 ;
  assign n14595 = n14593 | n14594 ;
  assign n14596 = x105 & n4795 ;
  assign n14597 = n14595 | n14596 ;
  assign n14598 = ( ~x44 & n14591 ) | ( ~x44 & n14597 ) | ( n14591 & n14597 ) ;
  assign n14599 = x44 & ~n14597 ;
  assign n14600 = ( ~n14592 & n14598 ) | ( ~n14592 & n14599 ) | ( n14598 & n14599 ) ;
  assign n14601 = n3957 & n5223 ;
  assign n14602 = x47 & n14601 ;
  assign n14603 = x104 & n5230 ;
  assign n14604 = x103 & n5227 ;
  assign n14605 = n14603 | n14604 ;
  assign n14606 = x102 & n5434 ;
  assign n14607 = n14605 | n14606 ;
  assign n14608 = ( ~x47 & n14601 ) | ( ~x47 & n14607 ) | ( n14601 & n14607 ) ;
  assign n14609 = x47 & ~n14607 ;
  assign n14610 = ( ~n14602 & n14608 ) | ( ~n14602 & n14609 ) | ( n14608 & n14609 ) ;
  assign n14611 = n3591 & n5858 ;
  assign n14612 = x50 & n14611 ;
  assign n14613 = x101 & n5865 ;
  assign n14614 = x100 & n5862 ;
  assign n14615 = n14613 | n14614 ;
  assign n14616 = x99 & n6092 ;
  assign n14617 = n14615 | n14616 ;
  assign n14618 = ( ~x50 & n14611 ) | ( ~x50 & n14617 ) | ( n14611 & n14617 ) ;
  assign n14619 = x50 & ~n14617 ;
  assign n14620 = ( ~n14612 & n14618 ) | ( ~n14612 & n14619 ) | ( n14618 & n14619 ) ;
  assign n14621 = n2939 & n6546 ;
  assign n14622 = x53 & n14621 ;
  assign n14623 = x98 & n6553 ;
  assign n14624 = x97 & n6550 ;
  assign n14625 = n14623 | n14624 ;
  assign n14626 = x96 & n6787 ;
  assign n14627 = n14625 | n14626 ;
  assign n14628 = ( ~x53 & n14621 ) | ( ~x53 & n14627 ) | ( n14621 & n14627 ) ;
  assign n14629 = x53 & ~n14627 ;
  assign n14630 = ( ~n14622 & n14628 ) | ( ~n14622 & n14629 ) | ( n14628 & n14629 ) ;
  assign n14631 = n2492 & n7277 ;
  assign n14632 = x56 & n14631 ;
  assign n14633 = x95 & n7545 ;
  assign n14634 = x94 & n7273 ;
  assign n14635 = n14633 | n14634 ;
  assign n14636 = x93 & n7552 ;
  assign n14637 = n14635 | n14636 ;
  assign n14638 = ( ~x56 & n14631 ) | ( ~x56 & n14637 ) | ( n14631 & n14637 ) ;
  assign n14639 = x56 & ~n14637 ;
  assign n14640 = ( ~n14632 & n14638 ) | ( ~n14632 & n14639 ) | ( n14638 & n14639 ) ;
  assign n14641 = n2083 & n8067 ;
  assign n14642 = x59 & n14641 ;
  assign n14643 = x92 & n8074 ;
  assign n14644 = x91 & n8071 ;
  assign n14645 = n14643 | n14644 ;
  assign n14646 = x90 & n8298 ;
  assign n14647 = n14645 | n14646 ;
  assign n14648 = ( ~x59 & n14641 ) | ( ~x59 & n14647 ) | ( n14641 & n14647 ) ;
  assign n14649 = x59 & ~n14647 ;
  assign n14650 = ( ~n14642 & n14648 ) | ( ~n14642 & n14649 ) | ( n14648 & n14649 ) ;
  assign n14651 = n1822 & n8859 ;
  assign n14652 = x62 & n14651 ;
  assign n14653 = x89 & n8866 ;
  assign n14654 = x88 & n8863 ;
  assign n14655 = n14653 | n14654 ;
  assign n14656 = x87 & n9125 ;
  assign n14657 = n14655 | n14656 ;
  assign n14658 = ( ~x62 & n14651 ) | ( ~x62 & n14657 ) | ( n14651 & n14657 ) ;
  assign n14659 = x62 & ~n14657 ;
  assign n14660 = ( ~n14652 & n14658 ) | ( ~n14652 & n14659 ) | ( n14658 & n14659 ) ;
  assign n14661 = ( x62 & x63 ) | ( x62 & x86 ) | ( x63 & x86 ) ;
  assign n14662 = ( x62 & x85 ) | ( x62 & ~n9394 ) | ( x85 & ~n9394 ) ;
  assign n14663 = ( x85 & n14661 ) | ( x85 & ~n14662 ) | ( n14661 & ~n14662 ) ;
  assign n14664 = ( n14466 & n14660 ) | ( n14466 & ~n14663 ) | ( n14660 & ~n14663 ) ;
  assign n14665 = ( ~n14466 & n14660 ) | ( ~n14466 & n14663 ) | ( n14660 & n14663 ) ;
  assign n14666 = ( ~n14660 & n14664 ) | ( ~n14660 & n14665 ) | ( n14664 & n14665 ) ;
  assign n14667 = ( n14468 & n14650 ) | ( n14468 & ~n14666 ) | ( n14650 & ~n14666 ) ;
  assign n14668 = ( ~n14468 & n14650 ) | ( ~n14468 & n14666 ) | ( n14650 & n14666 ) ;
  assign n14669 = ( ~n14650 & n14667 ) | ( ~n14650 & n14668 ) | ( n14667 & n14668 ) ;
  assign n14670 = ( n14471 & n14640 ) | ( n14471 & ~n14669 ) | ( n14640 & ~n14669 ) ;
  assign n14671 = ( ~n14471 & n14640 ) | ( ~n14471 & n14669 ) | ( n14640 & n14669 ) ;
  assign n14672 = ( ~n14640 & n14670 ) | ( ~n14640 & n14671 ) | ( n14670 & n14671 ) ;
  assign n14673 = ( n14474 & n14630 ) | ( n14474 & ~n14672 ) | ( n14630 & ~n14672 ) ;
  assign n14674 = ( ~n14474 & n14630 ) | ( ~n14474 & n14672 ) | ( n14630 & n14672 ) ;
  assign n14675 = ( ~n14630 & n14673 ) | ( ~n14630 & n14674 ) | ( n14673 & n14674 ) ;
  assign n14676 = ( n14477 & n14620 ) | ( n14477 & ~n14675 ) | ( n14620 & ~n14675 ) ;
  assign n14677 = ( ~n14477 & n14620 ) | ( ~n14477 & n14675 ) | ( n14620 & n14675 ) ;
  assign n14678 = ( ~n14620 & n14676 ) | ( ~n14620 & n14677 ) | ( n14676 & n14677 ) ;
  assign n14679 = ( n14490 & n14610 ) | ( n14490 & ~n14678 ) | ( n14610 & ~n14678 ) ;
  assign n14680 = ( ~n14490 & n14610 ) | ( ~n14490 & n14678 ) | ( n14610 & n14678 ) ;
  assign n14681 = ( ~n14610 & n14679 ) | ( ~n14610 & n14680 ) | ( n14679 & n14680 ) ;
  assign n14682 = ( n14493 & n14600 ) | ( n14493 & ~n14681 ) | ( n14600 & ~n14681 ) ;
  assign n14683 = ( ~n14493 & n14600 ) | ( ~n14493 & n14681 ) | ( n14600 & n14681 ) ;
  assign n14684 = ( ~n14600 & n14682 ) | ( ~n14600 & n14683 ) | ( n14682 & n14683 ) ;
  assign n14685 = ( ~n14496 & n14590 ) | ( ~n14496 & n14684 ) | ( n14590 & n14684 ) ;
  assign n14686 = ( n14496 & n14590 ) | ( n14496 & ~n14684 ) | ( n14590 & ~n14684 ) ;
  assign n14687 = ( ~n14590 & n14685 ) | ( ~n14590 & n14686 ) | ( n14685 & n14686 ) ;
  assign n14688 = ( n14499 & n14580 ) | ( n14499 & ~n14687 ) | ( n14580 & ~n14687 ) ;
  assign n14689 = ( ~n14499 & n14580 ) | ( ~n14499 & n14687 ) | ( n14580 & n14687 ) ;
  assign n14690 = ( ~n14580 & n14688 ) | ( ~n14580 & n14689 ) | ( n14688 & n14689 ) ;
  assign n14691 = ( n14503 & ~n14570 ) | ( n14503 & n14690 ) | ( ~n14570 & n14690 ) ;
  assign n14692 = ( n14503 & n14570 ) | ( n14503 & n14690 ) | ( n14570 & n14690 ) ;
  assign n14693 = ( n14570 & n14691 ) | ( n14570 & ~n14692 ) | ( n14691 & ~n14692 ) ;
  assign n14694 = ( n14505 & n14560 ) | ( n14505 & n14693 ) | ( n14560 & n14693 ) ;
  assign n14695 = ( n14505 & ~n14560 ) | ( n14505 & n14693 ) | ( ~n14560 & n14693 ) ;
  assign n14696 = ( n14560 & ~n14694 ) | ( n14560 & n14695 ) | ( ~n14694 & n14695 ) ;
  assign n14697 = ( n14508 & n14550 ) | ( n14508 & n14696 ) | ( n14550 & n14696 ) ;
  assign n14698 = ( n14508 & ~n14550 ) | ( n14508 & n14696 ) | ( ~n14550 & n14696 ) ;
  assign n14699 = ( n14550 & ~n14697 ) | ( n14550 & n14698 ) | ( ~n14697 & n14698 ) ;
  assign n14700 = ( n14511 & n14540 ) | ( n14511 & n14699 ) | ( n14540 & n14699 ) ;
  assign n14701 = ( n14511 & ~n14540 ) | ( n14511 & n14699 ) | ( ~n14540 & n14699 ) ;
  assign n14702 = ( n14540 & ~n14700 ) | ( n14540 & n14701 ) | ( ~n14700 & n14701 ) ;
  assign n14703 = ( n14514 & n14530 ) | ( n14514 & n14702 ) | ( n14530 & n14702 ) ;
  assign n14704 = ( n14514 & ~n14530 ) | ( n14514 & n14702 ) | ( ~n14530 & n14702 ) ;
  assign n14705 = ( n14530 & ~n14703 ) | ( n14530 & n14704 ) | ( ~n14703 & n14704 ) ;
  assign n14706 = ( n14517 & n14521 ) | ( n14517 & n14705 ) | ( n14521 & n14705 ) ;
  assign n14707 = ( n14517 & ~n14521 ) | ( n14517 & n14705 ) | ( ~n14521 & n14705 ) ;
  assign n14708 = ( n14521 & ~n14706 ) | ( n14521 & n14707 ) | ( ~n14706 & n14707 ) ;
  assign n14709 = n1755 & n9038 ;
  assign n14710 = x26 & n14709 ;
  assign n14711 = x126 & n1762 ;
  assign n14712 = x125 & n1759 ;
  assign n14713 = n14711 | n14712 ;
  assign n14714 = x124 & n1895 ;
  assign n14715 = n14713 | n14714 ;
  assign n14716 = ( ~x26 & n14709 ) | ( ~x26 & n14715 ) | ( n14709 & n14715 ) ;
  assign n14717 = x26 & ~n14715 ;
  assign n14718 = ( ~n14710 & n14716 ) | ( ~n14710 & n14717 ) | ( n14716 & n14717 ) ;
  assign n14719 = n2137 & n8461 ;
  assign n14720 = x29 & n14719 ;
  assign n14721 = x123 & n2144 ;
  assign n14722 = x122 & n2141 ;
  assign n14723 = n14721 | n14722 ;
  assign n14724 = x121 & n2267 ;
  assign n14725 = n14723 | n14724 ;
  assign n14726 = ( ~x29 & n14719 ) | ( ~x29 & n14725 ) | ( n14719 & n14725 ) ;
  assign n14727 = x29 & ~n14725 ;
  assign n14728 = ( ~n14720 & n14726 ) | ( ~n14720 & n14727 ) | ( n14726 & n14727 ) ;
  assign n14729 = n2545 & n7444 ;
  assign n14730 = x32 & n14729 ;
  assign n14731 = x120 & n2552 ;
  assign n14732 = x119 & n2549 ;
  assign n14733 = n14731 | n14732 ;
  assign n14734 = x118 & n2696 ;
  assign n14735 = n14733 | n14734 ;
  assign n14736 = ( ~x32 & n14729 ) | ( ~x32 & n14735 ) | ( n14729 & n14735 ) ;
  assign n14737 = x32 & ~n14735 ;
  assign n14738 = ( ~n14730 & n14736 ) | ( ~n14730 & n14737 ) | ( n14736 & n14737 ) ;
  assign n14739 = n2982 & n6924 ;
  assign n14740 = x35 & n14739 ;
  assign n14741 = x117 & n2989 ;
  assign n14742 = x116 & n2986 ;
  assign n14743 = n14741 | n14742 ;
  assign n14744 = x115 & n3159 ;
  assign n14745 = n14743 | n14744 ;
  assign n14746 = ( ~x35 & n14739 ) | ( ~x35 & n14745 ) | ( n14739 & n14745 ) ;
  assign n14747 = x35 & ~n14745 ;
  assign n14748 = ( ~n14740 & n14746 ) | ( ~n14740 & n14747 ) | ( n14746 & n14747 ) ;
  assign n14749 = n3492 & n6002 ;
  assign n14750 = x38 & n14749 ;
  assign n14751 = x114 & n3499 ;
  assign n14752 = x113 & n3496 ;
  assign n14753 = n14751 | n14752 ;
  assign n14754 = x112 & n3662 ;
  assign n14755 = n14753 | n14754 ;
  assign n14756 = ( ~x38 & n14749 ) | ( ~x38 & n14755 ) | ( n14749 & n14755 ) ;
  assign n14757 = x38 & ~n14755 ;
  assign n14758 = ( ~n14750 & n14756 ) | ( ~n14750 & n14757 ) | ( n14756 & n14757 ) ;
  assign n14759 = n4020 & n5347 ;
  assign n14760 = x41 & n14759 ;
  assign n14761 = x111 & n4027 ;
  assign n14762 = x110 & n4024 ;
  assign n14763 = n14761 | n14762 ;
  assign n14764 = x109 & n4223 ;
  assign n14765 = n14763 | n14764 ;
  assign n14766 = ( ~x41 & n14759 ) | ( ~x41 & n14765 ) | ( n14759 & n14765 ) ;
  assign n14767 = x41 & ~n14765 ;
  assign n14768 = ( ~n14760 & n14766 ) | ( ~n14760 & n14767 ) | ( n14766 & n14767 ) ;
  assign n14769 = n4625 & n4914 ;
  assign n14770 = x44 & n14769 ;
  assign n14771 = x108 & n4791 ;
  assign n14772 = x107 & n4621 ;
  assign n14773 = n14771 | n14772 ;
  assign n14774 = x106 & n4795 ;
  assign n14775 = n14773 | n14774 ;
  assign n14776 = ( ~x44 & n14769 ) | ( ~x44 & n14775 ) | ( n14769 & n14775 ) ;
  assign n14777 = x44 & ~n14775 ;
  assign n14778 = ( ~n14770 & n14776 ) | ( ~n14770 & n14777 ) | ( n14776 & n14777 ) ;
  assign n14779 = x104 & n5227 ;
  assign n14780 = x103 | n14779 ;
  assign n14781 = ( n5434 & n14779 ) | ( n5434 & n14780 ) | ( n14779 & n14780 ) ;
  assign n14782 = n4145 & n5223 ;
  assign n14783 = n14781 | n14782 ;
  assign n14784 = x105 & n5230 ;
  assign n14785 = ( ~x47 & n14783 ) | ( ~x47 & n14784 ) | ( n14783 & n14784 ) ;
  assign n14786 = ( x47 & ~n14783 ) | ( x47 & n14784 ) | ( ~n14783 & n14784 ) ;
  assign n14787 = ~n14784 & n14786 ;
  assign n14788 = n14785 | n14787 ;
  assign n14789 = n3764 & n5858 ;
  assign n14790 = x50 & n14789 ;
  assign n14791 = x102 & n5865 ;
  assign n14792 = x101 & n5862 ;
  assign n14793 = n14791 | n14792 ;
  assign n14794 = x100 & n6092 ;
  assign n14795 = n14793 | n14794 ;
  assign n14796 = ( ~x50 & n14789 ) | ( ~x50 & n14795 ) | ( n14789 & n14795 ) ;
  assign n14797 = x50 & ~n14795 ;
  assign n14798 = ( ~n14790 & n14796 ) | ( ~n14790 & n14797 ) | ( n14796 & n14797 ) ;
  assign n14799 = n3248 & n6546 ;
  assign n14800 = x53 & n14799 ;
  assign n14801 = x99 & n6553 ;
  assign n14802 = x98 & n6550 ;
  assign n14803 = n14801 | n14802 ;
  assign n14804 = x97 & n6787 ;
  assign n14805 = n14803 | n14804 ;
  assign n14806 = ( ~x53 & n14799 ) | ( ~x53 & n14805 ) | ( n14799 & n14805 ) ;
  assign n14807 = x53 & ~n14805 ;
  assign n14808 = ( ~n14800 & n14806 ) | ( ~n14800 & n14807 ) | ( n14806 & n14807 ) ;
  assign n14809 = n2772 & n7277 ;
  assign n14810 = x56 & n14809 ;
  assign n14811 = x96 & n7545 ;
  assign n14812 = x95 & n7273 ;
  assign n14813 = n14811 | n14812 ;
  assign n14814 = x94 & n7552 ;
  assign n14815 = n14813 | n14814 ;
  assign n14816 = ( ~x56 & n14809 ) | ( ~x56 & n14815 ) | ( n14809 & n14815 ) ;
  assign n14817 = x56 & ~n14815 ;
  assign n14818 = ( ~n14810 & n14816 ) | ( ~n14810 & n14817 ) | ( n14816 & n14817 ) ;
  assign n14819 = n2220 & n8067 ;
  assign n14820 = x59 & n14819 ;
  assign n14821 = x93 & n8074 ;
  assign n14822 = x92 & n8071 ;
  assign n14823 = n14821 | n14822 ;
  assign n14824 = x91 & n8298 ;
  assign n14825 = n14823 | n14824 ;
  assign n14826 = ( ~x59 & n14819 ) | ( ~x59 & n14825 ) | ( n14819 & n14825 ) ;
  assign n14827 = x59 & ~n14825 ;
  assign n14828 = ( ~n14820 & n14826 ) | ( ~n14820 & n14827 ) | ( n14826 & n14827 ) ;
  assign n14829 = ( x62 & x63 ) | ( x62 & x87 ) | ( x63 & x87 ) ;
  assign n14830 = ( x62 & x86 ) | ( x62 & ~n9394 ) | ( x86 & ~n9394 ) ;
  assign n14831 = ( x86 & n14829 ) | ( x86 & ~n14830 ) | ( n14829 & ~n14830 ) ;
  assign n14832 = n1838 & n8859 ;
  assign n14833 = x62 & n14832 ;
  assign n14834 = x90 & n8866 ;
  assign n14835 = x89 & n8863 ;
  assign n14836 = n14834 | n14835 ;
  assign n14837 = x88 & n9125 ;
  assign n14838 = n14836 | n14837 ;
  assign n14839 = ( ~x62 & n14832 ) | ( ~x62 & n14838 ) | ( n14832 & n14838 ) ;
  assign n14840 = x62 & ~n14838 ;
  assign n14841 = ( ~n14833 & n14839 ) | ( ~n14833 & n14840 ) | ( n14839 & n14840 ) ;
  assign n14842 = ( n14663 & n14831 ) | ( n14663 & n14841 ) | ( n14831 & n14841 ) ;
  assign n14843 = ( n14663 & ~n14831 ) | ( n14663 & n14841 ) | ( ~n14831 & n14841 ) ;
  assign n14844 = ( n14831 & ~n14842 ) | ( n14831 & n14843 ) | ( ~n14842 & n14843 ) ;
  assign n14845 = ( n14664 & n14828 ) | ( n14664 & ~n14844 ) | ( n14828 & ~n14844 ) ;
  assign n14846 = ( ~n14664 & n14828 ) | ( ~n14664 & n14844 ) | ( n14828 & n14844 ) ;
  assign n14847 = ( ~n14828 & n14845 ) | ( ~n14828 & n14846 ) | ( n14845 & n14846 ) ;
  assign n14848 = ( ~n14667 & n14818 ) | ( ~n14667 & n14847 ) | ( n14818 & n14847 ) ;
  assign n14849 = ( n14667 & n14818 ) | ( n14667 & ~n14847 ) | ( n14818 & ~n14847 ) ;
  assign n14850 = ( ~n14818 & n14848 ) | ( ~n14818 & n14849 ) | ( n14848 & n14849 ) ;
  assign n14851 = ( n14670 & n14808 ) | ( n14670 & ~n14850 ) | ( n14808 & ~n14850 ) ;
  assign n14852 = ( ~n14670 & n14808 ) | ( ~n14670 & n14850 ) | ( n14808 & n14850 ) ;
  assign n14853 = ( ~n14808 & n14851 ) | ( ~n14808 & n14852 ) | ( n14851 & n14852 ) ;
  assign n14854 = ( n14673 & n14798 ) | ( n14673 & ~n14853 ) | ( n14798 & ~n14853 ) ;
  assign n14855 = ( ~n14673 & n14798 ) | ( ~n14673 & n14853 ) | ( n14798 & n14853 ) ;
  assign n14856 = ( ~n14798 & n14854 ) | ( ~n14798 & n14855 ) | ( n14854 & n14855 ) ;
  assign n14857 = ( n14676 & n14788 ) | ( n14676 & ~n14856 ) | ( n14788 & ~n14856 ) ;
  assign n14858 = ( ~n14676 & n14788 ) | ( ~n14676 & n14856 ) | ( n14788 & n14856 ) ;
  assign n14859 = ( ~n14788 & n14857 ) | ( ~n14788 & n14858 ) | ( n14857 & n14858 ) ;
  assign n14860 = ( ~n14679 & n14778 ) | ( ~n14679 & n14859 ) | ( n14778 & n14859 ) ;
  assign n14861 = ( n14679 & n14778 ) | ( n14679 & ~n14859 ) | ( n14778 & ~n14859 ) ;
  assign n14862 = ( ~n14778 & n14860 ) | ( ~n14778 & n14861 ) | ( n14860 & n14861 ) ;
  assign n14863 = ( n14682 & n14768 ) | ( n14682 & ~n14862 ) | ( n14768 & ~n14862 ) ;
  assign n14864 = ( ~n14682 & n14768 ) | ( ~n14682 & n14862 ) | ( n14768 & n14862 ) ;
  assign n14865 = ( ~n14768 & n14863 ) | ( ~n14768 & n14864 ) | ( n14863 & n14864 ) ;
  assign n14866 = ( n14686 & n14758 ) | ( n14686 & ~n14865 ) | ( n14758 & ~n14865 ) ;
  assign n14867 = ( ~n14686 & n14758 ) | ( ~n14686 & n14865 ) | ( n14758 & n14865 ) ;
  assign n14868 = ( ~n14758 & n14866 ) | ( ~n14758 & n14867 ) | ( n14866 & n14867 ) ;
  assign n14869 = ( n14688 & n14748 ) | ( n14688 & ~n14868 ) | ( n14748 & ~n14868 ) ;
  assign n14870 = ( ~n14688 & n14748 ) | ( ~n14688 & n14868 ) | ( n14748 & n14868 ) ;
  assign n14871 = ( ~n14748 & n14869 ) | ( ~n14748 & n14870 ) | ( n14869 & n14870 ) ;
  assign n14872 = ( n14691 & ~n14738 ) | ( n14691 & n14871 ) | ( ~n14738 & n14871 ) ;
  assign n14873 = ( n14691 & n14738 ) | ( n14691 & n14871 ) | ( n14738 & n14871 ) ;
  assign n14874 = ( n14738 & n14872 ) | ( n14738 & ~n14873 ) | ( n14872 & ~n14873 ) ;
  assign n14875 = ( n14694 & n14728 ) | ( n14694 & n14874 ) | ( n14728 & n14874 ) ;
  assign n14876 = ( n14694 & ~n14728 ) | ( n14694 & n14874 ) | ( ~n14728 & n14874 ) ;
  assign n14877 = ( n14728 & ~n14875 ) | ( n14728 & n14876 ) | ( ~n14875 & n14876 ) ;
  assign n14878 = ( n14697 & n14718 ) | ( n14697 & n14877 ) | ( n14718 & n14877 ) ;
  assign n14879 = ( n14697 & ~n14718 ) | ( n14697 & n14877 ) | ( ~n14718 & n14877 ) ;
  assign n14880 = ( n14718 & ~n14878 ) | ( n14718 & n14879 ) | ( ~n14878 & n14879 ) ;
  assign n14881 = x127 & n1531 ;
  assign n14882 = n1427 | n14881 ;
  assign n14883 = ( n9865 & n14881 ) | ( n9865 & n14882 ) | ( n14881 & n14882 ) ;
  assign n14884 = x23 & ~n14883 ;
  assign n14885 = ~x23 & n14883 ;
  assign n14886 = n14884 | n14885 ;
  assign n14887 = ( n14700 & n14880 ) | ( n14700 & n14886 ) | ( n14880 & n14886 ) ;
  assign n14888 = ( n14700 & ~n14880 ) | ( n14700 & n14886 ) | ( ~n14880 & n14886 ) ;
  assign n14889 = ( n14880 & ~n14887 ) | ( n14880 & n14888 ) | ( ~n14887 & n14888 ) ;
  assign n14890 = ( n14703 & n14706 ) | ( n14703 & n14889 ) | ( n14706 & n14889 ) ;
  assign n14891 = ( n14703 & ~n14706 ) | ( n14703 & n14889 ) | ( ~n14706 & n14889 ) ;
  assign n14892 = ( n14706 & ~n14890 ) | ( n14706 & n14891 ) | ( ~n14890 & n14891 ) ;
  assign n14893 = n2982 & n6940 ;
  assign n14894 = x35 & n14893 ;
  assign n14895 = x118 & n2989 ;
  assign n14896 = x117 & n2986 ;
  assign n14897 = n14895 | n14896 ;
  assign n14898 = x116 & n3159 ;
  assign n14899 = n14897 | n14898 ;
  assign n14900 = ( ~x35 & n14893 ) | ( ~x35 & n14899 ) | ( n14893 & n14899 ) ;
  assign n14901 = x35 & ~n14899 ;
  assign n14902 = ( ~n14894 & n14900 ) | ( ~n14894 & n14901 ) | ( n14900 & n14901 ) ;
  assign n14903 = n3492 & n6446 ;
  assign n14904 = x38 & n14903 ;
  assign n14905 = x115 & n3499 ;
  assign n14906 = x114 & n3496 ;
  assign n14907 = n14905 | n14906 ;
  assign n14908 = x113 & n3662 ;
  assign n14909 = n14907 | n14908 ;
  assign n14910 = ( ~x38 & n14903 ) | ( ~x38 & n14909 ) | ( n14903 & n14909 ) ;
  assign n14911 = x38 & ~n14909 ;
  assign n14912 = ( ~n14904 & n14910 ) | ( ~n14904 & n14911 ) | ( n14910 & n14911 ) ;
  assign n14913 = n4020 & n5558 ;
  assign n14914 = x41 & n14913 ;
  assign n14915 = x112 & n4027 ;
  assign n14916 = x111 & n4024 ;
  assign n14917 = n14915 | n14916 ;
  assign n14918 = x110 & n4223 ;
  assign n14919 = n14917 | n14918 ;
  assign n14920 = ( ~x41 & n14913 ) | ( ~x41 & n14919 ) | ( n14913 & n14919 ) ;
  assign n14921 = x41 & ~n14919 ;
  assign n14922 = ( ~n14914 & n14920 ) | ( ~n14914 & n14921 ) | ( n14920 & n14921 ) ;
  assign n14923 = n4625 & n4930 ;
  assign n14924 = x44 & n14923 ;
  assign n14925 = x109 & n4791 ;
  assign n14926 = x108 & n4621 ;
  assign n14927 = n14925 | n14926 ;
  assign n14928 = x107 & n4795 ;
  assign n14929 = n14927 | n14928 ;
  assign n14930 = ( ~x44 & n14923 ) | ( ~x44 & n14929 ) | ( n14923 & n14929 ) ;
  assign n14931 = x44 & ~n14929 ;
  assign n14932 = ( ~n14924 & n14930 ) | ( ~n14924 & n14931 ) | ( n14930 & n14931 ) ;
  assign n14933 = n4331 & n5223 ;
  assign n14934 = x47 & n14933 ;
  assign n14935 = x106 & n5230 ;
  assign n14936 = x105 & n5227 ;
  assign n14937 = n14935 | n14936 ;
  assign n14938 = x104 & n5434 ;
  assign n14939 = n14937 | n14938 ;
  assign n14940 = ( ~x47 & n14933 ) | ( ~x47 & n14939 ) | ( n14933 & n14939 ) ;
  assign n14941 = x47 & ~n14939 ;
  assign n14942 = ( ~n14934 & n14940 ) | ( ~n14934 & n14941 ) | ( n14940 & n14941 ) ;
  assign n14943 = n3941 & n5858 ;
  assign n14944 = x50 & n14943 ;
  assign n14945 = x103 & n5865 ;
  assign n14946 = x102 & n5862 ;
  assign n14947 = n14945 | n14946 ;
  assign n14948 = x101 & n6092 ;
  assign n14949 = n14947 | n14948 ;
  assign n14950 = ( ~x50 & n14943 ) | ( ~x50 & n14949 ) | ( n14943 & n14949 ) ;
  assign n14951 = x50 & ~n14949 ;
  assign n14952 = ( ~n14944 & n14950 ) | ( ~n14944 & n14951 ) | ( n14950 & n14951 ) ;
  assign n14953 = n3264 & n6546 ;
  assign n14954 = x53 & n14953 ;
  assign n14955 = x100 & n6553 ;
  assign n14956 = x99 & n6550 ;
  assign n14957 = n14955 | n14956 ;
  assign n14958 = x98 & n6787 ;
  assign n14959 = n14957 | n14958 ;
  assign n14960 = ( ~x53 & n14953 ) | ( ~x53 & n14959 ) | ( n14953 & n14959 ) ;
  assign n14961 = x53 & ~n14959 ;
  assign n14962 = ( ~n14954 & n14960 ) | ( ~n14954 & n14961 ) | ( n14960 & n14961 ) ;
  assign n14963 = n2788 & n7277 ;
  assign n14964 = x56 & n14963 ;
  assign n14965 = x97 & n7545 ;
  assign n14966 = x96 & n7273 ;
  assign n14967 = n14965 | n14966 ;
  assign n14968 = x95 & n7552 ;
  assign n14969 = n14967 | n14968 ;
  assign n14970 = ( ~x56 & n14963 ) | ( ~x56 & n14969 ) | ( n14963 & n14969 ) ;
  assign n14971 = x56 & ~n14969 ;
  assign n14972 = ( ~n14964 & n14970 ) | ( ~n14964 & n14971 ) | ( n14970 & n14971 ) ;
  assign n14973 = n2476 & n8067 ;
  assign n14974 = x59 & n14973 ;
  assign n14975 = x94 & n8074 ;
  assign n14976 = x93 & n8071 ;
  assign n14977 = n14975 | n14976 ;
  assign n14978 = x92 & n8298 ;
  assign n14979 = n14977 | n14978 ;
  assign n14980 = ( ~x59 & n14973 ) | ( ~x59 & n14979 ) | ( n14973 & n14979 ) ;
  assign n14981 = x59 & ~n14979 ;
  assign n14982 = ( ~n14974 & n14980 ) | ( ~n14974 & n14981 ) | ( n14980 & n14981 ) ;
  assign n14983 = n1959 & n8859 ;
  assign n14984 = x62 & n14983 ;
  assign n14985 = x91 & n8866 ;
  assign n14986 = x90 & n8863 ;
  assign n14987 = n14985 | n14986 ;
  assign n14988 = x89 & n9125 ;
  assign n14989 = n14987 | n14988 ;
  assign n14990 = ( ~x62 & n14983 ) | ( ~x62 & n14989 ) | ( n14983 & n14989 ) ;
  assign n14991 = x62 & ~n14989 ;
  assign n14992 = ( ~n14984 & n14990 ) | ( ~n14984 & n14991 ) | ( n14990 & n14991 ) ;
  assign n14993 = ( x62 & x63 ) | ( x62 & x88 ) | ( x63 & x88 ) ;
  assign n14994 = ( x62 & x87 ) | ( x62 & ~n9394 ) | ( x87 & ~n9394 ) ;
  assign n14995 = ( x87 & n14993 ) | ( x87 & ~n14994 ) | ( n14993 & ~n14994 ) ;
  assign n14996 = ( x23 & n14831 ) | ( x23 & n14995 ) | ( n14831 & n14995 ) ;
  assign n14997 = ( ~x23 & n14831 ) | ( ~x23 & n14995 ) | ( n14831 & n14995 ) ;
  assign n14998 = ( x23 & ~n14996 ) | ( x23 & n14997 ) | ( ~n14996 & n14997 ) ;
  assign n14999 = ( n14843 & n14992 ) | ( n14843 & ~n14998 ) | ( n14992 & ~n14998 ) ;
  assign n15000 = ( ~n14843 & n14992 ) | ( ~n14843 & n14998 ) | ( n14992 & n14998 ) ;
  assign n15001 = ( ~n14992 & n14999 ) | ( ~n14992 & n15000 ) | ( n14999 & n15000 ) ;
  assign n15002 = ( n14845 & n14982 ) | ( n14845 & ~n15001 ) | ( n14982 & ~n15001 ) ;
  assign n15003 = ( n14845 & ~n14982 ) | ( n14845 & n15001 ) | ( ~n14982 & n15001 ) ;
  assign n15004 = ( ~n14845 & n15002 ) | ( ~n14845 & n15003 ) | ( n15002 & n15003 ) ;
  assign n15005 = ( n14849 & n14972 ) | ( n14849 & ~n15004 ) | ( n14972 & ~n15004 ) ;
  assign n15006 = ( ~n14849 & n14972 ) | ( ~n14849 & n15004 ) | ( n14972 & n15004 ) ;
  assign n15007 = ( ~n14972 & n15005 ) | ( ~n14972 & n15006 ) | ( n15005 & n15006 ) ;
  assign n15008 = ( n14851 & n14962 ) | ( n14851 & ~n15007 ) | ( n14962 & ~n15007 ) ;
  assign n15009 = ( n14851 & ~n14962 ) | ( n14851 & n15007 ) | ( ~n14962 & n15007 ) ;
  assign n15010 = ( ~n14851 & n15008 ) | ( ~n14851 & n15009 ) | ( n15008 & n15009 ) ;
  assign n15011 = ( n14854 & n14952 ) | ( n14854 & ~n15010 ) | ( n14952 & ~n15010 ) ;
  assign n15012 = ( n14854 & ~n14952 ) | ( n14854 & n15010 ) | ( ~n14952 & n15010 ) ;
  assign n15013 = ( ~n14854 & n15011 ) | ( ~n14854 & n15012 ) | ( n15011 & n15012 ) ;
  assign n15014 = ( n14857 & n14942 ) | ( n14857 & ~n15013 ) | ( n14942 & ~n15013 ) ;
  assign n15015 = ( n14857 & ~n14942 ) | ( n14857 & n15013 ) | ( ~n14942 & n15013 ) ;
  assign n15016 = ( ~n14857 & n15014 ) | ( ~n14857 & n15015 ) | ( n15014 & n15015 ) ;
  assign n15017 = ( n14861 & n14932 ) | ( n14861 & ~n15016 ) | ( n14932 & ~n15016 ) ;
  assign n15018 = ( n14861 & ~n14932 ) | ( n14861 & n15016 ) | ( ~n14932 & n15016 ) ;
  assign n15019 = ( ~n14861 & n15017 ) | ( ~n14861 & n15018 ) | ( n15017 & n15018 ) ;
  assign n15020 = ( n14863 & n14922 ) | ( n14863 & ~n15019 ) | ( n14922 & ~n15019 ) ;
  assign n15021 = ( ~n14863 & n14922 ) | ( ~n14863 & n15019 ) | ( n14922 & n15019 ) ;
  assign n15022 = ( ~n14922 & n15020 ) | ( ~n14922 & n15021 ) | ( n15020 & n15021 ) ;
  assign n15023 = ( ~n14866 & n14912 ) | ( ~n14866 & n15022 ) | ( n14912 & n15022 ) ;
  assign n15024 = ( n14866 & n14912 ) | ( n14866 & ~n15022 ) | ( n14912 & ~n15022 ) ;
  assign n15025 = ( ~n14912 & n15023 ) | ( ~n14912 & n15024 ) | ( n15023 & n15024 ) ;
  assign n15026 = ( n14869 & n14902 ) | ( n14869 & ~n15025 ) | ( n14902 & ~n15025 ) ;
  assign n15027 = ( ~n14869 & n14902 ) | ( ~n14869 & n15025 ) | ( n14902 & n15025 ) ;
  assign n15028 = ( ~n14902 & n15026 ) | ( ~n14902 & n15027 ) | ( n15026 & n15027 ) ;
  assign n15029 = n2545 & n7696 ;
  assign n15030 = x32 & n15029 ;
  assign n15031 = x121 & n2552 ;
  assign n15032 = x120 & n2549 ;
  assign n15033 = n15031 | n15032 ;
  assign n15034 = x119 & n2696 ;
  assign n15035 = n15033 | n15034 ;
  assign n15036 = ( ~x32 & n15029 ) | ( ~x32 & n15035 ) | ( n15029 & n15035 ) ;
  assign n15037 = x32 & ~n15035 ;
  assign n15038 = ( ~n15030 & n15036 ) | ( ~n15030 & n15037 ) | ( n15036 & n15037 ) ;
  assign n15039 = ( n14872 & n15028 ) | ( n14872 & ~n15038 ) | ( n15028 & ~n15038 ) ;
  assign n15040 = ( n14872 & ~n15028 ) | ( n14872 & n15038 ) | ( ~n15028 & n15038 ) ;
  assign n15041 = ( ~n14872 & n15039 ) | ( ~n14872 & n15040 ) | ( n15039 & n15040 ) ;
  assign n15042 = n2137 & n8729 ;
  assign n15043 = x29 & n15042 ;
  assign n15044 = x124 & n2144 ;
  assign n15045 = x123 & n2141 ;
  assign n15046 = n15044 | n15045 ;
  assign n15047 = x122 & n2267 ;
  assign n15048 = n15046 | n15047 ;
  assign n15049 = ( ~x29 & n15042 ) | ( ~x29 & n15048 ) | ( n15042 & n15048 ) ;
  assign n15050 = x29 & ~n15048 ;
  assign n15051 = ( ~n15043 & n15049 ) | ( ~n15043 & n15050 ) | ( n15049 & n15050 ) ;
  assign n15052 = ( n14875 & ~n15041 ) | ( n14875 & n15051 ) | ( ~n15041 & n15051 ) ;
  assign n15053 = ( n14875 & n15041 ) | ( n14875 & n15051 ) | ( n15041 & n15051 ) ;
  assign n15054 = ( n15041 & n15052 ) | ( n15041 & ~n15053 ) | ( n15052 & ~n15053 ) ;
  assign n15055 = n1755 & n9576 ;
  assign n15056 = x26 & n15055 ;
  assign n15057 = x127 & n1762 ;
  assign n15058 = x126 & n1759 ;
  assign n15059 = n15057 | n15058 ;
  assign n15060 = x125 & n1895 ;
  assign n15061 = n15059 | n15060 ;
  assign n15062 = ( ~x26 & n15055 ) | ( ~x26 & n15061 ) | ( n15055 & n15061 ) ;
  assign n15063 = x26 & ~n15061 ;
  assign n15064 = ( ~n15056 & n15062 ) | ( ~n15056 & n15063 ) | ( n15062 & n15063 ) ;
  assign n15065 = ( n14878 & n15054 ) | ( n14878 & n15064 ) | ( n15054 & n15064 ) ;
  assign n15066 = ( ~n14878 & n15054 ) | ( ~n14878 & n15064 ) | ( n15054 & n15064 ) ;
  assign n15067 = ( n14878 & ~n15065 ) | ( n14878 & n15066 ) | ( ~n15065 & n15066 ) ;
  assign n15068 = ( n14887 & ~n14890 ) | ( n14887 & n15067 ) | ( ~n14890 & n15067 ) ;
  assign n15069 = ( n14887 & n14890 ) | ( n14887 & n15067 ) | ( n14890 & n15067 ) ;
  assign n15070 = ( n14890 & n15068 ) | ( n14890 & ~n15069 ) | ( n15068 & ~n15069 ) ;
  assign n15071 = x126 & n1895 ;
  assign n15072 = x26 & n15071 ;
  assign n15073 = x127 & n1759 ;
  assign n15074 = n1755 | n15073 ;
  assign n15075 = ( n9867 & n15073 ) | ( n9867 & n15074 ) | ( n15073 & n15074 ) ;
  assign n15076 = ( ~x26 & n15071 ) | ( ~x26 & n15075 ) | ( n15071 & n15075 ) ;
  assign n15077 = x26 & ~n15075 ;
  assign n15078 = ( ~n15072 & n15076 ) | ( ~n15072 & n15077 ) | ( n15076 & n15077 ) ;
  assign n15079 = n2137 & n9009 ;
  assign n15080 = x29 & n15079 ;
  assign n15081 = x125 & n2144 ;
  assign n15082 = x124 & n2141 ;
  assign n15083 = n15081 | n15082 ;
  assign n15084 = x123 & n2267 ;
  assign n15085 = n15083 | n15084 ;
  assign n15086 = ( ~x29 & n15079 ) | ( ~x29 & n15085 ) | ( n15079 & n15085 ) ;
  assign n15087 = x29 & ~n15085 ;
  assign n15088 = ( ~n15080 & n15086 ) | ( ~n15080 & n15087 ) | ( n15086 & n15087 ) ;
  assign n15089 = n2545 & n8207 ;
  assign n15090 = x32 & n15089 ;
  assign n15091 = x122 & n2552 ;
  assign n15092 = x121 & n2549 ;
  assign n15093 = n15091 | n15092 ;
  assign n15094 = x120 & n2696 ;
  assign n15095 = n15093 | n15094 ;
  assign n15096 = ( ~x32 & n15089 ) | ( ~x32 & n15095 ) | ( n15089 & n15095 ) ;
  assign n15097 = x32 & ~n15095 ;
  assign n15098 = ( ~n15090 & n15096 ) | ( ~n15090 & n15097 ) | ( n15096 & n15097 ) ;
  assign n15099 = n2982 & n7181 ;
  assign n15100 = x35 & n15099 ;
  assign n15101 = x119 & n2989 ;
  assign n15102 = x118 & n2986 ;
  assign n15103 = n15101 | n15102 ;
  assign n15104 = x117 & n3159 ;
  assign n15105 = n15103 | n15104 ;
  assign n15106 = ( ~x35 & n15099 ) | ( ~x35 & n15105 ) | ( n15099 & n15105 ) ;
  assign n15107 = x35 & ~n15105 ;
  assign n15108 = ( ~n15100 & n15106 ) | ( ~n15100 & n15107 ) | ( n15106 & n15107 ) ;
  assign n15109 = n3492 & n6462 ;
  assign n15110 = x38 & n15109 ;
  assign n15111 = x116 & n3499 ;
  assign n15112 = x115 & n3496 ;
  assign n15113 = n15111 | n15112 ;
  assign n15114 = x114 & n3662 ;
  assign n15115 = n15113 | n15114 ;
  assign n15116 = ( ~x38 & n15109 ) | ( ~x38 & n15115 ) | ( n15109 & n15115 ) ;
  assign n15117 = x38 & ~n15115 ;
  assign n15118 = ( ~n15110 & n15116 ) | ( ~n15110 & n15117 ) | ( n15116 & n15117 ) ;
  assign n15119 = n4020 & n5774 ;
  assign n15120 = x41 & n15119 ;
  assign n15121 = x113 & n4027 ;
  assign n15122 = x112 & n4024 ;
  assign n15123 = n15121 | n15122 ;
  assign n15124 = x111 & n4223 ;
  assign n15125 = n15123 | n15124 ;
  assign n15126 = ( ~x41 & n15119 ) | ( ~x41 & n15125 ) | ( n15119 & n15125 ) ;
  assign n15127 = x41 & ~n15125 ;
  assign n15128 = ( ~n15120 & n15126 ) | ( ~n15120 & n15127 ) | ( n15126 & n15127 ) ;
  assign n15129 = n4625 & n5331 ;
  assign n15130 = x44 & n15129 ;
  assign n15131 = x110 & n4791 ;
  assign n15132 = x109 & n4621 ;
  assign n15133 = n15131 | n15132 ;
  assign n15134 = x108 & n4795 ;
  assign n15135 = n15133 | n15134 ;
  assign n15136 = ( ~x44 & n15129 ) | ( ~x44 & n15135 ) | ( n15129 & n15135 ) ;
  assign n15137 = x44 & ~n15135 ;
  assign n15138 = ( ~n15130 & n15136 ) | ( ~n15130 & n15137 ) | ( n15136 & n15137 ) ;
  assign n15139 = n4523 & n5223 ;
  assign n15140 = x47 & n15139 ;
  assign n15141 = x107 & n5230 ;
  assign n15142 = x106 & n5227 ;
  assign n15143 = n15141 | n15142 ;
  assign n15144 = x105 & n5434 ;
  assign n15145 = n15143 | n15144 ;
  assign n15146 = ( ~x47 & n15139 ) | ( ~x47 & n15145 ) | ( n15139 & n15145 ) ;
  assign n15147 = x47 & ~n15145 ;
  assign n15148 = ( ~n15140 & n15146 ) | ( ~n15140 & n15147 ) | ( n15146 & n15147 ) ;
  assign n15149 = n3957 & n5858 ;
  assign n15150 = x50 & n15149 ;
  assign n15151 = x104 & n5865 ;
  assign n15152 = x103 & n5862 ;
  assign n15153 = n15151 | n15152 ;
  assign n15154 = x102 & n6092 ;
  assign n15155 = n15153 | n15154 ;
  assign n15156 = ( ~x50 & n15149 ) | ( ~x50 & n15155 ) | ( n15149 & n15155 ) ;
  assign n15157 = x50 & ~n15155 ;
  assign n15158 = ( ~n15150 & n15156 ) | ( ~n15150 & n15157 ) | ( n15156 & n15157 ) ;
  assign n15159 = n3591 & n6546 ;
  assign n15160 = x53 & n15159 ;
  assign n15161 = x101 & n6553 ;
  assign n15162 = x100 & n6550 ;
  assign n15163 = n15161 | n15162 ;
  assign n15164 = x99 & n6787 ;
  assign n15165 = n15163 | n15164 ;
  assign n15166 = ( ~x53 & n15159 ) | ( ~x53 & n15165 ) | ( n15159 & n15165 ) ;
  assign n15167 = x53 & ~n15165 ;
  assign n15168 = ( ~n15160 & n15166 ) | ( ~n15160 & n15167 ) | ( n15166 & n15167 ) ;
  assign n15169 = n2492 & n8067 ;
  assign n15170 = x59 & n15169 ;
  assign n15171 = x95 & n8074 ;
  assign n15172 = x94 & n8071 ;
  assign n15173 = n15171 | n15172 ;
  assign n15174 = x93 & n8298 ;
  assign n15175 = n15173 | n15174 ;
  assign n15176 = ( ~x59 & n15169 ) | ( ~x59 & n15175 ) | ( n15169 & n15175 ) ;
  assign n15177 = x59 & ~n15175 ;
  assign n15178 = ( ~n15170 & n15176 ) | ( ~n15170 & n15177 ) | ( n15176 & n15177 ) ;
  assign n15179 = n2083 & n8859 ;
  assign n15180 = x62 & n15179 ;
  assign n15181 = x92 & n8866 ;
  assign n15182 = x91 & n8863 ;
  assign n15183 = n15181 | n15182 ;
  assign n15184 = x90 & n9125 ;
  assign n15185 = n15183 | n15184 ;
  assign n15186 = ( ~x62 & n15179 ) | ( ~x62 & n15185 ) | ( n15179 & n15185 ) ;
  assign n15187 = x62 & ~n15185 ;
  assign n15188 = ( ~n15180 & n15186 ) | ( ~n15180 & n15187 ) | ( n15186 & n15187 ) ;
  assign n15189 = ( x62 & x63 ) | ( x62 & x89 ) | ( x63 & x89 ) ;
  assign n15190 = ( x62 & x88 ) | ( x62 & ~n9394 ) | ( x88 & ~n9394 ) ;
  assign n15191 = ( x88 & n15189 ) | ( x88 & ~n15190 ) | ( n15189 & ~n15190 ) ;
  assign n15192 = ( n14997 & n15188 ) | ( n14997 & ~n15191 ) | ( n15188 & ~n15191 ) ;
  assign n15193 = ( ~n14997 & n15188 ) | ( ~n14997 & n15191 ) | ( n15188 & n15191 ) ;
  assign n15194 = ( ~n15188 & n15192 ) | ( ~n15188 & n15193 ) | ( n15192 & n15193 ) ;
  assign n15195 = ( n14999 & n15178 ) | ( n14999 & ~n15194 ) | ( n15178 & ~n15194 ) ;
  assign n15196 = ( ~n14999 & n15178 ) | ( ~n14999 & n15194 ) | ( n15178 & n15194 ) ;
  assign n15197 = ( ~n15178 & n15195 ) | ( ~n15178 & n15196 ) | ( n15195 & n15196 ) ;
  assign n15198 = n2939 & n7277 ;
  assign n15199 = x56 & n15198 ;
  assign n15200 = x98 & n7545 ;
  assign n15201 = x97 & n7273 ;
  assign n15202 = n15200 | n15201 ;
  assign n15203 = x96 & n7552 ;
  assign n15204 = n15202 | n15203 ;
  assign n15205 = ( ~x56 & n15198 ) | ( ~x56 & n15204 ) | ( n15198 & n15204 ) ;
  assign n15206 = x56 & ~n15204 ;
  assign n15207 = ( ~n15199 & n15205 ) | ( ~n15199 & n15206 ) | ( n15205 & n15206 ) ;
  assign n15208 = ( n15002 & ~n15197 ) | ( n15002 & n15207 ) | ( ~n15197 & n15207 ) ;
  assign n15209 = ( n15002 & n15197 ) | ( n15002 & n15207 ) | ( n15197 & n15207 ) ;
  assign n15210 = ( n15197 & n15208 ) | ( n15197 & ~n15209 ) | ( n15208 & ~n15209 ) ;
  assign n15211 = ( n15005 & n15168 ) | ( n15005 & ~n15210 ) | ( n15168 & ~n15210 ) ;
  assign n15212 = ( ~n15005 & n15168 ) | ( ~n15005 & n15210 ) | ( n15168 & n15210 ) ;
  assign n15213 = ( ~n15168 & n15211 ) | ( ~n15168 & n15212 ) | ( n15211 & n15212 ) ;
  assign n15214 = ( n15008 & n15158 ) | ( n15008 & ~n15213 ) | ( n15158 & ~n15213 ) ;
  assign n15215 = ( ~n15008 & n15158 ) | ( ~n15008 & n15213 ) | ( n15158 & n15213 ) ;
  assign n15216 = ( ~n15158 & n15214 ) | ( ~n15158 & n15215 ) | ( n15214 & n15215 ) ;
  assign n15217 = ( n15011 & n15148 ) | ( n15011 & ~n15216 ) | ( n15148 & ~n15216 ) ;
  assign n15218 = ( ~n15011 & n15148 ) | ( ~n15011 & n15216 ) | ( n15148 & n15216 ) ;
  assign n15219 = ( ~n15148 & n15217 ) | ( ~n15148 & n15218 ) | ( n15217 & n15218 ) ;
  assign n15220 = ( n15014 & n15138 ) | ( n15014 & ~n15219 ) | ( n15138 & ~n15219 ) ;
  assign n15221 = ( ~n15014 & n15138 ) | ( ~n15014 & n15219 ) | ( n15138 & n15219 ) ;
  assign n15222 = ( ~n15138 & n15220 ) | ( ~n15138 & n15221 ) | ( n15220 & n15221 ) ;
  assign n15223 = ( n15017 & n15128 ) | ( n15017 & ~n15222 ) | ( n15128 & ~n15222 ) ;
  assign n15224 = ( ~n15017 & n15128 ) | ( ~n15017 & n15222 ) | ( n15128 & n15222 ) ;
  assign n15225 = ( ~n15128 & n15223 ) | ( ~n15128 & n15224 ) | ( n15223 & n15224 ) ;
  assign n15226 = ( ~n15020 & n15118 ) | ( ~n15020 & n15225 ) | ( n15118 & n15225 ) ;
  assign n15227 = ( n15020 & n15118 ) | ( n15020 & ~n15225 ) | ( n15118 & ~n15225 ) ;
  assign n15228 = ( ~n15118 & n15226 ) | ( ~n15118 & n15227 ) | ( n15226 & n15227 ) ;
  assign n15229 = ( n15024 & n15108 ) | ( n15024 & ~n15228 ) | ( n15108 & ~n15228 ) ;
  assign n15230 = ( ~n15024 & n15108 ) | ( ~n15024 & n15228 ) | ( n15108 & n15228 ) ;
  assign n15231 = ( ~n15108 & n15229 ) | ( ~n15108 & n15230 ) | ( n15229 & n15230 ) ;
  assign n15232 = ( n15026 & n15098 ) | ( n15026 & ~n15231 ) | ( n15098 & ~n15231 ) ;
  assign n15233 = ( ~n15026 & n15098 ) | ( ~n15026 & n15231 ) | ( n15098 & n15231 ) ;
  assign n15234 = ( ~n15098 & n15232 ) | ( ~n15098 & n15233 ) | ( n15232 & n15233 ) ;
  assign n15235 = ( n15039 & n15088 ) | ( n15039 & n15234 ) | ( n15088 & n15234 ) ;
  assign n15236 = ( n15039 & ~n15088 ) | ( n15039 & n15234 ) | ( ~n15088 & n15234 ) ;
  assign n15237 = ( n15088 & ~n15235 ) | ( n15088 & n15236 ) | ( ~n15235 & n15236 ) ;
  assign n15238 = ( n15053 & ~n15078 ) | ( n15053 & n15237 ) | ( ~n15078 & n15237 ) ;
  assign n15239 = ( n15053 & n15078 ) | ( n15053 & n15237 ) | ( n15078 & n15237 ) ;
  assign n15240 = ( n15078 & n15238 ) | ( n15078 & ~n15239 ) | ( n15238 & ~n15239 ) ;
  assign n15241 = ( n15065 & n15069 ) | ( n15065 & n15240 ) | ( n15069 & n15240 ) ;
  assign n15242 = ( n15065 & ~n15069 ) | ( n15065 & n15240 ) | ( ~n15069 & n15240 ) ;
  assign n15243 = ( n15069 & ~n15241 ) | ( n15069 & n15242 ) | ( ~n15241 & n15242 ) ;
  assign n15244 = x25 | n1759 ;
  assign n15245 = ( x127 & n1894 ) | ( x127 & n9865 ) | ( n1894 & n9865 ) ;
  assign n15246 = n15244 & n15245 ;
  assign n15247 = ( n1759 & ~n15244 ) | ( n1759 & n15245 ) | ( ~n15244 & n15245 ) ;
  assign n15248 = ( x26 & n15246 ) | ( x26 & ~n15247 ) | ( n15246 & ~n15247 ) ;
  assign n15249 = n2137 & n9038 ;
  assign n15250 = x29 & n15249 ;
  assign n15251 = x126 & n2144 ;
  assign n15252 = x125 & n2141 ;
  assign n15253 = n15251 | n15252 ;
  assign n15254 = x124 & n2267 ;
  assign n15255 = n15253 | n15254 ;
  assign n15256 = ( ~x29 & n15249 ) | ( ~x29 & n15255 ) | ( n15249 & n15255 ) ;
  assign n15257 = x29 & ~n15255 ;
  assign n15258 = ( ~n15250 & n15256 ) | ( ~n15250 & n15257 ) | ( n15256 & n15257 ) ;
  assign n15259 = n2545 & n8461 ;
  assign n15260 = x32 & n15259 ;
  assign n15261 = x123 & n2552 ;
  assign n15262 = x122 & n2549 ;
  assign n15263 = n15261 | n15262 ;
  assign n15264 = x121 & n2696 ;
  assign n15265 = n15263 | n15264 ;
  assign n15266 = ( ~x32 & n15259 ) | ( ~x32 & n15265 ) | ( n15259 & n15265 ) ;
  assign n15267 = x32 & ~n15265 ;
  assign n15268 = ( ~n15260 & n15266 ) | ( ~n15260 & n15267 ) | ( n15266 & n15267 ) ;
  assign n15269 = n2982 & n7444 ;
  assign n15270 = x35 & n15269 ;
  assign n15271 = x120 & n2989 ;
  assign n15272 = x119 & n2986 ;
  assign n15273 = n15271 | n15272 ;
  assign n15274 = x118 & n3159 ;
  assign n15275 = n15273 | n15274 ;
  assign n15276 = ( ~x35 & n15269 ) | ( ~x35 & n15275 ) | ( n15269 & n15275 ) ;
  assign n15277 = x35 & ~n15275 ;
  assign n15278 = ( ~n15270 & n15276 ) | ( ~n15270 & n15277 ) | ( n15276 & n15277 ) ;
  assign n15279 = n3492 & n6924 ;
  assign n15280 = x38 & n15279 ;
  assign n15281 = x117 & n3499 ;
  assign n15282 = x116 & n3496 ;
  assign n15283 = n15281 | n15282 ;
  assign n15284 = x115 & n3662 ;
  assign n15285 = n15283 | n15284 ;
  assign n15286 = ( ~x38 & n15279 ) | ( ~x38 & n15285 ) | ( n15279 & n15285 ) ;
  assign n15287 = x38 & ~n15285 ;
  assign n15288 = ( ~n15280 & n15286 ) | ( ~n15280 & n15287 ) | ( n15286 & n15287 ) ;
  assign n15289 = n4020 & n6002 ;
  assign n15290 = x41 & n15289 ;
  assign n15291 = x114 & n4027 ;
  assign n15292 = x113 & n4024 ;
  assign n15293 = n15291 | n15292 ;
  assign n15294 = x112 & n4223 ;
  assign n15295 = n15293 | n15294 ;
  assign n15296 = ( ~x41 & n15289 ) | ( ~x41 & n15295 ) | ( n15289 & n15295 ) ;
  assign n15297 = x41 & ~n15295 ;
  assign n15298 = ( ~n15290 & n15296 ) | ( ~n15290 & n15297 ) | ( n15296 & n15297 ) ;
  assign n15299 = n4625 & n5347 ;
  assign n15300 = x44 & n15299 ;
  assign n15301 = x111 & n4791 ;
  assign n15302 = x110 & n4621 ;
  assign n15303 = n15301 | n15302 ;
  assign n15304 = x109 & n4795 ;
  assign n15305 = n15303 | n15304 ;
  assign n15306 = ( ~x44 & n15299 ) | ( ~x44 & n15305 ) | ( n15299 & n15305 ) ;
  assign n15307 = x44 & ~n15305 ;
  assign n15308 = ( ~n15300 & n15306 ) | ( ~n15300 & n15307 ) | ( n15306 & n15307 ) ;
  assign n15309 = n4914 & n5223 ;
  assign n15310 = x47 & n15309 ;
  assign n15311 = x108 & n5230 ;
  assign n15312 = x107 & n5227 ;
  assign n15313 = n15311 | n15312 ;
  assign n15314 = x106 & n5434 ;
  assign n15315 = n15313 | n15314 ;
  assign n15316 = ( ~x47 & n15309 ) | ( ~x47 & n15315 ) | ( n15309 & n15315 ) ;
  assign n15317 = x47 & ~n15315 ;
  assign n15318 = ( ~n15310 & n15316 ) | ( ~n15310 & n15317 ) | ( n15316 & n15317 ) ;
  assign n15319 = n4145 & n5858 ;
  assign n15320 = x50 & n15319 ;
  assign n15321 = x105 & n5865 ;
  assign n15322 = x104 & n5862 ;
  assign n15323 = n15321 | n15322 ;
  assign n15324 = x103 & n6092 ;
  assign n15325 = n15323 | n15324 ;
  assign n15326 = ( ~x50 & n15319 ) | ( ~x50 & n15325 ) | ( n15319 & n15325 ) ;
  assign n15327 = x50 & ~n15325 ;
  assign n15328 = ( ~n15320 & n15326 ) | ( ~n15320 & n15327 ) | ( n15326 & n15327 ) ;
  assign n15329 = n3764 & n6546 ;
  assign n15330 = x53 & n15329 ;
  assign n15331 = x102 & n6553 ;
  assign n15332 = x101 & n6550 ;
  assign n15333 = n15331 | n15332 ;
  assign n15334 = x100 & n6787 ;
  assign n15335 = n15333 | n15334 ;
  assign n15336 = ( ~x53 & n15329 ) | ( ~x53 & n15335 ) | ( n15329 & n15335 ) ;
  assign n15337 = x53 & ~n15335 ;
  assign n15338 = ( ~n15330 & n15336 ) | ( ~n15330 & n15337 ) | ( n15336 & n15337 ) ;
  assign n15339 = n3248 & n7277 ;
  assign n15340 = x56 & n15339 ;
  assign n15341 = x99 & n7545 ;
  assign n15342 = x98 & n7273 ;
  assign n15343 = n15341 | n15342 ;
  assign n15344 = x97 & n7552 ;
  assign n15345 = n15343 | n15344 ;
  assign n15346 = ( ~x56 & n15339 ) | ( ~x56 & n15345 ) | ( n15339 & n15345 ) ;
  assign n15347 = x56 & ~n15345 ;
  assign n15348 = ( ~n15340 & n15346 ) | ( ~n15340 & n15347 ) | ( n15346 & n15347 ) ;
  assign n15349 = n2772 & n8067 ;
  assign n15350 = x59 & n15349 ;
  assign n15351 = x96 & n8074 ;
  assign n15352 = x95 & n8071 ;
  assign n15353 = n15351 | n15352 ;
  assign n15354 = x94 & n8298 ;
  assign n15355 = n15353 | n15354 ;
  assign n15356 = ( ~x59 & n15349 ) | ( ~x59 & n15355 ) | ( n15349 & n15355 ) ;
  assign n15357 = x59 & ~n15355 ;
  assign n15358 = ( ~n15350 & n15356 ) | ( ~n15350 & n15357 ) | ( n15356 & n15357 ) ;
  assign n15359 = ( x62 & x63 ) | ( x62 & x90 ) | ( x63 & x90 ) ;
  assign n15360 = ( x62 & x89 ) | ( x62 & ~n9394 ) | ( x89 & ~n9394 ) ;
  assign n15361 = ( x89 & n15359 ) | ( x89 & ~n15360 ) | ( n15359 & ~n15360 ) ;
  assign n15362 = n2220 & n8859 ;
  assign n15363 = x62 & n15362 ;
  assign n15364 = x93 & n8866 ;
  assign n15365 = x92 & n8863 ;
  assign n15366 = n15364 | n15365 ;
  assign n15367 = x91 & n9125 ;
  assign n15368 = n15366 | n15367 ;
  assign n15369 = ( ~x62 & n15362 ) | ( ~x62 & n15368 ) | ( n15362 & n15368 ) ;
  assign n15370 = x62 & ~n15368 ;
  assign n15371 = ( ~n15363 & n15369 ) | ( ~n15363 & n15370 ) | ( n15369 & n15370 ) ;
  assign n15372 = ( n15191 & n15361 ) | ( n15191 & n15371 ) | ( n15361 & n15371 ) ;
  assign n15373 = ( n15191 & ~n15361 ) | ( n15191 & n15371 ) | ( ~n15361 & n15371 ) ;
  assign n15374 = ( n15361 & ~n15372 ) | ( n15361 & n15373 ) | ( ~n15372 & n15373 ) ;
  assign n15375 = ( n15192 & n15358 ) | ( n15192 & ~n15374 ) | ( n15358 & ~n15374 ) ;
  assign n15376 = ( ~n15192 & n15358 ) | ( ~n15192 & n15374 ) | ( n15358 & n15374 ) ;
  assign n15377 = ( ~n15358 & n15375 ) | ( ~n15358 & n15376 ) | ( n15375 & n15376 ) ;
  assign n15378 = ( n15195 & n15348 ) | ( n15195 & ~n15377 ) | ( n15348 & ~n15377 ) ;
  assign n15379 = ( ~n15195 & n15348 ) | ( ~n15195 & n15377 ) | ( n15348 & n15377 ) ;
  assign n15380 = ( ~n15348 & n15378 ) | ( ~n15348 & n15379 ) | ( n15378 & n15379 ) ;
  assign n15381 = ( n15208 & n15338 ) | ( n15208 & ~n15380 ) | ( n15338 & ~n15380 ) ;
  assign n15382 = ( ~n15208 & n15338 ) | ( ~n15208 & n15380 ) | ( n15338 & n15380 ) ;
  assign n15383 = ( ~n15338 & n15381 ) | ( ~n15338 & n15382 ) | ( n15381 & n15382 ) ;
  assign n15384 = ( n15211 & n15328 ) | ( n15211 & ~n15383 ) | ( n15328 & ~n15383 ) ;
  assign n15385 = ( ~n15211 & n15328 ) | ( ~n15211 & n15383 ) | ( n15328 & n15383 ) ;
  assign n15386 = ( ~n15328 & n15384 ) | ( ~n15328 & n15385 ) | ( n15384 & n15385 ) ;
  assign n15387 = ( n15214 & n15318 ) | ( n15214 & ~n15386 ) | ( n15318 & ~n15386 ) ;
  assign n15388 = ( ~n15214 & n15318 ) | ( ~n15214 & n15386 ) | ( n15318 & n15386 ) ;
  assign n15389 = ( ~n15318 & n15387 ) | ( ~n15318 & n15388 ) | ( n15387 & n15388 ) ;
  assign n15390 = ( n15217 & n15308 ) | ( n15217 & ~n15389 ) | ( n15308 & ~n15389 ) ;
  assign n15391 = ( ~n15217 & n15308 ) | ( ~n15217 & n15389 ) | ( n15308 & n15389 ) ;
  assign n15392 = ( ~n15308 & n15390 ) | ( ~n15308 & n15391 ) | ( n15390 & n15391 ) ;
  assign n15393 = ( n15220 & n15298 ) | ( n15220 & ~n15392 ) | ( n15298 & ~n15392 ) ;
  assign n15394 = ( ~n15220 & n15298 ) | ( ~n15220 & n15392 ) | ( n15298 & n15392 ) ;
  assign n15395 = ( ~n15298 & n15393 ) | ( ~n15298 & n15394 ) | ( n15393 & n15394 ) ;
  assign n15396 = ( n15223 & n15288 ) | ( n15223 & ~n15395 ) | ( n15288 & ~n15395 ) ;
  assign n15397 = ( ~n15223 & n15288 ) | ( ~n15223 & n15395 ) | ( n15288 & n15395 ) ;
  assign n15398 = ( ~n15288 & n15396 ) | ( ~n15288 & n15397 ) | ( n15396 & n15397 ) ;
  assign n15399 = ( n15227 & n15278 ) | ( n15227 & ~n15398 ) | ( n15278 & ~n15398 ) ;
  assign n15400 = ( ~n15227 & n15278 ) | ( ~n15227 & n15398 ) | ( n15278 & n15398 ) ;
  assign n15401 = ( ~n15278 & n15399 ) | ( ~n15278 & n15400 ) | ( n15399 & n15400 ) ;
  assign n15402 = ( n15229 & n15268 ) | ( n15229 & ~n15401 ) | ( n15268 & ~n15401 ) ;
  assign n15403 = ( ~n15229 & n15268 ) | ( ~n15229 & n15401 ) | ( n15268 & n15401 ) ;
  assign n15404 = ( ~n15268 & n15402 ) | ( ~n15268 & n15403 ) | ( n15402 & n15403 ) ;
  assign n15405 = ( n15232 & n15258 ) | ( n15232 & ~n15404 ) | ( n15258 & ~n15404 ) ;
  assign n15406 = ( ~n15232 & n15258 ) | ( ~n15232 & n15404 ) | ( n15258 & n15404 ) ;
  assign n15407 = ( ~n15258 & n15405 ) | ( ~n15258 & n15406 ) | ( n15405 & n15406 ) ;
  assign n15408 = ( n15236 & n15248 ) | ( n15236 & n15407 ) | ( n15248 & n15407 ) ;
  assign n15409 = ( n15236 & ~n15248 ) | ( n15236 & n15407 ) | ( ~n15248 & n15407 ) ;
  assign n15410 = ( n15248 & ~n15408 ) | ( n15248 & n15409 ) | ( ~n15408 & n15409 ) ;
  assign n15411 = ( n15239 & n15241 ) | ( n15239 & n15410 ) | ( n15241 & n15410 ) ;
  assign n15412 = ( n15239 & ~n15241 ) | ( n15239 & n15410 ) | ( ~n15241 & n15410 ) ;
  assign n15413 = ( n15241 & ~n15411 ) | ( n15241 & n15412 ) | ( ~n15411 & n15412 ) ;
  assign n15414 = n2545 & n8729 ;
  assign n15415 = x32 & n15414 ;
  assign n15416 = x124 & n2552 ;
  assign n15417 = x123 & n2549 ;
  assign n15418 = n15416 | n15417 ;
  assign n15419 = x122 & n2696 ;
  assign n15420 = n15418 | n15419 ;
  assign n15421 = ( ~x32 & n15414 ) | ( ~x32 & n15420 ) | ( n15414 & n15420 ) ;
  assign n15422 = x32 & ~n15420 ;
  assign n15423 = ( ~n15415 & n15421 ) | ( ~n15415 & n15422 ) | ( n15421 & n15422 ) ;
  assign n15424 = n2982 & n7696 ;
  assign n15425 = x35 & n15424 ;
  assign n15426 = x121 & n2989 ;
  assign n15427 = x120 & n2986 ;
  assign n15428 = n15426 | n15427 ;
  assign n15429 = x119 & n3159 ;
  assign n15430 = n15428 | n15429 ;
  assign n15431 = ( ~x35 & n15424 ) | ( ~x35 & n15430 ) | ( n15424 & n15430 ) ;
  assign n15432 = x35 & ~n15430 ;
  assign n15433 = ( ~n15425 & n15431 ) | ( ~n15425 & n15432 ) | ( n15431 & n15432 ) ;
  assign n15434 = n3492 & n6940 ;
  assign n15435 = x38 & n15434 ;
  assign n15436 = x118 & n3499 ;
  assign n15437 = x117 & n3496 ;
  assign n15438 = n15436 | n15437 ;
  assign n15439 = x116 & n3662 ;
  assign n15440 = n15438 | n15439 ;
  assign n15441 = ( ~x38 & n15434 ) | ( ~x38 & n15440 ) | ( n15434 & n15440 ) ;
  assign n15442 = x38 & ~n15440 ;
  assign n15443 = ( ~n15435 & n15441 ) | ( ~n15435 & n15442 ) | ( n15441 & n15442 ) ;
  assign n15444 = n4020 & n6446 ;
  assign n15445 = x41 & n15444 ;
  assign n15446 = x115 & n4027 ;
  assign n15447 = x114 & n4024 ;
  assign n15448 = n15446 | n15447 ;
  assign n15449 = x113 & n4223 ;
  assign n15450 = n15448 | n15449 ;
  assign n15451 = ( ~x41 & n15444 ) | ( ~x41 & n15450 ) | ( n15444 & n15450 ) ;
  assign n15452 = x41 & ~n15450 ;
  assign n15453 = ( ~n15445 & n15451 ) | ( ~n15445 & n15452 ) | ( n15451 & n15452 ) ;
  assign n15454 = n4625 & n5558 ;
  assign n15455 = x44 & n15454 ;
  assign n15456 = x112 & n4791 ;
  assign n15457 = x111 & n4621 ;
  assign n15458 = n15456 | n15457 ;
  assign n15459 = x110 & n4795 ;
  assign n15460 = n15458 | n15459 ;
  assign n15461 = ( ~x44 & n15454 ) | ( ~x44 & n15460 ) | ( n15454 & n15460 ) ;
  assign n15462 = x44 & ~n15460 ;
  assign n15463 = ( ~n15455 & n15461 ) | ( ~n15455 & n15462 ) | ( n15461 & n15462 ) ;
  assign n15464 = n4930 & n5223 ;
  assign n15465 = x47 & n15464 ;
  assign n15466 = x109 & n5230 ;
  assign n15467 = x108 & n5227 ;
  assign n15468 = n15466 | n15467 ;
  assign n15469 = x107 & n5434 ;
  assign n15470 = n15468 | n15469 ;
  assign n15471 = ( ~x47 & n15464 ) | ( ~x47 & n15470 ) | ( n15464 & n15470 ) ;
  assign n15472 = x47 & ~n15470 ;
  assign n15473 = ( ~n15465 & n15471 ) | ( ~n15465 & n15472 ) | ( n15471 & n15472 ) ;
  assign n15474 = n4331 & n5858 ;
  assign n15475 = x50 & n15474 ;
  assign n15476 = x106 & n5865 ;
  assign n15477 = x105 & n5862 ;
  assign n15478 = n15476 | n15477 ;
  assign n15479 = x104 & n6092 ;
  assign n15480 = n15478 | n15479 ;
  assign n15481 = ( ~x50 & n15474 ) | ( ~x50 & n15480 ) | ( n15474 & n15480 ) ;
  assign n15482 = x50 & ~n15480 ;
  assign n15483 = ( ~n15475 & n15481 ) | ( ~n15475 & n15482 ) | ( n15481 & n15482 ) ;
  assign n15484 = n3941 & n6546 ;
  assign n15485 = x53 & n15484 ;
  assign n15486 = x103 & n6553 ;
  assign n15487 = x102 & n6550 ;
  assign n15488 = n15486 | n15487 ;
  assign n15489 = x101 & n6787 ;
  assign n15490 = n15488 | n15489 ;
  assign n15491 = ( ~x53 & n15484 ) | ( ~x53 & n15490 ) | ( n15484 & n15490 ) ;
  assign n15492 = x53 & ~n15490 ;
  assign n15493 = ( ~n15485 & n15491 ) | ( ~n15485 & n15492 ) | ( n15491 & n15492 ) ;
  assign n15494 = n3264 & n7277 ;
  assign n15495 = x56 & n15494 ;
  assign n15496 = x100 & n7545 ;
  assign n15497 = x99 & n7273 ;
  assign n15498 = n15496 | n15497 ;
  assign n15499 = x98 & n7552 ;
  assign n15500 = n15498 | n15499 ;
  assign n15501 = ( ~x56 & n15494 ) | ( ~x56 & n15500 ) | ( n15494 & n15500 ) ;
  assign n15502 = x56 & ~n15500 ;
  assign n15503 = ( ~n15495 & n15501 ) | ( ~n15495 & n15502 ) | ( n15501 & n15502 ) ;
  assign n15504 = n2788 & n8067 ;
  assign n15505 = x59 & n15504 ;
  assign n15506 = x97 & n8074 ;
  assign n15507 = x96 & n8071 ;
  assign n15508 = n15506 | n15507 ;
  assign n15509 = x95 & n8298 ;
  assign n15510 = n15508 | n15509 ;
  assign n15511 = ( ~x59 & n15504 ) | ( ~x59 & n15510 ) | ( n15504 & n15510 ) ;
  assign n15512 = x59 & ~n15510 ;
  assign n15513 = ( ~n15505 & n15511 ) | ( ~n15505 & n15512 ) | ( n15511 & n15512 ) ;
  assign n15514 = n2476 & n8859 ;
  assign n15515 = x62 & n15514 ;
  assign n15516 = x94 & n8866 ;
  assign n15517 = x93 & n8863 ;
  assign n15518 = n15516 | n15517 ;
  assign n15519 = x92 & n9125 ;
  assign n15520 = n15518 | n15519 ;
  assign n15521 = ( ~x62 & n15514 ) | ( ~x62 & n15520 ) | ( n15514 & n15520 ) ;
  assign n15522 = x62 & ~n15520 ;
  assign n15523 = ( ~n15515 & n15521 ) | ( ~n15515 & n15522 ) | ( n15521 & n15522 ) ;
  assign n15524 = ( x62 & x63 ) | ( x62 & x91 ) | ( x63 & x91 ) ;
  assign n15525 = ( x62 & x90 ) | ( x62 & ~n9394 ) | ( x90 & ~n9394 ) ;
  assign n15526 = ( x90 & n15524 ) | ( x90 & ~n15525 ) | ( n15524 & ~n15525 ) ;
  assign n15527 = ( x26 & n15361 ) | ( x26 & n15526 ) | ( n15361 & n15526 ) ;
  assign n15528 = ( ~x26 & n15361 ) | ( ~x26 & n15526 ) | ( n15361 & n15526 ) ;
  assign n15529 = ( x26 & ~n15527 ) | ( x26 & n15528 ) | ( ~n15527 & n15528 ) ;
  assign n15530 = ( n15373 & n15523 ) | ( n15373 & ~n15529 ) | ( n15523 & ~n15529 ) ;
  assign n15531 = ( n15373 & ~n15523 ) | ( n15373 & n15529 ) | ( ~n15523 & n15529 ) ;
  assign n15532 = ( ~n15373 & n15530 ) | ( ~n15373 & n15531 ) | ( n15530 & n15531 ) ;
  assign n15533 = ( n15375 & n15513 ) | ( n15375 & ~n15532 ) | ( n15513 & ~n15532 ) ;
  assign n15534 = ( n15375 & ~n15513 ) | ( n15375 & n15532 ) | ( ~n15513 & n15532 ) ;
  assign n15535 = ( ~n15375 & n15533 ) | ( ~n15375 & n15534 ) | ( n15533 & n15534 ) ;
  assign n15536 = ( n15378 & n15503 ) | ( n15378 & ~n15535 ) | ( n15503 & ~n15535 ) ;
  assign n15537 = ( n15378 & ~n15503 ) | ( n15378 & n15535 ) | ( ~n15503 & n15535 ) ;
  assign n15538 = ( ~n15378 & n15536 ) | ( ~n15378 & n15537 ) | ( n15536 & n15537 ) ;
  assign n15539 = ( n15381 & n15493 ) | ( n15381 & ~n15538 ) | ( n15493 & ~n15538 ) ;
  assign n15540 = ( n15381 & ~n15493 ) | ( n15381 & n15538 ) | ( ~n15493 & n15538 ) ;
  assign n15541 = ( ~n15381 & n15539 ) | ( ~n15381 & n15540 ) | ( n15539 & n15540 ) ;
  assign n15542 = ( n15384 & n15483 ) | ( n15384 & ~n15541 ) | ( n15483 & ~n15541 ) ;
  assign n15543 = ( n15384 & ~n15483 ) | ( n15384 & n15541 ) | ( ~n15483 & n15541 ) ;
  assign n15544 = ( ~n15384 & n15542 ) | ( ~n15384 & n15543 ) | ( n15542 & n15543 ) ;
  assign n15545 = ( n15387 & n15473 ) | ( n15387 & ~n15544 ) | ( n15473 & ~n15544 ) ;
  assign n15546 = ( n15387 & ~n15473 ) | ( n15387 & n15544 ) | ( ~n15473 & n15544 ) ;
  assign n15547 = ( ~n15387 & n15545 ) | ( ~n15387 & n15546 ) | ( n15545 & n15546 ) ;
  assign n15548 = ( n15390 & n15463 ) | ( n15390 & ~n15547 ) | ( n15463 & ~n15547 ) ;
  assign n15549 = ( n15390 & ~n15463 ) | ( n15390 & n15547 ) | ( ~n15463 & n15547 ) ;
  assign n15550 = ( ~n15390 & n15548 ) | ( ~n15390 & n15549 ) | ( n15548 & n15549 ) ;
  assign n15551 = ( n15393 & ~n15453 ) | ( n15393 & n15550 ) | ( ~n15453 & n15550 ) ;
  assign n15552 = ( n15393 & n15453 ) | ( n15393 & ~n15550 ) | ( n15453 & ~n15550 ) ;
  assign n15553 = ( ~n15393 & n15551 ) | ( ~n15393 & n15552 ) | ( n15551 & n15552 ) ;
  assign n15554 = ( n15396 & n15443 ) | ( n15396 & ~n15553 ) | ( n15443 & ~n15553 ) ;
  assign n15555 = ( n15396 & ~n15443 ) | ( n15396 & n15553 ) | ( ~n15443 & n15553 ) ;
  assign n15556 = ( ~n15396 & n15554 ) | ( ~n15396 & n15555 ) | ( n15554 & n15555 ) ;
  assign n15557 = ( n15399 & n15433 ) | ( n15399 & ~n15556 ) | ( n15433 & ~n15556 ) ;
  assign n15558 = ( n15399 & ~n15433 ) | ( n15399 & n15556 ) | ( ~n15433 & n15556 ) ;
  assign n15559 = ( ~n15399 & n15557 ) | ( ~n15399 & n15558 ) | ( n15557 & n15558 ) ;
  assign n15560 = ( n15402 & n15423 ) | ( n15402 & ~n15559 ) | ( n15423 & ~n15559 ) ;
  assign n15561 = ( n15402 & ~n15423 ) | ( n15402 & n15559 ) | ( ~n15423 & n15559 ) ;
  assign n15562 = ( ~n15402 & n15560 ) | ( ~n15402 & n15561 ) | ( n15560 & n15561 ) ;
  assign n15563 = x127 & n2144 ;
  assign n15564 = n2137 | n15563 ;
  assign n15565 = ( n9576 & n15563 ) | ( n9576 & n15564 ) | ( n15563 & n15564 ) ;
  assign n15566 = x125 & n2267 ;
  assign n15567 = n15565 | n15566 ;
  assign n15568 = x126 & n2141 ;
  assign n15569 = ( ~x29 & n15567 ) | ( ~x29 & n15568 ) | ( n15567 & n15568 ) ;
  assign n15570 = ( x29 & ~n15567 ) | ( x29 & n15568 ) | ( ~n15567 & n15568 ) ;
  assign n15571 = ~n15568 & n15570 ;
  assign n15572 = n15569 | n15571 ;
  assign n15573 = ( n15405 & n15562 ) | ( n15405 & ~n15572 ) | ( n15562 & ~n15572 ) ;
  assign n15574 = ( n15405 & ~n15562 ) | ( n15405 & n15572 ) | ( ~n15562 & n15572 ) ;
  assign n15575 = ( ~n15405 & n15573 ) | ( ~n15405 & n15574 ) | ( n15573 & n15574 ) ;
  assign n15576 = ( n15409 & n15411 ) | ( n15409 & n15575 ) | ( n15411 & n15575 ) ;
  assign n15577 = ( n15409 & ~n15411 ) | ( n15409 & n15575 ) | ( ~n15411 & n15575 ) ;
  assign n15578 = ( n15411 & ~n15576 ) | ( n15411 & n15577 ) | ( ~n15576 & n15577 ) ;
  assign n15579 = x127 & n2141 ;
  assign n15580 = n2137 | n15579 ;
  assign n15581 = ( n9867 & n15579 ) | ( n9867 & n15580 ) | ( n15579 & n15580 ) ;
  assign n15582 = x126 & n2267 ;
  assign n15583 = ( ~x29 & n15581 ) | ( ~x29 & n15582 ) | ( n15581 & n15582 ) ;
  assign n15584 = ( x29 & ~n15581 ) | ( x29 & n15582 ) | ( ~n15581 & n15582 ) ;
  assign n15585 = ~n15582 & n15584 ;
  assign n15586 = n15583 | n15585 ;
  assign n15587 = n2545 & n9009 ;
  assign n15588 = x32 & n15587 ;
  assign n15589 = x125 & n2552 ;
  assign n15590 = x124 & n2549 ;
  assign n15591 = n15589 | n15590 ;
  assign n15592 = x123 & n2696 ;
  assign n15593 = n15591 | n15592 ;
  assign n15594 = ( ~x32 & n15587 ) | ( ~x32 & n15593 ) | ( n15587 & n15593 ) ;
  assign n15595 = x32 & ~n15593 ;
  assign n15596 = ( ~n15588 & n15594 ) | ( ~n15588 & n15595 ) | ( n15594 & n15595 ) ;
  assign n15597 = n2982 & n8207 ;
  assign n15598 = x35 & n15597 ;
  assign n15599 = x122 & n2989 ;
  assign n15600 = x121 & n2986 ;
  assign n15601 = n15599 | n15600 ;
  assign n15602 = x120 & n3159 ;
  assign n15603 = n15601 | n15602 ;
  assign n15604 = ( ~x35 & n15597 ) | ( ~x35 & n15603 ) | ( n15597 & n15603 ) ;
  assign n15605 = x35 & ~n15603 ;
  assign n15606 = ( ~n15598 & n15604 ) | ( ~n15598 & n15605 ) | ( n15604 & n15605 ) ;
  assign n15607 = n3492 & n7181 ;
  assign n15608 = x38 & n15607 ;
  assign n15609 = x119 & n3499 ;
  assign n15610 = x118 & n3496 ;
  assign n15611 = n15609 | n15610 ;
  assign n15612 = x117 & n3662 ;
  assign n15613 = n15611 | n15612 ;
  assign n15614 = ( ~x38 & n15607 ) | ( ~x38 & n15613 ) | ( n15607 & n15613 ) ;
  assign n15615 = x38 & ~n15613 ;
  assign n15616 = ( ~n15608 & n15614 ) | ( ~n15608 & n15615 ) | ( n15614 & n15615 ) ;
  assign n15617 = n4625 & n5774 ;
  assign n15618 = x44 & n15617 ;
  assign n15619 = x113 & n4791 ;
  assign n15620 = x112 & n4621 ;
  assign n15621 = n15619 | n15620 ;
  assign n15622 = x111 & n4795 ;
  assign n15623 = n15621 | n15622 ;
  assign n15624 = ( ~x44 & n15617 ) | ( ~x44 & n15623 ) | ( n15617 & n15623 ) ;
  assign n15625 = x44 & ~n15623 ;
  assign n15626 = ( ~n15618 & n15624 ) | ( ~n15618 & n15625 ) | ( n15624 & n15625 ) ;
  assign n15627 = n5223 & n5331 ;
  assign n15628 = x47 & n15627 ;
  assign n15629 = x110 & n5230 ;
  assign n15630 = x109 & n5227 ;
  assign n15631 = n15629 | n15630 ;
  assign n15632 = x108 & n5434 ;
  assign n15633 = n15631 | n15632 ;
  assign n15634 = ( ~x47 & n15627 ) | ( ~x47 & n15633 ) | ( n15627 & n15633 ) ;
  assign n15635 = x47 & ~n15633 ;
  assign n15636 = ( ~n15628 & n15634 ) | ( ~n15628 & n15635 ) | ( n15634 & n15635 ) ;
  assign n15637 = n4523 & n5858 ;
  assign n15638 = x50 & n15637 ;
  assign n15639 = x107 & n5865 ;
  assign n15640 = x106 & n5862 ;
  assign n15641 = n15639 | n15640 ;
  assign n15642 = x105 & n6092 ;
  assign n15643 = n15641 | n15642 ;
  assign n15644 = ( ~x50 & n15637 ) | ( ~x50 & n15643 ) | ( n15637 & n15643 ) ;
  assign n15645 = x50 & ~n15643 ;
  assign n15646 = ( ~n15638 & n15644 ) | ( ~n15638 & n15645 ) | ( n15644 & n15645 ) ;
  assign n15647 = n3957 & n6546 ;
  assign n15648 = x53 & n15647 ;
  assign n15649 = x104 & n6553 ;
  assign n15650 = x103 & n6550 ;
  assign n15651 = n15649 | n15650 ;
  assign n15652 = x102 & n6787 ;
  assign n15653 = n15651 | n15652 ;
  assign n15654 = ( ~x53 & n15647 ) | ( ~x53 & n15653 ) | ( n15647 & n15653 ) ;
  assign n15655 = x53 & ~n15653 ;
  assign n15656 = ( ~n15648 & n15654 ) | ( ~n15648 & n15655 ) | ( n15654 & n15655 ) ;
  assign n15657 = n3591 & n7277 ;
  assign n15658 = x56 & n15657 ;
  assign n15659 = x101 & n7545 ;
  assign n15660 = x100 & n7273 ;
  assign n15661 = n15659 | n15660 ;
  assign n15662 = x99 & n7552 ;
  assign n15663 = n15661 | n15662 ;
  assign n15664 = ( ~x56 & n15657 ) | ( ~x56 & n15663 ) | ( n15657 & n15663 ) ;
  assign n15665 = x56 & ~n15663 ;
  assign n15666 = ( ~n15658 & n15664 ) | ( ~n15658 & n15665 ) | ( n15664 & n15665 ) ;
  assign n15667 = n2939 & n8067 ;
  assign n15668 = x59 & n15667 ;
  assign n15669 = x98 & n8074 ;
  assign n15670 = x97 & n8071 ;
  assign n15671 = n15669 | n15670 ;
  assign n15672 = x96 & n8298 ;
  assign n15673 = n15671 | n15672 ;
  assign n15674 = ( ~x59 & n15667 ) | ( ~x59 & n15673 ) | ( n15667 & n15673 ) ;
  assign n15675 = x59 & ~n15673 ;
  assign n15676 = ( ~n15668 & n15674 ) | ( ~n15668 & n15675 ) | ( n15674 & n15675 ) ;
  assign n15677 = ( x62 & x63 ) | ( x62 & x92 ) | ( x63 & x92 ) ;
  assign n15678 = ( x62 & x91 ) | ( x62 & ~n9394 ) | ( x91 & ~n9394 ) ;
  assign n15679 = ( x91 & n15677 ) | ( x91 & ~n15678 ) | ( n15677 & ~n15678 ) ;
  assign n15680 = n2492 & n8859 ;
  assign n15681 = x62 & n15680 ;
  assign n15682 = x95 & n8866 ;
  assign n15683 = x94 & n8863 ;
  assign n15684 = n15682 | n15683 ;
  assign n15685 = x93 & n9125 ;
  assign n15686 = n15684 | n15685 ;
  assign n15687 = ( ~x62 & n15680 ) | ( ~x62 & n15686 ) | ( n15680 & n15686 ) ;
  assign n15688 = x62 & ~n15686 ;
  assign n15689 = ( ~n15681 & n15687 ) | ( ~n15681 & n15688 ) | ( n15687 & n15688 ) ;
  assign n15690 = ( ~n15528 & n15679 ) | ( ~n15528 & n15689 ) | ( n15679 & n15689 ) ;
  assign n15691 = ( n15528 & n15679 ) | ( n15528 & ~n15689 ) | ( n15679 & ~n15689 ) ;
  assign n15692 = ( ~n15679 & n15690 ) | ( ~n15679 & n15691 ) | ( n15690 & n15691 ) ;
  assign n15693 = ( n15530 & n15676 ) | ( n15530 & ~n15692 ) | ( n15676 & ~n15692 ) ;
  assign n15694 = ( ~n15530 & n15676 ) | ( ~n15530 & n15692 ) | ( n15676 & n15692 ) ;
  assign n15695 = ( ~n15676 & n15693 ) | ( ~n15676 & n15694 ) | ( n15693 & n15694 ) ;
  assign n15696 = ( n15533 & n15666 ) | ( n15533 & ~n15695 ) | ( n15666 & ~n15695 ) ;
  assign n15697 = ( ~n15533 & n15666 ) | ( ~n15533 & n15695 ) | ( n15666 & n15695 ) ;
  assign n15698 = ( ~n15666 & n15696 ) | ( ~n15666 & n15697 ) | ( n15696 & n15697 ) ;
  assign n15699 = ( n15536 & n15656 ) | ( n15536 & ~n15698 ) | ( n15656 & ~n15698 ) ;
  assign n15700 = ( ~n15536 & n15656 ) | ( ~n15536 & n15698 ) | ( n15656 & n15698 ) ;
  assign n15701 = ( ~n15656 & n15699 ) | ( ~n15656 & n15700 ) | ( n15699 & n15700 ) ;
  assign n15702 = ( n15539 & n15646 ) | ( n15539 & ~n15701 ) | ( n15646 & ~n15701 ) ;
  assign n15703 = ( ~n15539 & n15646 ) | ( ~n15539 & n15701 ) | ( n15646 & n15701 ) ;
  assign n15704 = ( ~n15646 & n15702 ) | ( ~n15646 & n15703 ) | ( n15702 & n15703 ) ;
  assign n15705 = ( ~n15542 & n15636 ) | ( ~n15542 & n15704 ) | ( n15636 & n15704 ) ;
  assign n15706 = ( n15542 & n15636 ) | ( n15542 & ~n15704 ) | ( n15636 & ~n15704 ) ;
  assign n15707 = ( ~n15636 & n15705 ) | ( ~n15636 & n15706 ) | ( n15705 & n15706 ) ;
  assign n15708 = ( n15545 & n15626 ) | ( n15545 & ~n15707 ) | ( n15626 & ~n15707 ) ;
  assign n15709 = ( ~n15545 & n15626 ) | ( ~n15545 & n15707 ) | ( n15626 & n15707 ) ;
  assign n15710 = ( ~n15626 & n15708 ) | ( ~n15626 & n15709 ) | ( n15708 & n15709 ) ;
  assign n15711 = n4020 & n6462 ;
  assign n15712 = x41 & n15711 ;
  assign n15713 = x116 & n4027 ;
  assign n15714 = x115 & n4024 ;
  assign n15715 = n15713 | n15714 ;
  assign n15716 = x114 & n4223 ;
  assign n15717 = n15715 | n15716 ;
  assign n15718 = ( ~x41 & n15711 ) | ( ~x41 & n15717 ) | ( n15711 & n15717 ) ;
  assign n15719 = x41 & ~n15717 ;
  assign n15720 = ( ~n15712 & n15718 ) | ( ~n15712 & n15719 ) | ( n15718 & n15719 ) ;
  assign n15721 = ( n15548 & ~n15710 ) | ( n15548 & n15720 ) | ( ~n15710 & n15720 ) ;
  assign n15722 = ( n15548 & n15710 ) | ( n15548 & n15720 ) | ( n15710 & n15720 ) ;
  assign n15723 = ( n15710 & n15721 ) | ( n15710 & ~n15722 ) | ( n15721 & ~n15722 ) ;
  assign n15724 = ( n15552 & n15616 ) | ( n15552 & ~n15723 ) | ( n15616 & ~n15723 ) ;
  assign n15725 = ( ~n15552 & n15616 ) | ( ~n15552 & n15723 ) | ( n15616 & n15723 ) ;
  assign n15726 = ( ~n15616 & n15724 ) | ( ~n15616 & n15725 ) | ( n15724 & n15725 ) ;
  assign n15727 = ( n15554 & n15606 ) | ( n15554 & ~n15726 ) | ( n15606 & ~n15726 ) ;
  assign n15728 = ( ~n15554 & n15606 ) | ( ~n15554 & n15726 ) | ( n15606 & n15726 ) ;
  assign n15729 = ( ~n15606 & n15727 ) | ( ~n15606 & n15728 ) | ( n15727 & n15728 ) ;
  assign n15730 = ( n15557 & n15596 ) | ( n15557 & ~n15729 ) | ( n15596 & ~n15729 ) ;
  assign n15731 = ( ~n15557 & n15596 ) | ( ~n15557 & n15729 ) | ( n15596 & n15729 ) ;
  assign n15732 = ( ~n15596 & n15730 ) | ( ~n15596 & n15731 ) | ( n15730 & n15731 ) ;
  assign n15733 = ( n15560 & n15586 ) | ( n15560 & ~n15732 ) | ( n15586 & ~n15732 ) ;
  assign n15734 = ( ~n15560 & n15586 ) | ( ~n15560 & n15732 ) | ( n15586 & n15732 ) ;
  assign n15735 = ( ~n15586 & n15733 ) | ( ~n15586 & n15734 ) | ( n15733 & n15734 ) ;
  assign n15736 = ( ~n15574 & n15577 ) | ( ~n15574 & n15735 ) | ( n15577 & n15735 ) ;
  assign n15737 = ( n15574 & n15577 ) | ( n15574 & ~n15735 ) | ( n15577 & ~n15735 ) ;
  assign n15738 = ( ~n15577 & n15736 ) | ( ~n15577 & n15737 ) | ( n15736 & n15737 ) ;
  assign n15739 = n2545 & n9038 ;
  assign n15740 = x32 & n15739 ;
  assign n15741 = x126 & n2552 ;
  assign n15742 = x125 & n2549 ;
  assign n15743 = n15741 | n15742 ;
  assign n15744 = x124 & n2696 ;
  assign n15745 = n15743 | n15744 ;
  assign n15746 = ( ~x32 & n15739 ) | ( ~x32 & n15745 ) | ( n15739 & n15745 ) ;
  assign n15747 = x32 & ~n15745 ;
  assign n15748 = ( ~n15740 & n15746 ) | ( ~n15740 & n15747 ) | ( n15746 & n15747 ) ;
  assign n15749 = n2982 & n8461 ;
  assign n15750 = x35 & n15749 ;
  assign n15751 = x123 & n2989 ;
  assign n15752 = x122 & n2986 ;
  assign n15753 = n15751 | n15752 ;
  assign n15754 = x121 & n3159 ;
  assign n15755 = n15753 | n15754 ;
  assign n15756 = ( ~x35 & n15749 ) | ( ~x35 & n15755 ) | ( n15749 & n15755 ) ;
  assign n15757 = x35 & ~n15755 ;
  assign n15758 = ( ~n15750 & n15756 ) | ( ~n15750 & n15757 ) | ( n15756 & n15757 ) ;
  assign n15759 = n3492 & n7444 ;
  assign n15760 = x38 & n15759 ;
  assign n15761 = x120 & n3499 ;
  assign n15762 = x119 & n3496 ;
  assign n15763 = n15761 | n15762 ;
  assign n15764 = x118 & n3662 ;
  assign n15765 = n15763 | n15764 ;
  assign n15766 = ( ~x38 & n15759 ) | ( ~x38 & n15765 ) | ( n15759 & n15765 ) ;
  assign n15767 = x38 & ~n15765 ;
  assign n15768 = ( ~n15760 & n15766 ) | ( ~n15760 & n15767 ) | ( n15766 & n15767 ) ;
  assign n15769 = n4020 & n6924 ;
  assign n15770 = x41 & n15769 ;
  assign n15771 = x117 & n4027 ;
  assign n15772 = x116 & n4024 ;
  assign n15773 = n15771 | n15772 ;
  assign n15774 = x115 & n4223 ;
  assign n15775 = n15773 | n15774 ;
  assign n15776 = ( ~x41 & n15769 ) | ( ~x41 & n15775 ) | ( n15769 & n15775 ) ;
  assign n15777 = x41 & ~n15775 ;
  assign n15778 = ( ~n15770 & n15776 ) | ( ~n15770 & n15777 ) | ( n15776 & n15777 ) ;
  assign n15779 = n4625 & n6002 ;
  assign n15780 = x44 & n15779 ;
  assign n15781 = x114 & n4791 ;
  assign n15782 = x113 & n4621 ;
  assign n15783 = n15781 | n15782 ;
  assign n15784 = x112 & n4795 ;
  assign n15785 = n15783 | n15784 ;
  assign n15786 = ( ~x44 & n15779 ) | ( ~x44 & n15785 ) | ( n15779 & n15785 ) ;
  assign n15787 = x44 & ~n15785 ;
  assign n15788 = ( ~n15780 & n15786 ) | ( ~n15780 & n15787 ) | ( n15786 & n15787 ) ;
  assign n15789 = n5223 & n5347 ;
  assign n15790 = x47 & n15789 ;
  assign n15791 = x111 & n5230 ;
  assign n15792 = x110 & n5227 ;
  assign n15793 = n15791 | n15792 ;
  assign n15794 = x109 & n5434 ;
  assign n15795 = n15793 | n15794 ;
  assign n15796 = ( ~x47 & n15789 ) | ( ~x47 & n15795 ) | ( n15789 & n15795 ) ;
  assign n15797 = x47 & ~n15795 ;
  assign n15798 = ( ~n15790 & n15796 ) | ( ~n15790 & n15797 ) | ( n15796 & n15797 ) ;
  assign n15799 = n4914 & n5858 ;
  assign n15800 = x50 & n15799 ;
  assign n15801 = x108 & n5865 ;
  assign n15802 = x107 & n5862 ;
  assign n15803 = n15801 | n15802 ;
  assign n15804 = x106 & n6092 ;
  assign n15805 = n15803 | n15804 ;
  assign n15806 = ( ~x50 & n15799 ) | ( ~x50 & n15805 ) | ( n15799 & n15805 ) ;
  assign n15807 = x50 & ~n15805 ;
  assign n15808 = ( ~n15800 & n15806 ) | ( ~n15800 & n15807 ) | ( n15806 & n15807 ) ;
  assign n15809 = n4145 & n6546 ;
  assign n15810 = x53 & n15809 ;
  assign n15811 = x105 & n6553 ;
  assign n15812 = x104 & n6550 ;
  assign n15813 = n15811 | n15812 ;
  assign n15814 = x103 & n6787 ;
  assign n15815 = n15813 | n15814 ;
  assign n15816 = ( ~x53 & n15809 ) | ( ~x53 & n15815 ) | ( n15809 & n15815 ) ;
  assign n15817 = x53 & ~n15815 ;
  assign n15818 = ( ~n15810 & n15816 ) | ( ~n15810 & n15817 ) | ( n15816 & n15817 ) ;
  assign n15819 = n3764 & n7277 ;
  assign n15820 = x56 & n15819 ;
  assign n15821 = x102 & n7545 ;
  assign n15822 = x101 & n7273 ;
  assign n15823 = n15821 | n15822 ;
  assign n15824 = x100 & n7552 ;
  assign n15825 = n15823 | n15824 ;
  assign n15826 = ( ~x56 & n15819 ) | ( ~x56 & n15825 ) | ( n15819 & n15825 ) ;
  assign n15827 = x56 & ~n15825 ;
  assign n15828 = ( ~n15820 & n15826 ) | ( ~n15820 & n15827 ) | ( n15826 & n15827 ) ;
  assign n15829 = n3248 & n8067 ;
  assign n15830 = x59 & n15829 ;
  assign n15831 = x99 & n8074 ;
  assign n15832 = x98 & n8071 ;
  assign n15833 = n15831 | n15832 ;
  assign n15834 = x97 & n8298 ;
  assign n15835 = n15833 | n15834 ;
  assign n15836 = ( ~x59 & n15829 ) | ( ~x59 & n15835 ) | ( n15829 & n15835 ) ;
  assign n15837 = x59 & ~n15835 ;
  assign n15838 = ( ~n15830 & n15836 ) | ( ~n15830 & n15837 ) | ( n15836 & n15837 ) ;
  assign n15839 = n2772 & n8859 ;
  assign n15840 = x62 & n15839 ;
  assign n15841 = x96 & n8866 ;
  assign n15842 = x95 & n8863 ;
  assign n15843 = n15841 | n15842 ;
  assign n15844 = x94 & n9125 ;
  assign n15845 = n15843 | n15844 ;
  assign n15846 = ( ~x62 & n15839 ) | ( ~x62 & n15845 ) | ( n15839 & n15845 ) ;
  assign n15847 = x62 & ~n15845 ;
  assign n15848 = ( ~n15840 & n15846 ) | ( ~n15840 & n15847 ) | ( n15846 & n15847 ) ;
  assign n15849 = ( x62 & x63 ) | ( x62 & x93 ) | ( x63 & x93 ) ;
  assign n15850 = ( x62 & x92 ) | ( x62 & ~n9394 ) | ( x92 & ~n9394 ) ;
  assign n15851 = ( x92 & n15849 ) | ( x92 & ~n15850 ) | ( n15849 & ~n15850 ) ;
  assign n15852 = ( n15689 & ~n15691 ) | ( n15689 & n15851 ) | ( ~n15691 & n15851 ) ;
  assign n15853 = ( n15528 & n15690 ) | ( n15528 & ~n15851 ) | ( n15690 & ~n15851 ) ;
  assign n15854 = ( ~n15689 & n15852 ) | ( ~n15689 & n15853 ) | ( n15852 & n15853 ) ;
  assign n15855 = ( n15838 & ~n15848 ) | ( n15838 & n15854 ) | ( ~n15848 & n15854 ) ;
  assign n15856 = ( n15838 & n15848 ) | ( n15838 & ~n15854 ) | ( n15848 & ~n15854 ) ;
  assign n15857 = ( ~n15838 & n15855 ) | ( ~n15838 & n15856 ) | ( n15855 & n15856 ) ;
  assign n15858 = ( n15693 & n15828 ) | ( n15693 & ~n15857 ) | ( n15828 & ~n15857 ) ;
  assign n15859 = ( ~n15693 & n15828 ) | ( ~n15693 & n15857 ) | ( n15828 & n15857 ) ;
  assign n15860 = ( ~n15828 & n15858 ) | ( ~n15828 & n15859 ) | ( n15858 & n15859 ) ;
  assign n15861 = ( n15696 & n15818 ) | ( n15696 & ~n15860 ) | ( n15818 & ~n15860 ) ;
  assign n15862 = ( ~n15696 & n15818 ) | ( ~n15696 & n15860 ) | ( n15818 & n15860 ) ;
  assign n15863 = ( ~n15818 & n15861 ) | ( ~n15818 & n15862 ) | ( n15861 & n15862 ) ;
  assign n15864 = ( ~n15699 & n15808 ) | ( ~n15699 & n15863 ) | ( n15808 & n15863 ) ;
  assign n15865 = ( n15699 & n15808 ) | ( n15699 & ~n15863 ) | ( n15808 & ~n15863 ) ;
  assign n15866 = ( ~n15808 & n15864 ) | ( ~n15808 & n15865 ) | ( n15864 & n15865 ) ;
  assign n15867 = ( n15702 & n15798 ) | ( n15702 & ~n15866 ) | ( n15798 & ~n15866 ) ;
  assign n15868 = ( ~n15702 & n15798 ) | ( ~n15702 & n15866 ) | ( n15798 & n15866 ) ;
  assign n15869 = ( ~n15798 & n15867 ) | ( ~n15798 & n15868 ) | ( n15867 & n15868 ) ;
  assign n15870 = ( n15706 & n15788 ) | ( n15706 & ~n15869 ) | ( n15788 & ~n15869 ) ;
  assign n15871 = ( ~n15706 & n15788 ) | ( ~n15706 & n15869 ) | ( n15788 & n15869 ) ;
  assign n15872 = ( ~n15788 & n15870 ) | ( ~n15788 & n15871 ) | ( n15870 & n15871 ) ;
  assign n15873 = ( ~n15708 & n15778 ) | ( ~n15708 & n15872 ) | ( n15778 & n15872 ) ;
  assign n15874 = ( n15708 & n15778 ) | ( n15708 & ~n15872 ) | ( n15778 & ~n15872 ) ;
  assign n15875 = ( ~n15778 & n15873 ) | ( ~n15778 & n15874 ) | ( n15873 & n15874 ) ;
  assign n15876 = ( n15721 & n15768 ) | ( n15721 & ~n15875 ) | ( n15768 & ~n15875 ) ;
  assign n15877 = ( ~n15721 & n15768 ) | ( ~n15721 & n15875 ) | ( n15768 & n15875 ) ;
  assign n15878 = ( ~n15768 & n15876 ) | ( ~n15768 & n15877 ) | ( n15876 & n15877 ) ;
  assign n15879 = ( ~n15724 & n15758 ) | ( ~n15724 & n15878 ) | ( n15758 & n15878 ) ;
  assign n15880 = ( n15724 & n15758 ) | ( n15724 & ~n15878 ) | ( n15758 & ~n15878 ) ;
  assign n15881 = ( ~n15758 & n15879 ) | ( ~n15758 & n15880 ) | ( n15879 & n15880 ) ;
  assign n15882 = ( n15727 & n15748 ) | ( n15727 & ~n15881 ) | ( n15748 & ~n15881 ) ;
  assign n15883 = ( ~n15727 & n15748 ) | ( ~n15727 & n15881 ) | ( n15748 & n15881 ) ;
  assign n15884 = ( ~n15748 & n15882 ) | ( ~n15748 & n15883 ) | ( n15882 & n15883 ) ;
  assign n15885 = x127 & n2267 ;
  assign n15886 = n2137 | n15885 ;
  assign n15887 = ( n9865 & n15885 ) | ( n9865 & n15886 ) | ( n15885 & n15886 ) ;
  assign n15888 = x29 & ~n15887 ;
  assign n15889 = ~x29 & n15887 ;
  assign n15890 = n15888 | n15889 ;
  assign n15891 = ( n15730 & n15884 ) | ( n15730 & n15890 ) | ( n15884 & n15890 ) ;
  assign n15892 = ( n15730 & ~n15884 ) | ( n15730 & n15890 ) | ( ~n15884 & n15890 ) ;
  assign n15893 = ( n15884 & ~n15891 ) | ( n15884 & n15892 ) | ( ~n15891 & n15892 ) ;
  assign n15894 = ( ~n15733 & n15736 ) | ( ~n15733 & n15893 ) | ( n15736 & n15893 ) ;
  assign n15895 = ( n15733 & n15736 ) | ( n15733 & ~n15893 ) | ( n15736 & ~n15893 ) ;
  assign n15896 = ( ~n15736 & n15894 ) | ( ~n15736 & n15895 ) | ( n15894 & n15895 ) ;
  assign n15897 = n2545 & n9576 ;
  assign n15898 = x32 & n15897 ;
  assign n15899 = x127 & n2552 ;
  assign n15900 = x126 & n2549 ;
  assign n15901 = n15899 | n15900 ;
  assign n15902 = x125 & n2696 ;
  assign n15903 = n15901 | n15902 ;
  assign n15904 = ( ~x32 & n15897 ) | ( ~x32 & n15903 ) | ( n15897 & n15903 ) ;
  assign n15905 = x32 & ~n15903 ;
  assign n15906 = ( ~n15898 & n15904 ) | ( ~n15898 & n15905 ) | ( n15904 & n15905 ) ;
  assign n15907 = n2982 & n8729 ;
  assign n15908 = x35 & n15907 ;
  assign n15909 = x124 & n2989 ;
  assign n15910 = x123 & n2986 ;
  assign n15911 = n15909 | n15910 ;
  assign n15912 = x122 & n3159 ;
  assign n15913 = n15911 | n15912 ;
  assign n15914 = ( ~x35 & n15907 ) | ( ~x35 & n15913 ) | ( n15907 & n15913 ) ;
  assign n15915 = x35 & ~n15913 ;
  assign n15916 = ( ~n15908 & n15914 ) | ( ~n15908 & n15915 ) | ( n15914 & n15915 ) ;
  assign n15917 = n3492 & n7696 ;
  assign n15918 = x38 & n15917 ;
  assign n15919 = x121 & n3499 ;
  assign n15920 = x120 & n3496 ;
  assign n15921 = n15919 | n15920 ;
  assign n15922 = x119 & n3662 ;
  assign n15923 = n15921 | n15922 ;
  assign n15924 = ( ~x38 & n15917 ) | ( ~x38 & n15923 ) | ( n15917 & n15923 ) ;
  assign n15925 = x38 & ~n15923 ;
  assign n15926 = ( ~n15918 & n15924 ) | ( ~n15918 & n15925 ) | ( n15924 & n15925 ) ;
  assign n15927 = n4020 & n6940 ;
  assign n15928 = x41 & n15927 ;
  assign n15929 = x118 & n4027 ;
  assign n15930 = x117 & n4024 ;
  assign n15931 = n15929 | n15930 ;
  assign n15932 = x116 & n4223 ;
  assign n15933 = n15931 | n15932 ;
  assign n15934 = ( ~x41 & n15927 ) | ( ~x41 & n15933 ) | ( n15927 & n15933 ) ;
  assign n15935 = x41 & ~n15933 ;
  assign n15936 = ( ~n15928 & n15934 ) | ( ~n15928 & n15935 ) | ( n15934 & n15935 ) ;
  assign n15937 = n4625 & n6446 ;
  assign n15938 = x44 & n15937 ;
  assign n15939 = x115 & n4791 ;
  assign n15940 = x114 & n4621 ;
  assign n15941 = n15939 | n15940 ;
  assign n15942 = x113 & n4795 ;
  assign n15943 = n15941 | n15942 ;
  assign n15944 = ( ~x44 & n15937 ) | ( ~x44 & n15943 ) | ( n15937 & n15943 ) ;
  assign n15945 = x44 & ~n15943 ;
  assign n15946 = ( ~n15938 & n15944 ) | ( ~n15938 & n15945 ) | ( n15944 & n15945 ) ;
  assign n15947 = n5223 & n5558 ;
  assign n15948 = x47 & n15947 ;
  assign n15949 = x112 & n5230 ;
  assign n15950 = x111 & n5227 ;
  assign n15951 = n15949 | n15950 ;
  assign n15952 = x110 & n5434 ;
  assign n15953 = n15951 | n15952 ;
  assign n15954 = ( ~x47 & n15947 ) | ( ~x47 & n15953 ) | ( n15947 & n15953 ) ;
  assign n15955 = x47 & ~n15953 ;
  assign n15956 = ( ~n15948 & n15954 ) | ( ~n15948 & n15955 ) | ( n15954 & n15955 ) ;
  assign n15957 = n4930 & n5858 ;
  assign n15958 = x50 & n15957 ;
  assign n15959 = x109 & n5865 ;
  assign n15960 = x108 & n5862 ;
  assign n15961 = n15959 | n15960 ;
  assign n15962 = x107 & n6092 ;
  assign n15963 = n15961 | n15962 ;
  assign n15964 = ( ~x50 & n15957 ) | ( ~x50 & n15963 ) | ( n15957 & n15963 ) ;
  assign n15965 = x50 & ~n15963 ;
  assign n15966 = ( ~n15958 & n15964 ) | ( ~n15958 & n15965 ) | ( n15964 & n15965 ) ;
  assign n15967 = n3941 & n7277 ;
  assign n15968 = x56 & n15967 ;
  assign n15969 = x103 & n7545 ;
  assign n15970 = x102 & n7273 ;
  assign n15971 = n15969 | n15970 ;
  assign n15972 = x101 & n7552 ;
  assign n15973 = n15971 | n15972 ;
  assign n15974 = ( ~x56 & n15967 ) | ( ~x56 & n15973 ) | ( n15967 & n15973 ) ;
  assign n15975 = x56 & ~n15973 ;
  assign n15976 = ( ~n15968 & n15974 ) | ( ~n15968 & n15975 ) | ( n15974 & n15975 ) ;
  assign n15977 = n3264 & n8067 ;
  assign n15978 = x59 & n15977 ;
  assign n15979 = x100 & n8074 ;
  assign n15980 = x99 & n8071 ;
  assign n15981 = n15979 | n15980 ;
  assign n15982 = x98 & n8298 ;
  assign n15983 = n15981 | n15982 ;
  assign n15984 = ( ~x59 & n15977 ) | ( ~x59 & n15983 ) | ( n15977 & n15983 ) ;
  assign n15985 = x59 & ~n15983 ;
  assign n15986 = ( ~n15978 & n15984 ) | ( ~n15978 & n15985 ) | ( n15984 & n15985 ) ;
  assign n15987 = n2788 & n8859 ;
  assign n15988 = x62 & n15987 ;
  assign n15989 = x97 & n8866 ;
  assign n15990 = x96 & n8863 ;
  assign n15991 = n15989 | n15990 ;
  assign n15992 = x95 & n9125 ;
  assign n15993 = n15991 | n15992 ;
  assign n15994 = ( ~x62 & n15987 ) | ( ~x62 & n15993 ) | ( n15987 & n15993 ) ;
  assign n15995 = x62 & ~n15993 ;
  assign n15996 = ( ~n15988 & n15994 ) | ( ~n15988 & n15995 ) | ( n15994 & n15995 ) ;
  assign n15997 = ( x62 & x63 ) | ( x62 & x94 ) | ( x63 & x94 ) ;
  assign n15998 = ( x62 & x93 ) | ( x62 & ~n9394 ) | ( x93 & ~n9394 ) ;
  assign n15999 = ( x93 & n15997 ) | ( x93 & ~n15998 ) | ( n15997 & ~n15998 ) ;
  assign n16000 = ( x29 & n15851 ) | ( x29 & n15999 ) | ( n15851 & n15999 ) ;
  assign n16001 = ( ~x29 & n15851 ) | ( ~x29 & n15999 ) | ( n15851 & n15999 ) ;
  assign n16002 = ( x29 & ~n16000 ) | ( x29 & n16001 ) | ( ~n16000 & n16001 ) ;
  assign n16003 = ( n15853 & n15996 ) | ( n15853 & ~n16002 ) | ( n15996 & ~n16002 ) ;
  assign n16004 = ( ~n15853 & n15996 ) | ( ~n15853 & n16002 ) | ( n15996 & n16002 ) ;
  assign n16005 = ( ~n15996 & n16003 ) | ( ~n15996 & n16004 ) | ( n16003 & n16004 ) ;
  assign n16006 = ( n15856 & n15986 ) | ( n15856 & ~n16005 ) | ( n15986 & ~n16005 ) ;
  assign n16007 = ( n15856 & ~n15986 ) | ( n15856 & n16005 ) | ( ~n15986 & n16005 ) ;
  assign n16008 = ( ~n15856 & n16006 ) | ( ~n15856 & n16007 ) | ( n16006 & n16007 ) ;
  assign n16009 = ( n15858 & ~n15976 ) | ( n15858 & n16008 ) | ( ~n15976 & n16008 ) ;
  assign n16010 = ( n15858 & n15976 ) | ( n15858 & ~n16008 ) | ( n15976 & ~n16008 ) ;
  assign n16011 = ( ~n15858 & n16009 ) | ( ~n15858 & n16010 ) | ( n16009 & n16010 ) ;
  assign n16012 = n4331 & n6546 ;
  assign n16013 = x53 & n16012 ;
  assign n16014 = x106 & n6553 ;
  assign n16015 = x105 & n6550 ;
  assign n16016 = n16014 | n16015 ;
  assign n16017 = x104 & n6787 ;
  assign n16018 = n16016 | n16017 ;
  assign n16019 = ( ~x53 & n16012 ) | ( ~x53 & n16018 ) | ( n16012 & n16018 ) ;
  assign n16020 = x53 & ~n16018 ;
  assign n16021 = ( ~n16013 & n16019 ) | ( ~n16013 & n16020 ) | ( n16019 & n16020 ) ;
  assign n16022 = ( n15861 & n16011 ) | ( n15861 & ~n16021 ) | ( n16011 & ~n16021 ) ;
  assign n16023 = ( n15861 & ~n16011 ) | ( n15861 & n16021 ) | ( ~n16011 & n16021 ) ;
  assign n16024 = ( ~n15861 & n16022 ) | ( ~n15861 & n16023 ) | ( n16022 & n16023 ) ;
  assign n16025 = ( n15865 & n15966 ) | ( n15865 & ~n16024 ) | ( n15966 & ~n16024 ) ;
  assign n16026 = ( n15865 & ~n15966 ) | ( n15865 & n16024 ) | ( ~n15966 & n16024 ) ;
  assign n16027 = ( ~n15865 & n16025 ) | ( ~n15865 & n16026 ) | ( n16025 & n16026 ) ;
  assign n16028 = ( n15867 & n15956 ) | ( n15867 & ~n16027 ) | ( n15956 & ~n16027 ) ;
  assign n16029 = ( n15867 & ~n15956 ) | ( n15867 & n16027 ) | ( ~n15956 & n16027 ) ;
  assign n16030 = ( ~n15867 & n16028 ) | ( ~n15867 & n16029 ) | ( n16028 & n16029 ) ;
  assign n16031 = ( n15870 & n15946 ) | ( n15870 & ~n16030 ) | ( n15946 & ~n16030 ) ;
  assign n16032 = ( n15870 & ~n15946 ) | ( n15870 & n16030 ) | ( ~n15946 & n16030 ) ;
  assign n16033 = ( ~n15870 & n16031 ) | ( ~n15870 & n16032 ) | ( n16031 & n16032 ) ;
  assign n16034 = ( n15874 & n15936 ) | ( n15874 & ~n16033 ) | ( n15936 & ~n16033 ) ;
  assign n16035 = ( n15874 & ~n15936 ) | ( n15874 & n16033 ) | ( ~n15936 & n16033 ) ;
  assign n16036 = ( ~n15874 & n16034 ) | ( ~n15874 & n16035 ) | ( n16034 & n16035 ) ;
  assign n16037 = ( n15876 & n15926 ) | ( n15876 & ~n16036 ) | ( n15926 & ~n16036 ) ;
  assign n16038 = ( n15876 & ~n15926 ) | ( n15876 & n16036 ) | ( ~n15926 & n16036 ) ;
  assign n16039 = ( ~n15876 & n16037 ) | ( ~n15876 & n16038 ) | ( n16037 & n16038 ) ;
  assign n16040 = ( n15880 & n15916 ) | ( n15880 & ~n16039 ) | ( n15916 & ~n16039 ) ;
  assign n16041 = ( n15880 & ~n15916 ) | ( n15880 & n16039 ) | ( ~n15916 & n16039 ) ;
  assign n16042 = ( ~n15880 & n16040 ) | ( ~n15880 & n16041 ) | ( n16040 & n16041 ) ;
  assign n16043 = ( n15882 & n15906 ) | ( n15882 & ~n16042 ) | ( n15906 & ~n16042 ) ;
  assign n16044 = ( n15882 & ~n15906 ) | ( n15882 & n16042 ) | ( ~n15906 & n16042 ) ;
  assign n16045 = ( ~n15882 & n16043 ) | ( ~n15882 & n16044 ) | ( n16043 & n16044 ) ;
  assign n16046 = ( ~n15892 & n15894 ) | ( ~n15892 & n16045 ) | ( n15894 & n16045 ) ;
  assign n16047 = ( n15892 & n15894 ) | ( n15892 & ~n16045 ) | ( n15894 & ~n16045 ) ;
  assign n16048 = ( ~n15894 & n16046 ) | ( ~n15894 & n16047 ) | ( n16046 & n16047 ) ;
  assign n16049 = x127 & n2549 ;
  assign n16050 = n2545 | n16049 ;
  assign n16051 = ( n9867 & n16049 ) | ( n9867 & n16050 ) | ( n16049 & n16050 ) ;
  assign n16052 = x126 & n2696 ;
  assign n16053 = ( ~x32 & n16051 ) | ( ~x32 & n16052 ) | ( n16051 & n16052 ) ;
  assign n16054 = ( x32 & ~n16051 ) | ( x32 & n16052 ) | ( ~n16051 & n16052 ) ;
  assign n16055 = ~n16052 & n16054 ;
  assign n16056 = n16053 | n16055 ;
  assign n16057 = n2982 & n9009 ;
  assign n16058 = x35 & n16057 ;
  assign n16059 = x125 & n2989 ;
  assign n16060 = x124 & n2986 ;
  assign n16061 = n16059 | n16060 ;
  assign n16062 = x123 & n3159 ;
  assign n16063 = n16061 | n16062 ;
  assign n16064 = ( ~x35 & n16057 ) | ( ~x35 & n16063 ) | ( n16057 & n16063 ) ;
  assign n16065 = x35 & ~n16063 ;
  assign n16066 = ( ~n16058 & n16064 ) | ( ~n16058 & n16065 ) | ( n16064 & n16065 ) ;
  assign n16067 = n3492 & n8207 ;
  assign n16068 = x38 & n16067 ;
  assign n16069 = x122 & n3499 ;
  assign n16070 = x121 & n3496 ;
  assign n16071 = n16069 | n16070 ;
  assign n16072 = x120 & n3662 ;
  assign n16073 = n16071 | n16072 ;
  assign n16074 = ( ~x38 & n16067 ) | ( ~x38 & n16073 ) | ( n16067 & n16073 ) ;
  assign n16075 = x38 & ~n16073 ;
  assign n16076 = ( ~n16068 & n16074 ) | ( ~n16068 & n16075 ) | ( n16074 & n16075 ) ;
  assign n16077 = n4020 & n7181 ;
  assign n16078 = x41 & n16077 ;
  assign n16079 = x119 & n4027 ;
  assign n16080 = x118 & n4024 ;
  assign n16081 = n16079 | n16080 ;
  assign n16082 = x117 & n4223 ;
  assign n16083 = n16081 | n16082 ;
  assign n16084 = ( ~x41 & n16077 ) | ( ~x41 & n16083 ) | ( n16077 & n16083 ) ;
  assign n16085 = x41 & ~n16083 ;
  assign n16086 = ( ~n16078 & n16084 ) | ( ~n16078 & n16085 ) | ( n16084 & n16085 ) ;
  assign n16087 = n4625 & n6462 ;
  assign n16088 = x44 & n16087 ;
  assign n16089 = x116 & n4791 ;
  assign n16090 = x115 & n4621 ;
  assign n16091 = n16089 | n16090 ;
  assign n16092 = x114 & n4795 ;
  assign n16093 = n16091 | n16092 ;
  assign n16094 = ( ~x44 & n16087 ) | ( ~x44 & n16093 ) | ( n16087 & n16093 ) ;
  assign n16095 = x44 & ~n16093 ;
  assign n16096 = ( ~n16088 & n16094 ) | ( ~n16088 & n16095 ) | ( n16094 & n16095 ) ;
  assign n16097 = n5223 & n5774 ;
  assign n16098 = x47 & n16097 ;
  assign n16099 = x113 & n5230 ;
  assign n16100 = x112 & n5227 ;
  assign n16101 = n16099 | n16100 ;
  assign n16102 = x111 & n5434 ;
  assign n16103 = n16101 | n16102 ;
  assign n16104 = ( ~x47 & n16097 ) | ( ~x47 & n16103 ) | ( n16097 & n16103 ) ;
  assign n16105 = x47 & ~n16103 ;
  assign n16106 = ( ~n16098 & n16104 ) | ( ~n16098 & n16105 ) | ( n16104 & n16105 ) ;
  assign n16107 = n5331 & n5858 ;
  assign n16108 = x50 & n16107 ;
  assign n16109 = x110 & n5865 ;
  assign n16110 = x109 & n5862 ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = x108 & n6092 ;
  assign n16113 = n16111 | n16112 ;
  assign n16114 = ( ~x50 & n16107 ) | ( ~x50 & n16113 ) | ( n16107 & n16113 ) ;
  assign n16115 = x50 & ~n16113 ;
  assign n16116 = ( ~n16108 & n16114 ) | ( ~n16108 & n16115 ) | ( n16114 & n16115 ) ;
  assign n16117 = n4523 & n6546 ;
  assign n16118 = x53 & n16117 ;
  assign n16119 = x107 & n6553 ;
  assign n16120 = x106 & n6550 ;
  assign n16121 = n16119 | n16120 ;
  assign n16122 = x105 & n6787 ;
  assign n16123 = n16121 | n16122 ;
  assign n16124 = ( ~x53 & n16117 ) | ( ~x53 & n16123 ) | ( n16117 & n16123 ) ;
  assign n16125 = x53 & ~n16123 ;
  assign n16126 = ( ~n16118 & n16124 ) | ( ~n16118 & n16125 ) | ( n16124 & n16125 ) ;
  assign n16127 = n3957 & n7277 ;
  assign n16128 = x56 & n16127 ;
  assign n16129 = x104 & n7545 ;
  assign n16130 = x103 & n7273 ;
  assign n16131 = n16129 | n16130 ;
  assign n16132 = x102 & n7552 ;
  assign n16133 = n16131 | n16132 ;
  assign n16134 = ( ~x56 & n16127 ) | ( ~x56 & n16133 ) | ( n16127 & n16133 ) ;
  assign n16135 = x56 & ~n16133 ;
  assign n16136 = ( ~n16128 & n16134 ) | ( ~n16128 & n16135 ) | ( n16134 & n16135 ) ;
  assign n16137 = n3591 & n8067 ;
  assign n16138 = x59 & n16137 ;
  assign n16139 = x101 & n8074 ;
  assign n16140 = x100 & n8071 ;
  assign n16141 = n16139 | n16140 ;
  assign n16142 = x99 & n8298 ;
  assign n16143 = n16141 | n16142 ;
  assign n16144 = ( ~x59 & n16137 ) | ( ~x59 & n16143 ) | ( n16137 & n16143 ) ;
  assign n16145 = x59 & ~n16143 ;
  assign n16146 = ( ~n16138 & n16144 ) | ( ~n16138 & n16145 ) | ( n16144 & n16145 ) ;
  assign n16147 = ( x62 & x63 ) | ( x62 & x95 ) | ( x63 & x95 ) ;
  assign n16148 = ( x62 & x94 ) | ( x62 & ~n9394 ) | ( x94 & ~n9394 ) ;
  assign n16149 = ( x94 & n16147 ) | ( x94 & ~n16148 ) | ( n16147 & ~n16148 ) ;
  assign n16150 = n2939 & n8859 ;
  assign n16151 = x62 & n16150 ;
  assign n16152 = x98 & n8866 ;
  assign n16153 = x97 & n8863 ;
  assign n16154 = n16152 | n16153 ;
  assign n16155 = x96 & n9125 ;
  assign n16156 = n16154 | n16155 ;
  assign n16157 = ( ~x62 & n16150 ) | ( ~x62 & n16156 ) | ( n16150 & n16156 ) ;
  assign n16158 = x62 & ~n16156 ;
  assign n16159 = ( ~n16151 & n16157 ) | ( ~n16151 & n16158 ) | ( n16157 & n16158 ) ;
  assign n16160 = ( ~n16001 & n16149 ) | ( ~n16001 & n16159 ) | ( n16149 & n16159 ) ;
  assign n16161 = ( n16001 & n16149 ) | ( n16001 & ~n16159 ) | ( n16149 & ~n16159 ) ;
  assign n16162 = ( ~n16149 & n16160 ) | ( ~n16149 & n16161 ) | ( n16160 & n16161 ) ;
  assign n16163 = ( n16003 & n16146 ) | ( n16003 & ~n16162 ) | ( n16146 & ~n16162 ) ;
  assign n16164 = ( ~n16003 & n16146 ) | ( ~n16003 & n16162 ) | ( n16146 & n16162 ) ;
  assign n16165 = ( ~n16146 & n16163 ) | ( ~n16146 & n16164 ) | ( n16163 & n16164 ) ;
  assign n16166 = ( n16006 & n16136 ) | ( n16006 & ~n16165 ) | ( n16136 & ~n16165 ) ;
  assign n16167 = ( ~n16006 & n16136 ) | ( ~n16006 & n16165 ) | ( n16136 & n16165 ) ;
  assign n16168 = ( ~n16136 & n16166 ) | ( ~n16136 & n16167 ) | ( n16166 & n16167 ) ;
  assign n16169 = ( n16010 & n16126 ) | ( n16010 & ~n16168 ) | ( n16126 & ~n16168 ) ;
  assign n16170 = ( ~n16010 & n16126 ) | ( ~n16010 & n16168 ) | ( n16126 & n16168 ) ;
  assign n16171 = ( ~n16126 & n16169 ) | ( ~n16126 & n16170 ) | ( n16169 & n16170 ) ;
  assign n16172 = ( n16023 & n16116 ) | ( n16023 & ~n16171 ) | ( n16116 & ~n16171 ) ;
  assign n16173 = ( ~n16023 & n16116 ) | ( ~n16023 & n16171 ) | ( n16116 & n16171 ) ;
  assign n16174 = ( ~n16116 & n16172 ) | ( ~n16116 & n16173 ) | ( n16172 & n16173 ) ;
  assign n16175 = ( n16025 & n16106 ) | ( n16025 & ~n16174 ) | ( n16106 & ~n16174 ) ;
  assign n16176 = ( ~n16025 & n16106 ) | ( ~n16025 & n16174 ) | ( n16106 & n16174 ) ;
  assign n16177 = ( ~n16106 & n16175 ) | ( ~n16106 & n16176 ) | ( n16175 & n16176 ) ;
  assign n16178 = ( n16028 & n16096 ) | ( n16028 & ~n16177 ) | ( n16096 & ~n16177 ) ;
  assign n16179 = ( ~n16028 & n16096 ) | ( ~n16028 & n16177 ) | ( n16096 & n16177 ) ;
  assign n16180 = ( ~n16096 & n16178 ) | ( ~n16096 & n16179 ) | ( n16178 & n16179 ) ;
  assign n16181 = ( n16031 & n16086 ) | ( n16031 & ~n16180 ) | ( n16086 & ~n16180 ) ;
  assign n16182 = ( ~n16031 & n16086 ) | ( ~n16031 & n16180 ) | ( n16086 & n16180 ) ;
  assign n16183 = ( ~n16086 & n16181 ) | ( ~n16086 & n16182 ) | ( n16181 & n16182 ) ;
  assign n16184 = ( n16034 & n16076 ) | ( n16034 & ~n16183 ) | ( n16076 & ~n16183 ) ;
  assign n16185 = ( ~n16034 & n16076 ) | ( ~n16034 & n16183 ) | ( n16076 & n16183 ) ;
  assign n16186 = ( ~n16076 & n16184 ) | ( ~n16076 & n16185 ) | ( n16184 & n16185 ) ;
  assign n16187 = ( n16037 & n16066 ) | ( n16037 & ~n16186 ) | ( n16066 & ~n16186 ) ;
  assign n16188 = ( ~n16037 & n16066 ) | ( ~n16037 & n16186 ) | ( n16066 & n16186 ) ;
  assign n16189 = ( ~n16066 & n16187 ) | ( ~n16066 & n16188 ) | ( n16187 & n16188 ) ;
  assign n16190 = ( n16040 & n16056 ) | ( n16040 & ~n16189 ) | ( n16056 & ~n16189 ) ;
  assign n16191 = ( ~n16040 & n16056 ) | ( ~n16040 & n16189 ) | ( n16056 & n16189 ) ;
  assign n16192 = ( ~n16056 & n16190 ) | ( ~n16056 & n16191 ) | ( n16190 & n16191 ) ;
  assign n16193 = ( ~n16043 & n16046 ) | ( ~n16043 & n16192 ) | ( n16046 & n16192 ) ;
  assign n16194 = ( n16043 & n16046 ) | ( n16043 & ~n16192 ) | ( n16046 & ~n16192 ) ;
  assign n16195 = ( ~n16046 & n16193 ) | ( ~n16046 & n16194 ) | ( n16193 & n16194 ) ;
  assign n16196 = n2982 & n9038 ;
  assign n16197 = x35 & n16196 ;
  assign n16198 = x126 & n2989 ;
  assign n16199 = x125 & n2986 ;
  assign n16200 = n16198 | n16199 ;
  assign n16201 = x124 & n3159 ;
  assign n16202 = n16200 | n16201 ;
  assign n16203 = ( ~x35 & n16196 ) | ( ~x35 & n16202 ) | ( n16196 & n16202 ) ;
  assign n16204 = x35 & ~n16202 ;
  assign n16205 = ( ~n16197 & n16203 ) | ( ~n16197 & n16204 ) | ( n16203 & n16204 ) ;
  assign n16206 = n3492 & n8461 ;
  assign n16207 = x38 & n16206 ;
  assign n16208 = x123 & n3499 ;
  assign n16209 = x122 & n3496 ;
  assign n16210 = n16208 | n16209 ;
  assign n16211 = x121 & n3662 ;
  assign n16212 = n16210 | n16211 ;
  assign n16213 = ( ~x38 & n16206 ) | ( ~x38 & n16212 ) | ( n16206 & n16212 ) ;
  assign n16214 = x38 & ~n16212 ;
  assign n16215 = ( ~n16207 & n16213 ) | ( ~n16207 & n16214 ) | ( n16213 & n16214 ) ;
  assign n16216 = n4020 & n7444 ;
  assign n16217 = x41 & n16216 ;
  assign n16218 = x120 & n4027 ;
  assign n16219 = x119 & n4024 ;
  assign n16220 = n16218 | n16219 ;
  assign n16221 = x118 & n4223 ;
  assign n16222 = n16220 | n16221 ;
  assign n16223 = ( ~x41 & n16216 ) | ( ~x41 & n16222 ) | ( n16216 & n16222 ) ;
  assign n16224 = x41 & ~n16222 ;
  assign n16225 = ( ~n16217 & n16223 ) | ( ~n16217 & n16224 ) | ( n16223 & n16224 ) ;
  assign n16226 = n4625 & n6924 ;
  assign n16227 = x44 & n16226 ;
  assign n16228 = x117 & n4791 ;
  assign n16229 = x116 & n4621 ;
  assign n16230 = n16228 | n16229 ;
  assign n16231 = x115 & n4795 ;
  assign n16232 = n16230 | n16231 ;
  assign n16233 = ( ~x44 & n16226 ) | ( ~x44 & n16232 ) | ( n16226 & n16232 ) ;
  assign n16234 = x44 & ~n16232 ;
  assign n16235 = ( ~n16227 & n16233 ) | ( ~n16227 & n16234 ) | ( n16233 & n16234 ) ;
  assign n16236 = n5223 & n6002 ;
  assign n16237 = x47 & n16236 ;
  assign n16238 = x114 & n5230 ;
  assign n16239 = x113 & n5227 ;
  assign n16240 = n16238 | n16239 ;
  assign n16241 = x112 & n5434 ;
  assign n16242 = n16240 | n16241 ;
  assign n16243 = ( ~x47 & n16236 ) | ( ~x47 & n16242 ) | ( n16236 & n16242 ) ;
  assign n16244 = x47 & ~n16242 ;
  assign n16245 = ( ~n16237 & n16243 ) | ( ~n16237 & n16244 ) | ( n16243 & n16244 ) ;
  assign n16246 = n5347 & n5858 ;
  assign n16247 = x50 & n16246 ;
  assign n16248 = x111 & n5865 ;
  assign n16249 = x110 & n5862 ;
  assign n16250 = n16248 | n16249 ;
  assign n16251 = x109 & n6092 ;
  assign n16252 = n16250 | n16251 ;
  assign n16253 = ( ~x50 & n16246 ) | ( ~x50 & n16252 ) | ( n16246 & n16252 ) ;
  assign n16254 = x50 & ~n16252 ;
  assign n16255 = ( ~n16247 & n16253 ) | ( ~n16247 & n16254 ) | ( n16253 & n16254 ) ;
  assign n16256 = n4914 & n6546 ;
  assign n16257 = x53 & n16256 ;
  assign n16258 = x108 & n6553 ;
  assign n16259 = x107 & n6550 ;
  assign n16260 = n16258 | n16259 ;
  assign n16261 = x106 & n6787 ;
  assign n16262 = n16260 | n16261 ;
  assign n16263 = ( ~x53 & n16256 ) | ( ~x53 & n16262 ) | ( n16256 & n16262 ) ;
  assign n16264 = x53 & ~n16262 ;
  assign n16265 = ( ~n16257 & n16263 ) | ( ~n16257 & n16264 ) | ( n16263 & n16264 ) ;
  assign n16266 = n4145 & n7277 ;
  assign n16267 = x56 & n16266 ;
  assign n16268 = x105 & n7545 ;
  assign n16269 = x104 & n7273 ;
  assign n16270 = n16268 | n16269 ;
  assign n16271 = x103 & n7552 ;
  assign n16272 = n16270 | n16271 ;
  assign n16273 = ( ~x56 & n16266 ) | ( ~x56 & n16272 ) | ( n16266 & n16272 ) ;
  assign n16274 = x56 & ~n16272 ;
  assign n16275 = ( ~n16267 & n16273 ) | ( ~n16267 & n16274 ) | ( n16273 & n16274 ) ;
  assign n16276 = n3764 & n8067 ;
  assign n16277 = x59 & n16276 ;
  assign n16278 = x102 & n8074 ;
  assign n16279 = x101 & n8071 ;
  assign n16280 = n16278 | n16279 ;
  assign n16281 = x100 & n8298 ;
  assign n16282 = n16280 | n16281 ;
  assign n16283 = ( ~x59 & n16276 ) | ( ~x59 & n16282 ) | ( n16276 & n16282 ) ;
  assign n16284 = x59 & ~n16282 ;
  assign n16285 = ( ~n16277 & n16283 ) | ( ~n16277 & n16284 ) | ( n16283 & n16284 ) ;
  assign n16286 = n3248 & n8859 ;
  assign n16287 = x62 & n16286 ;
  assign n16288 = x99 & n8866 ;
  assign n16289 = x98 & n8863 ;
  assign n16290 = n16288 | n16289 ;
  assign n16291 = x97 & n9125 ;
  assign n16292 = n16290 | n16291 ;
  assign n16293 = ( ~x62 & n16286 ) | ( ~x62 & n16292 ) | ( n16286 & n16292 ) ;
  assign n16294 = x62 & ~n16292 ;
  assign n16295 = ( ~n16287 & n16293 ) | ( ~n16287 & n16294 ) | ( n16293 & n16294 ) ;
  assign n16296 = ( x62 & x63 ) | ( x62 & x96 ) | ( x63 & x96 ) ;
  assign n16297 = ( x62 & x95 ) | ( x62 & ~n9394 ) | ( x95 & ~n9394 ) ;
  assign n16298 = ( x95 & n16296 ) | ( x95 & ~n16297 ) | ( n16296 & ~n16297 ) ;
  assign n16299 = ( n16159 & ~n16161 ) | ( n16159 & n16298 ) | ( ~n16161 & n16298 ) ;
  assign n16300 = ( n16001 & n16160 ) | ( n16001 & ~n16298 ) | ( n16160 & ~n16298 ) ;
  assign n16301 = ( ~n16159 & n16299 ) | ( ~n16159 & n16300 ) | ( n16299 & n16300 ) ;
  assign n16302 = ( n16285 & ~n16295 ) | ( n16285 & n16301 ) | ( ~n16295 & n16301 ) ;
  assign n16303 = ( n16285 & n16295 ) | ( n16285 & ~n16301 ) | ( n16295 & ~n16301 ) ;
  assign n16304 = ( ~n16285 & n16302 ) | ( ~n16285 & n16303 ) | ( n16302 & n16303 ) ;
  assign n16305 = ( n16163 & n16275 ) | ( n16163 & ~n16304 ) | ( n16275 & ~n16304 ) ;
  assign n16306 = ( ~n16163 & n16275 ) | ( ~n16163 & n16304 ) | ( n16275 & n16304 ) ;
  assign n16307 = ( ~n16275 & n16305 ) | ( ~n16275 & n16306 ) | ( n16305 & n16306 ) ;
  assign n16308 = ( n16166 & n16265 ) | ( n16166 & ~n16307 ) | ( n16265 & ~n16307 ) ;
  assign n16309 = ( ~n16166 & n16265 ) | ( ~n16166 & n16307 ) | ( n16265 & n16307 ) ;
  assign n16310 = ( ~n16265 & n16308 ) | ( ~n16265 & n16309 ) | ( n16308 & n16309 ) ;
  assign n16311 = ( n16169 & n16255 ) | ( n16169 & ~n16310 ) | ( n16255 & ~n16310 ) ;
  assign n16312 = ( ~n16169 & n16255 ) | ( ~n16169 & n16310 ) | ( n16255 & n16310 ) ;
  assign n16313 = ( ~n16255 & n16311 ) | ( ~n16255 & n16312 ) | ( n16311 & n16312 ) ;
  assign n16314 = ( ~n16172 & n16245 ) | ( ~n16172 & n16313 ) | ( n16245 & n16313 ) ;
  assign n16315 = ( n16172 & n16245 ) | ( n16172 & ~n16313 ) | ( n16245 & ~n16313 ) ;
  assign n16316 = ( ~n16245 & n16314 ) | ( ~n16245 & n16315 ) | ( n16314 & n16315 ) ;
  assign n16317 = ( n16175 & n16235 ) | ( n16175 & ~n16316 ) | ( n16235 & ~n16316 ) ;
  assign n16318 = ( ~n16175 & n16235 ) | ( ~n16175 & n16316 ) | ( n16235 & n16316 ) ;
  assign n16319 = ( ~n16235 & n16317 ) | ( ~n16235 & n16318 ) | ( n16317 & n16318 ) ;
  assign n16320 = ( n16178 & n16225 ) | ( n16178 & ~n16319 ) | ( n16225 & ~n16319 ) ;
  assign n16321 = ( ~n16178 & n16225 ) | ( ~n16178 & n16319 ) | ( n16225 & n16319 ) ;
  assign n16322 = ( ~n16225 & n16320 ) | ( ~n16225 & n16321 ) | ( n16320 & n16321 ) ;
  assign n16323 = ( n16181 & n16215 ) | ( n16181 & ~n16322 ) | ( n16215 & ~n16322 ) ;
  assign n16324 = ( ~n16181 & n16215 ) | ( ~n16181 & n16322 ) | ( n16215 & n16322 ) ;
  assign n16325 = ( ~n16215 & n16323 ) | ( ~n16215 & n16324 ) | ( n16323 & n16324 ) ;
  assign n16326 = ( n16184 & n16205 ) | ( n16184 & ~n16325 ) | ( n16205 & ~n16325 ) ;
  assign n16327 = ( ~n16184 & n16205 ) | ( ~n16184 & n16325 ) | ( n16205 & n16325 ) ;
  assign n16328 = ( ~n16205 & n16326 ) | ( ~n16205 & n16327 ) | ( n16326 & n16327 ) ;
  assign n16329 = x127 & n2696 ;
  assign n16330 = n2545 | n16329 ;
  assign n16331 = ( n9865 & n16329 ) | ( n9865 & n16330 ) | ( n16329 & n16330 ) ;
  assign n16332 = x32 & ~n16331 ;
  assign n16333 = ~x32 & n16331 ;
  assign n16334 = n16332 | n16333 ;
  assign n16335 = ( n16187 & ~n16328 ) | ( n16187 & n16334 ) | ( ~n16328 & n16334 ) ;
  assign n16336 = ( n16187 & n16328 ) | ( n16187 & n16334 ) | ( n16328 & n16334 ) ;
  assign n16337 = ( n16328 & n16335 ) | ( n16328 & ~n16336 ) | ( n16335 & ~n16336 ) ;
  assign n16338 = ( ~n16190 & n16193 ) | ( ~n16190 & n16337 ) | ( n16193 & n16337 ) ;
  assign n16339 = ( n16190 & n16193 ) | ( n16190 & ~n16337 ) | ( n16193 & ~n16337 ) ;
  assign n16340 = ( ~n16193 & n16338 ) | ( ~n16193 & n16339 ) | ( n16338 & n16339 ) ;
  assign n16341 = n2982 & n9576 ;
  assign n16342 = x35 & n16341 ;
  assign n16343 = x127 & n2989 ;
  assign n16344 = x126 & n2986 ;
  assign n16345 = n16343 | n16344 ;
  assign n16346 = x125 & n3159 ;
  assign n16347 = n16345 | n16346 ;
  assign n16348 = ( ~x35 & n16341 ) | ( ~x35 & n16347 ) | ( n16341 & n16347 ) ;
  assign n16349 = x35 & ~n16347 ;
  assign n16350 = ( ~n16342 & n16348 ) | ( ~n16342 & n16349 ) | ( n16348 & n16349 ) ;
  assign n16351 = n3492 & n8729 ;
  assign n16352 = x38 & n16351 ;
  assign n16353 = x124 & n3499 ;
  assign n16354 = x123 & n3496 ;
  assign n16355 = n16353 | n16354 ;
  assign n16356 = x122 & n3662 ;
  assign n16357 = n16355 | n16356 ;
  assign n16358 = ( ~x38 & n16351 ) | ( ~x38 & n16357 ) | ( n16351 & n16357 ) ;
  assign n16359 = x38 & ~n16357 ;
  assign n16360 = ( ~n16352 & n16358 ) | ( ~n16352 & n16359 ) | ( n16358 & n16359 ) ;
  assign n16361 = n4020 & n7696 ;
  assign n16362 = x41 & n16361 ;
  assign n16363 = x121 & n4027 ;
  assign n16364 = x120 & n4024 ;
  assign n16365 = n16363 | n16364 ;
  assign n16366 = x119 & n4223 ;
  assign n16367 = n16365 | n16366 ;
  assign n16368 = ( ~x41 & n16361 ) | ( ~x41 & n16367 ) | ( n16361 & n16367 ) ;
  assign n16369 = x41 & ~n16367 ;
  assign n16370 = ( ~n16362 & n16368 ) | ( ~n16362 & n16369 ) | ( n16368 & n16369 ) ;
  assign n16371 = n4625 & n6940 ;
  assign n16372 = x44 & n16371 ;
  assign n16373 = x118 & n4791 ;
  assign n16374 = x117 & n4621 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = x116 & n4795 ;
  assign n16377 = n16375 | n16376 ;
  assign n16378 = ( ~x44 & n16371 ) | ( ~x44 & n16377 ) | ( n16371 & n16377 ) ;
  assign n16379 = x44 & ~n16377 ;
  assign n16380 = ( ~n16372 & n16378 ) | ( ~n16372 & n16379 ) | ( n16378 & n16379 ) ;
  assign n16381 = n5223 & n6446 ;
  assign n16382 = x47 & n16381 ;
  assign n16383 = x115 & n5230 ;
  assign n16384 = x114 & n5227 ;
  assign n16385 = n16383 | n16384 ;
  assign n16386 = x113 & n5434 ;
  assign n16387 = n16385 | n16386 ;
  assign n16388 = ( ~x47 & n16381 ) | ( ~x47 & n16387 ) | ( n16381 & n16387 ) ;
  assign n16389 = x47 & ~n16387 ;
  assign n16390 = ( ~n16382 & n16388 ) | ( ~n16382 & n16389 ) | ( n16388 & n16389 ) ;
  assign n16391 = n5558 & n5858 ;
  assign n16392 = x50 & n16391 ;
  assign n16393 = x112 & n5865 ;
  assign n16394 = x111 & n5862 ;
  assign n16395 = n16393 | n16394 ;
  assign n16396 = x110 & n6092 ;
  assign n16397 = n16395 | n16396 ;
  assign n16398 = ( ~x50 & n16391 ) | ( ~x50 & n16397 ) | ( n16391 & n16397 ) ;
  assign n16399 = x50 & ~n16397 ;
  assign n16400 = ( ~n16392 & n16398 ) | ( ~n16392 & n16399 ) | ( n16398 & n16399 ) ;
  assign n16401 = n4930 & n6546 ;
  assign n16402 = x53 & n16401 ;
  assign n16403 = x109 & n6553 ;
  assign n16404 = x108 & n6550 ;
  assign n16405 = n16403 | n16404 ;
  assign n16406 = x107 & n6787 ;
  assign n16407 = n16405 | n16406 ;
  assign n16408 = ( ~x53 & n16401 ) | ( ~x53 & n16407 ) | ( n16401 & n16407 ) ;
  assign n16409 = x53 & ~n16407 ;
  assign n16410 = ( ~n16402 & n16408 ) | ( ~n16402 & n16409 ) | ( n16408 & n16409 ) ;
  assign n16411 = n4331 & n7277 ;
  assign n16412 = x56 & n16411 ;
  assign n16413 = x106 & n7545 ;
  assign n16414 = x105 & n7273 ;
  assign n16415 = n16413 | n16414 ;
  assign n16416 = x104 & n7552 ;
  assign n16417 = n16415 | n16416 ;
  assign n16418 = ( ~x56 & n16411 ) | ( ~x56 & n16417 ) | ( n16411 & n16417 ) ;
  assign n16419 = x56 & ~n16417 ;
  assign n16420 = ( ~n16412 & n16418 ) | ( ~n16412 & n16419 ) | ( n16418 & n16419 ) ;
  assign n16421 = n3941 & n8067 ;
  assign n16422 = x59 & n16421 ;
  assign n16423 = x103 & n8074 ;
  assign n16424 = x102 & n8071 ;
  assign n16425 = n16423 | n16424 ;
  assign n16426 = x101 & n8298 ;
  assign n16427 = n16425 | n16426 ;
  assign n16428 = ( ~x59 & n16421 ) | ( ~x59 & n16427 ) | ( n16421 & n16427 ) ;
  assign n16429 = x59 & ~n16427 ;
  assign n16430 = ( ~n16422 & n16428 ) | ( ~n16422 & n16429 ) | ( n16428 & n16429 ) ;
  assign n16431 = n3264 & n8859 ;
  assign n16432 = x62 & n16431 ;
  assign n16433 = x100 & n8866 ;
  assign n16434 = x99 & n8863 ;
  assign n16435 = n16433 | n16434 ;
  assign n16436 = x98 & n9125 ;
  assign n16437 = n16435 | n16436 ;
  assign n16438 = ( ~x62 & n16431 ) | ( ~x62 & n16437 ) | ( n16431 & n16437 ) ;
  assign n16439 = x62 & ~n16437 ;
  assign n16440 = ( ~n16432 & n16438 ) | ( ~n16432 & n16439 ) | ( n16438 & n16439 ) ;
  assign n16441 = ( x62 & x63 ) | ( x62 & x97 ) | ( x63 & x97 ) ;
  assign n16442 = ( x62 & x96 ) | ( x62 & ~n9394 ) | ( x96 & ~n9394 ) ;
  assign n16443 = ( x96 & n16441 ) | ( x96 & ~n16442 ) | ( n16441 & ~n16442 ) ;
  assign n16444 = ( x32 & n16298 ) | ( x32 & n16443 ) | ( n16298 & n16443 ) ;
  assign n16445 = ( ~x32 & n16298 ) | ( ~x32 & n16443 ) | ( n16298 & n16443 ) ;
  assign n16446 = ( x32 & ~n16444 ) | ( x32 & n16445 ) | ( ~n16444 & n16445 ) ;
  assign n16447 = ( n16300 & n16440 ) | ( n16300 & ~n16446 ) | ( n16440 & ~n16446 ) ;
  assign n16448 = ( ~n16300 & n16440 ) | ( ~n16300 & n16446 ) | ( n16440 & n16446 ) ;
  assign n16449 = ( ~n16440 & n16447 ) | ( ~n16440 & n16448 ) | ( n16447 & n16448 ) ;
  assign n16450 = ( n16303 & n16430 ) | ( n16303 & ~n16449 ) | ( n16430 & ~n16449 ) ;
  assign n16451 = ( n16303 & ~n16430 ) | ( n16303 & n16449 ) | ( ~n16430 & n16449 ) ;
  assign n16452 = ( ~n16303 & n16450 ) | ( ~n16303 & n16451 ) | ( n16450 & n16451 ) ;
  assign n16453 = ( n16305 & n16420 ) | ( n16305 & ~n16452 ) | ( n16420 & ~n16452 ) ;
  assign n16454 = ( n16305 & ~n16420 ) | ( n16305 & n16452 ) | ( ~n16420 & n16452 ) ;
  assign n16455 = ( ~n16305 & n16453 ) | ( ~n16305 & n16454 ) | ( n16453 & n16454 ) ;
  assign n16456 = ( n16308 & n16410 ) | ( n16308 & ~n16455 ) | ( n16410 & ~n16455 ) ;
  assign n16457 = ( ~n16308 & n16410 ) | ( ~n16308 & n16455 ) | ( n16410 & n16455 ) ;
  assign n16458 = ( ~n16410 & n16456 ) | ( ~n16410 & n16457 ) | ( n16456 & n16457 ) ;
  assign n16459 = ( n16311 & n16400 ) | ( n16311 & ~n16458 ) | ( n16400 & ~n16458 ) ;
  assign n16460 = ( n16311 & ~n16400 ) | ( n16311 & n16458 ) | ( ~n16400 & n16458 ) ;
  assign n16461 = ( ~n16311 & n16459 ) | ( ~n16311 & n16460 ) | ( n16459 & n16460 ) ;
  assign n16462 = ( n16315 & n16390 ) | ( n16315 & ~n16461 ) | ( n16390 & ~n16461 ) ;
  assign n16463 = ( n16315 & ~n16390 ) | ( n16315 & n16461 ) | ( ~n16390 & n16461 ) ;
  assign n16464 = ( ~n16315 & n16462 ) | ( ~n16315 & n16463 ) | ( n16462 & n16463 ) ;
  assign n16465 = ( n16317 & n16380 ) | ( n16317 & ~n16464 ) | ( n16380 & ~n16464 ) ;
  assign n16466 = ( n16317 & ~n16380 ) | ( n16317 & n16464 ) | ( ~n16380 & n16464 ) ;
  assign n16467 = ( ~n16317 & n16465 ) | ( ~n16317 & n16466 ) | ( n16465 & n16466 ) ;
  assign n16468 = ( n16320 & n16370 ) | ( n16320 & ~n16467 ) | ( n16370 & ~n16467 ) ;
  assign n16469 = ( n16320 & ~n16370 ) | ( n16320 & n16467 ) | ( ~n16370 & n16467 ) ;
  assign n16470 = ( ~n16320 & n16468 ) | ( ~n16320 & n16469 ) | ( n16468 & n16469 ) ;
  assign n16471 = ( n16323 & n16360 ) | ( n16323 & ~n16470 ) | ( n16360 & ~n16470 ) ;
  assign n16472 = ( n16323 & ~n16360 ) | ( n16323 & n16470 ) | ( ~n16360 & n16470 ) ;
  assign n16473 = ( ~n16323 & n16471 ) | ( ~n16323 & n16472 ) | ( n16471 & n16472 ) ;
  assign n16474 = ( n16326 & n16350 ) | ( n16326 & ~n16473 ) | ( n16350 & ~n16473 ) ;
  assign n16475 = ( n16326 & ~n16350 ) | ( n16326 & n16473 ) | ( ~n16350 & n16473 ) ;
  assign n16476 = ( ~n16326 & n16474 ) | ( ~n16326 & n16475 ) | ( n16474 & n16475 ) ;
  assign n16477 = ( ~n16335 & n16338 ) | ( ~n16335 & n16476 ) | ( n16338 & n16476 ) ;
  assign n16478 = ( n16335 & n16338 ) | ( n16335 & ~n16476 ) | ( n16338 & ~n16476 ) ;
  assign n16479 = ( ~n16338 & n16477 ) | ( ~n16338 & n16478 ) | ( n16477 & n16478 ) ;
  assign n16480 = x126 & n3159 ;
  assign n16481 = x35 & n16480 ;
  assign n16482 = x127 & n2986 ;
  assign n16483 = n2982 | n16482 ;
  assign n16484 = ( n9867 & n16482 ) | ( n9867 & n16483 ) | ( n16482 & n16483 ) ;
  assign n16485 = ( ~x35 & n16480 ) | ( ~x35 & n16484 ) | ( n16480 & n16484 ) ;
  assign n16486 = x35 & ~n16484 ;
  assign n16487 = ( ~n16481 & n16485 ) | ( ~n16481 & n16486 ) | ( n16485 & n16486 ) ;
  assign n16488 = n3492 & n9009 ;
  assign n16489 = x38 & n16488 ;
  assign n16490 = x125 & n3499 ;
  assign n16491 = x124 & n3496 ;
  assign n16492 = n16490 | n16491 ;
  assign n16493 = x123 & n3662 ;
  assign n16494 = n16492 | n16493 ;
  assign n16495 = ( ~x38 & n16488 ) | ( ~x38 & n16494 ) | ( n16488 & n16494 ) ;
  assign n16496 = x38 & ~n16494 ;
  assign n16497 = ( ~n16489 & n16495 ) | ( ~n16489 & n16496 ) | ( n16495 & n16496 ) ;
  assign n16498 = n4020 & n8207 ;
  assign n16499 = x41 & n16498 ;
  assign n16500 = x122 & n4027 ;
  assign n16501 = x121 & n4024 ;
  assign n16502 = n16500 | n16501 ;
  assign n16503 = x120 & n4223 ;
  assign n16504 = n16502 | n16503 ;
  assign n16505 = ( ~x41 & n16498 ) | ( ~x41 & n16504 ) | ( n16498 & n16504 ) ;
  assign n16506 = x41 & ~n16504 ;
  assign n16507 = ( ~n16499 & n16505 ) | ( ~n16499 & n16506 ) | ( n16505 & n16506 ) ;
  assign n16508 = n4625 & n7181 ;
  assign n16509 = x44 & n16508 ;
  assign n16510 = x119 & n4791 ;
  assign n16511 = x118 & n4621 ;
  assign n16512 = n16510 | n16511 ;
  assign n16513 = x117 & n4795 ;
  assign n16514 = n16512 | n16513 ;
  assign n16515 = ( ~x44 & n16508 ) | ( ~x44 & n16514 ) | ( n16508 & n16514 ) ;
  assign n16516 = x44 & ~n16514 ;
  assign n16517 = ( ~n16509 & n16515 ) | ( ~n16509 & n16516 ) | ( n16515 & n16516 ) ;
  assign n16518 = n5223 & n6462 ;
  assign n16519 = x47 & n16518 ;
  assign n16520 = x116 & n5230 ;
  assign n16521 = x115 & n5227 ;
  assign n16522 = n16520 | n16521 ;
  assign n16523 = x114 & n5434 ;
  assign n16524 = n16522 | n16523 ;
  assign n16525 = ( ~x47 & n16518 ) | ( ~x47 & n16524 ) | ( n16518 & n16524 ) ;
  assign n16526 = x47 & ~n16524 ;
  assign n16527 = ( ~n16519 & n16525 ) | ( ~n16519 & n16526 ) | ( n16525 & n16526 ) ;
  assign n16528 = n5774 & n5858 ;
  assign n16529 = x50 & n16528 ;
  assign n16530 = x113 & n5865 ;
  assign n16531 = x112 & n5862 ;
  assign n16532 = n16530 | n16531 ;
  assign n16533 = x111 & n6092 ;
  assign n16534 = n16532 | n16533 ;
  assign n16535 = ( ~x50 & n16528 ) | ( ~x50 & n16534 ) | ( n16528 & n16534 ) ;
  assign n16536 = x50 & ~n16534 ;
  assign n16537 = ( ~n16529 & n16535 ) | ( ~n16529 & n16536 ) | ( n16535 & n16536 ) ;
  assign n16538 = n5331 & n6546 ;
  assign n16539 = x53 & n16538 ;
  assign n16540 = x110 & n6553 ;
  assign n16541 = x109 & n6550 ;
  assign n16542 = n16540 | n16541 ;
  assign n16543 = x108 & n6787 ;
  assign n16544 = n16542 | n16543 ;
  assign n16545 = ( ~x53 & n16538 ) | ( ~x53 & n16544 ) | ( n16538 & n16544 ) ;
  assign n16546 = x53 & ~n16544 ;
  assign n16547 = ( ~n16539 & n16545 ) | ( ~n16539 & n16546 ) | ( n16545 & n16546 ) ;
  assign n16548 = n4523 & n7277 ;
  assign n16549 = x56 & n16548 ;
  assign n16550 = x107 & n7545 ;
  assign n16551 = x106 & n7273 ;
  assign n16552 = n16550 | n16551 ;
  assign n16553 = x105 & n7552 ;
  assign n16554 = n16552 | n16553 ;
  assign n16555 = ( ~x56 & n16548 ) | ( ~x56 & n16554 ) | ( n16548 & n16554 ) ;
  assign n16556 = x56 & ~n16554 ;
  assign n16557 = ( ~n16549 & n16555 ) | ( ~n16549 & n16556 ) | ( n16555 & n16556 ) ;
  assign n16558 = n3957 & n8067 ;
  assign n16559 = x59 & n16558 ;
  assign n16560 = x104 & n8074 ;
  assign n16561 = x103 & n8071 ;
  assign n16562 = n16560 | n16561 ;
  assign n16563 = x102 & n8298 ;
  assign n16564 = n16562 | n16563 ;
  assign n16565 = ( ~x59 & n16558 ) | ( ~x59 & n16564 ) | ( n16558 & n16564 ) ;
  assign n16566 = x59 & ~n16564 ;
  assign n16567 = ( ~n16559 & n16565 ) | ( ~n16559 & n16566 ) | ( n16565 & n16566 ) ;
  assign n16568 = ( x62 & x63 ) | ( x62 & x98 ) | ( x63 & x98 ) ;
  assign n16569 = ( x62 & x97 ) | ( x62 & ~n9394 ) | ( x97 & ~n9394 ) ;
  assign n16570 = ( x97 & n16568 ) | ( x97 & ~n16569 ) | ( n16568 & ~n16569 ) ;
  assign n16571 = n3591 & n8859 ;
  assign n16572 = x62 & n16571 ;
  assign n16573 = x101 & n8866 ;
  assign n16574 = x100 & n8863 ;
  assign n16575 = n16573 | n16574 ;
  assign n16576 = x99 & n9125 ;
  assign n16577 = n16575 | n16576 ;
  assign n16578 = ( ~x62 & n16571 ) | ( ~x62 & n16577 ) | ( n16571 & n16577 ) ;
  assign n16579 = x62 & ~n16577 ;
  assign n16580 = ( ~n16572 & n16578 ) | ( ~n16572 & n16579 ) | ( n16578 & n16579 ) ;
  assign n16581 = ( ~n16445 & n16570 ) | ( ~n16445 & n16580 ) | ( n16570 & n16580 ) ;
  assign n16582 = ( n16445 & n16570 ) | ( n16445 & ~n16580 ) | ( n16570 & ~n16580 ) ;
  assign n16583 = ( ~n16570 & n16581 ) | ( ~n16570 & n16582 ) | ( n16581 & n16582 ) ;
  assign n16584 = ( ~n16447 & n16567 ) | ( ~n16447 & n16583 ) | ( n16567 & n16583 ) ;
  assign n16585 = ( n16447 & n16567 ) | ( n16447 & ~n16583 ) | ( n16567 & ~n16583 ) ;
  assign n16586 = ( ~n16567 & n16584 ) | ( ~n16567 & n16585 ) | ( n16584 & n16585 ) ;
  assign n16587 = ( n16450 & n16557 ) | ( n16450 & ~n16586 ) | ( n16557 & ~n16586 ) ;
  assign n16588 = ( ~n16450 & n16557 ) | ( ~n16450 & n16586 ) | ( n16557 & n16586 ) ;
  assign n16589 = ( ~n16557 & n16587 ) | ( ~n16557 & n16588 ) | ( n16587 & n16588 ) ;
  assign n16590 = ( n16453 & n16547 ) | ( n16453 & ~n16589 ) | ( n16547 & ~n16589 ) ;
  assign n16591 = ( ~n16453 & n16547 ) | ( ~n16453 & n16589 ) | ( n16547 & n16589 ) ;
  assign n16592 = ( ~n16547 & n16590 ) | ( ~n16547 & n16591 ) | ( n16590 & n16591 ) ;
  assign n16593 = ( n16456 & n16537 ) | ( n16456 & ~n16592 ) | ( n16537 & ~n16592 ) ;
  assign n16594 = ( ~n16456 & n16537 ) | ( ~n16456 & n16592 ) | ( n16537 & n16592 ) ;
  assign n16595 = ( ~n16537 & n16593 ) | ( ~n16537 & n16594 ) | ( n16593 & n16594 ) ;
  assign n16596 = ( n16459 & n16527 ) | ( n16459 & ~n16595 ) | ( n16527 & ~n16595 ) ;
  assign n16597 = ( ~n16459 & n16527 ) | ( ~n16459 & n16595 ) | ( n16527 & n16595 ) ;
  assign n16598 = ( ~n16527 & n16596 ) | ( ~n16527 & n16597 ) | ( n16596 & n16597 ) ;
  assign n16599 = ( n16462 & n16517 ) | ( n16462 & ~n16598 ) | ( n16517 & ~n16598 ) ;
  assign n16600 = ( ~n16462 & n16517 ) | ( ~n16462 & n16598 ) | ( n16517 & n16598 ) ;
  assign n16601 = ( ~n16517 & n16599 ) | ( ~n16517 & n16600 ) | ( n16599 & n16600 ) ;
  assign n16602 = ( n16465 & n16507 ) | ( n16465 & ~n16601 ) | ( n16507 & ~n16601 ) ;
  assign n16603 = ( ~n16465 & n16507 ) | ( ~n16465 & n16601 ) | ( n16507 & n16601 ) ;
  assign n16604 = ( ~n16507 & n16602 ) | ( ~n16507 & n16603 ) | ( n16602 & n16603 ) ;
  assign n16605 = ( n16468 & n16497 ) | ( n16468 & ~n16604 ) | ( n16497 & ~n16604 ) ;
  assign n16606 = ( ~n16468 & n16497 ) | ( ~n16468 & n16604 ) | ( n16497 & n16604 ) ;
  assign n16607 = ( ~n16497 & n16605 ) | ( ~n16497 & n16606 ) | ( n16605 & n16606 ) ;
  assign n16608 = ( n16471 & n16487 ) | ( n16471 & ~n16607 ) | ( n16487 & ~n16607 ) ;
  assign n16609 = ( ~n16471 & n16487 ) | ( ~n16471 & n16607 ) | ( n16487 & n16607 ) ;
  assign n16610 = ( ~n16487 & n16608 ) | ( ~n16487 & n16609 ) | ( n16608 & n16609 ) ;
  assign n16611 = ( ~n16474 & n16477 ) | ( ~n16474 & n16610 ) | ( n16477 & n16610 ) ;
  assign n16612 = ( n16474 & n16477 ) | ( n16474 & ~n16610 ) | ( n16477 & ~n16610 ) ;
  assign n16613 = ( ~n16477 & n16611 ) | ( ~n16477 & n16612 ) | ( n16611 & n16612 ) ;
  assign n16614 = n3492 & n9038 ;
  assign n16615 = x38 & n16614 ;
  assign n16616 = x126 & n3499 ;
  assign n16617 = x125 & n3496 ;
  assign n16618 = n16616 | n16617 ;
  assign n16619 = x124 & n3662 ;
  assign n16620 = n16618 | n16619 ;
  assign n16621 = ( ~x38 & n16614 ) | ( ~x38 & n16620 ) | ( n16614 & n16620 ) ;
  assign n16622 = x38 & ~n16620 ;
  assign n16623 = ( ~n16615 & n16621 ) | ( ~n16615 & n16622 ) | ( n16621 & n16622 ) ;
  assign n16624 = n4020 & n8461 ;
  assign n16625 = x41 & n16624 ;
  assign n16626 = x123 & n4027 ;
  assign n16627 = x122 & n4024 ;
  assign n16628 = n16626 | n16627 ;
  assign n16629 = x121 & n4223 ;
  assign n16630 = n16628 | n16629 ;
  assign n16631 = ( ~x41 & n16624 ) | ( ~x41 & n16630 ) | ( n16624 & n16630 ) ;
  assign n16632 = x41 & ~n16630 ;
  assign n16633 = ( ~n16625 & n16631 ) | ( ~n16625 & n16632 ) | ( n16631 & n16632 ) ;
  assign n16634 = n4625 & n7444 ;
  assign n16635 = x44 & n16634 ;
  assign n16636 = x120 & n4791 ;
  assign n16637 = x119 & n4621 ;
  assign n16638 = n16636 | n16637 ;
  assign n16639 = x118 & n4795 ;
  assign n16640 = n16638 | n16639 ;
  assign n16641 = ( ~x44 & n16634 ) | ( ~x44 & n16640 ) | ( n16634 & n16640 ) ;
  assign n16642 = x44 & ~n16640 ;
  assign n16643 = ( ~n16635 & n16641 ) | ( ~n16635 & n16642 ) | ( n16641 & n16642 ) ;
  assign n16644 = n5223 & n6924 ;
  assign n16645 = x47 & n16644 ;
  assign n16646 = x117 & n5230 ;
  assign n16647 = x116 & n5227 ;
  assign n16648 = n16646 | n16647 ;
  assign n16649 = x115 & n5434 ;
  assign n16650 = n16648 | n16649 ;
  assign n16651 = ( ~x47 & n16644 ) | ( ~x47 & n16650 ) | ( n16644 & n16650 ) ;
  assign n16652 = x47 & ~n16650 ;
  assign n16653 = ( ~n16645 & n16651 ) | ( ~n16645 & n16652 ) | ( n16651 & n16652 ) ;
  assign n16654 = n5858 & n6002 ;
  assign n16655 = x50 & n16654 ;
  assign n16656 = x114 & n5865 ;
  assign n16657 = x113 & n5862 ;
  assign n16658 = n16656 | n16657 ;
  assign n16659 = x112 & n6092 ;
  assign n16660 = n16658 | n16659 ;
  assign n16661 = ( ~x50 & n16654 ) | ( ~x50 & n16660 ) | ( n16654 & n16660 ) ;
  assign n16662 = x50 & ~n16660 ;
  assign n16663 = ( ~n16655 & n16661 ) | ( ~n16655 & n16662 ) | ( n16661 & n16662 ) ;
  assign n16664 = n5347 & n6546 ;
  assign n16665 = x53 & n16664 ;
  assign n16666 = x111 & n6553 ;
  assign n16667 = x110 & n6550 ;
  assign n16668 = n16666 | n16667 ;
  assign n16669 = x109 & n6787 ;
  assign n16670 = n16668 | n16669 ;
  assign n16671 = ( ~x53 & n16664 ) | ( ~x53 & n16670 ) | ( n16664 & n16670 ) ;
  assign n16672 = x53 & ~n16670 ;
  assign n16673 = ( ~n16665 & n16671 ) | ( ~n16665 & n16672 ) | ( n16671 & n16672 ) ;
  assign n16674 = n4914 & n7277 ;
  assign n16675 = x56 & n16674 ;
  assign n16676 = x108 & n7545 ;
  assign n16677 = x107 & n7273 ;
  assign n16678 = n16676 | n16677 ;
  assign n16679 = x106 & n7552 ;
  assign n16680 = n16678 | n16679 ;
  assign n16681 = ( ~x56 & n16674 ) | ( ~x56 & n16680 ) | ( n16674 & n16680 ) ;
  assign n16682 = x56 & ~n16680 ;
  assign n16683 = ( ~n16675 & n16681 ) | ( ~n16675 & n16682 ) | ( n16681 & n16682 ) ;
  assign n16684 = n4145 & n8067 ;
  assign n16685 = x59 & n16684 ;
  assign n16686 = x105 & n8074 ;
  assign n16687 = x104 & n8071 ;
  assign n16688 = n16686 | n16687 ;
  assign n16689 = x103 & n8298 ;
  assign n16690 = n16688 | n16689 ;
  assign n16691 = ( ~x59 & n16684 ) | ( ~x59 & n16690 ) | ( n16684 & n16690 ) ;
  assign n16692 = x59 & ~n16690 ;
  assign n16693 = ( ~n16685 & n16691 ) | ( ~n16685 & n16692 ) | ( n16691 & n16692 ) ;
  assign n16694 = n3764 & n8859 ;
  assign n16695 = x62 & n16694 ;
  assign n16696 = x102 & n8866 ;
  assign n16697 = x101 & n8863 ;
  assign n16698 = n16696 | n16697 ;
  assign n16699 = x100 & n9125 ;
  assign n16700 = n16698 | n16699 ;
  assign n16701 = ( ~x62 & n16694 ) | ( ~x62 & n16700 ) | ( n16694 & n16700 ) ;
  assign n16702 = x62 & ~n16700 ;
  assign n16703 = ( ~n16695 & n16701 ) | ( ~n16695 & n16702 ) | ( n16701 & n16702 ) ;
  assign n16704 = ( x62 & x63 ) | ( x62 & x99 ) | ( x63 & x99 ) ;
  assign n16705 = ( x62 & x98 ) | ( x62 & ~n9394 ) | ( x98 & ~n9394 ) ;
  assign n16706 = ( x98 & n16704 ) | ( x98 & ~n16705 ) | ( n16704 & ~n16705 ) ;
  assign n16707 = ( n16580 & ~n16582 ) | ( n16580 & n16706 ) | ( ~n16582 & n16706 ) ;
  assign n16708 = ( n16445 & n16581 ) | ( n16445 & ~n16706 ) | ( n16581 & ~n16706 ) ;
  assign n16709 = ( ~n16580 & n16707 ) | ( ~n16580 & n16708 ) | ( n16707 & n16708 ) ;
  assign n16710 = ( n16693 & ~n16703 ) | ( n16693 & n16709 ) | ( ~n16703 & n16709 ) ;
  assign n16711 = ( n16693 & n16703 ) | ( n16693 & ~n16709 ) | ( n16703 & ~n16709 ) ;
  assign n16712 = ( ~n16693 & n16710 ) | ( ~n16693 & n16711 ) | ( n16710 & n16711 ) ;
  assign n16713 = ( n16585 & n16683 ) | ( n16585 & ~n16712 ) | ( n16683 & ~n16712 ) ;
  assign n16714 = ( n16585 & ~n16683 ) | ( n16585 & n16712 ) | ( ~n16683 & n16712 ) ;
  assign n16715 = ( ~n16585 & n16713 ) | ( ~n16585 & n16714 ) | ( n16713 & n16714 ) ;
  assign n16716 = ( n16587 & n16673 ) | ( n16587 & ~n16715 ) | ( n16673 & ~n16715 ) ;
  assign n16717 = ( ~n16587 & n16673 ) | ( ~n16587 & n16715 ) | ( n16673 & n16715 ) ;
  assign n16718 = ( ~n16673 & n16716 ) | ( ~n16673 & n16717 ) | ( n16716 & n16717 ) ;
  assign n16719 = ( n16590 & n16663 ) | ( n16590 & ~n16718 ) | ( n16663 & ~n16718 ) ;
  assign n16720 = ( ~n16590 & n16663 ) | ( ~n16590 & n16718 ) | ( n16663 & n16718 ) ;
  assign n16721 = ( ~n16663 & n16719 ) | ( ~n16663 & n16720 ) | ( n16719 & n16720 ) ;
  assign n16722 = ( n16593 & n16653 ) | ( n16593 & ~n16721 ) | ( n16653 & ~n16721 ) ;
  assign n16723 = ( ~n16593 & n16653 ) | ( ~n16593 & n16721 ) | ( n16653 & n16721 ) ;
  assign n16724 = ( ~n16653 & n16722 ) | ( ~n16653 & n16723 ) | ( n16722 & n16723 ) ;
  assign n16725 = ( n16596 & n16643 ) | ( n16596 & ~n16724 ) | ( n16643 & ~n16724 ) ;
  assign n16726 = ( ~n16596 & n16643 ) | ( ~n16596 & n16724 ) | ( n16643 & n16724 ) ;
  assign n16727 = ( ~n16643 & n16725 ) | ( ~n16643 & n16726 ) | ( n16725 & n16726 ) ;
  assign n16728 = ( n16599 & n16633 ) | ( n16599 & ~n16727 ) | ( n16633 & ~n16727 ) ;
  assign n16729 = ( ~n16599 & n16633 ) | ( ~n16599 & n16727 ) | ( n16633 & n16727 ) ;
  assign n16730 = ( ~n16633 & n16728 ) | ( ~n16633 & n16729 ) | ( n16728 & n16729 ) ;
  assign n16731 = ( n16602 & n16623 ) | ( n16602 & ~n16730 ) | ( n16623 & ~n16730 ) ;
  assign n16732 = ( ~n16602 & n16623 ) | ( ~n16602 & n16730 ) | ( n16623 & n16730 ) ;
  assign n16733 = ( ~n16623 & n16731 ) | ( ~n16623 & n16732 ) | ( n16731 & n16732 ) ;
  assign n16734 = x127 & n3159 ;
  assign n16735 = n2982 | n16734 ;
  assign n16736 = ( n9865 & n16734 ) | ( n9865 & n16735 ) | ( n16734 & n16735 ) ;
  assign n16737 = x35 & ~n16736 ;
  assign n16738 = ~x35 & n16736 ;
  assign n16739 = n16737 | n16738 ;
  assign n16740 = ( n16605 & ~n16733 ) | ( n16605 & n16739 ) | ( ~n16733 & n16739 ) ;
  assign n16741 = ( n16605 & n16733 ) | ( n16605 & n16739 ) | ( n16733 & n16739 ) ;
  assign n16742 = ( n16733 & n16740 ) | ( n16733 & ~n16741 ) | ( n16740 & ~n16741 ) ;
  assign n16743 = ( ~n16608 & n16611 ) | ( ~n16608 & n16742 ) | ( n16611 & n16742 ) ;
  assign n16744 = ( n16608 & n16611 ) | ( n16608 & ~n16742 ) | ( n16611 & ~n16742 ) ;
  assign n16745 = ( ~n16611 & n16743 ) | ( ~n16611 & n16744 ) | ( n16743 & n16744 ) ;
  assign n16746 = n4020 & n8729 ;
  assign n16747 = x41 & n16746 ;
  assign n16748 = x124 & n4027 ;
  assign n16749 = x123 & n4024 ;
  assign n16750 = n16748 | n16749 ;
  assign n16751 = x122 & n4223 ;
  assign n16752 = n16750 | n16751 ;
  assign n16753 = ( ~x41 & n16746 ) | ( ~x41 & n16752 ) | ( n16746 & n16752 ) ;
  assign n16754 = x41 & ~n16752 ;
  assign n16755 = ( ~n16747 & n16753 ) | ( ~n16747 & n16754 ) | ( n16753 & n16754 ) ;
  assign n16756 = n4625 & n7696 ;
  assign n16757 = x44 & n16756 ;
  assign n16758 = x121 & n4791 ;
  assign n16759 = x120 & n4621 ;
  assign n16760 = n16758 | n16759 ;
  assign n16761 = x119 & n4795 ;
  assign n16762 = n16760 | n16761 ;
  assign n16763 = ( ~x44 & n16756 ) | ( ~x44 & n16762 ) | ( n16756 & n16762 ) ;
  assign n16764 = x44 & ~n16762 ;
  assign n16765 = ( ~n16757 & n16763 ) | ( ~n16757 & n16764 ) | ( n16763 & n16764 ) ;
  assign n16766 = n5223 & n6940 ;
  assign n16767 = x47 & n16766 ;
  assign n16768 = x118 & n5230 ;
  assign n16769 = x117 & n5227 ;
  assign n16770 = n16768 | n16769 ;
  assign n16771 = x116 & n5434 ;
  assign n16772 = n16770 | n16771 ;
  assign n16773 = ( ~x47 & n16766 ) | ( ~x47 & n16772 ) | ( n16766 & n16772 ) ;
  assign n16774 = x47 & ~n16772 ;
  assign n16775 = ( ~n16767 & n16773 ) | ( ~n16767 & n16774 ) | ( n16773 & n16774 ) ;
  assign n16776 = n5858 & n6446 ;
  assign n16777 = x50 & n16776 ;
  assign n16778 = x115 & n5865 ;
  assign n16779 = x114 & n5862 ;
  assign n16780 = n16778 | n16779 ;
  assign n16781 = x113 & n6092 ;
  assign n16782 = n16780 | n16781 ;
  assign n16783 = ( ~x50 & n16776 ) | ( ~x50 & n16782 ) | ( n16776 & n16782 ) ;
  assign n16784 = x50 & ~n16782 ;
  assign n16785 = ( ~n16777 & n16783 ) | ( ~n16777 & n16784 ) | ( n16783 & n16784 ) ;
  assign n16786 = n5558 & n6546 ;
  assign n16787 = x53 & n16786 ;
  assign n16788 = x112 & n6553 ;
  assign n16789 = x111 & n6550 ;
  assign n16790 = n16788 | n16789 ;
  assign n16791 = x110 & n6787 ;
  assign n16792 = n16790 | n16791 ;
  assign n16793 = ( ~x53 & n16786 ) | ( ~x53 & n16792 ) | ( n16786 & n16792 ) ;
  assign n16794 = x53 & ~n16792 ;
  assign n16795 = ( ~n16787 & n16793 ) | ( ~n16787 & n16794 ) | ( n16793 & n16794 ) ;
  assign n16796 = n4930 & n7277 ;
  assign n16797 = x56 & n16796 ;
  assign n16798 = x109 & n7545 ;
  assign n16799 = x108 & n7273 ;
  assign n16800 = n16798 | n16799 ;
  assign n16801 = x107 & n7552 ;
  assign n16802 = n16800 | n16801 ;
  assign n16803 = ( ~x56 & n16796 ) | ( ~x56 & n16802 ) | ( n16796 & n16802 ) ;
  assign n16804 = x56 & ~n16802 ;
  assign n16805 = ( ~n16797 & n16803 ) | ( ~n16797 & n16804 ) | ( n16803 & n16804 ) ;
  assign n16806 = n4331 & n8067 ;
  assign n16807 = x59 & n16806 ;
  assign n16808 = x106 & n8074 ;
  assign n16809 = x105 & n8071 ;
  assign n16810 = n16808 | n16809 ;
  assign n16811 = x104 & n8298 ;
  assign n16812 = n16810 | n16811 ;
  assign n16813 = ( ~x59 & n16806 ) | ( ~x59 & n16812 ) | ( n16806 & n16812 ) ;
  assign n16814 = x59 & ~n16812 ;
  assign n16815 = ( ~n16807 & n16813 ) | ( ~n16807 & n16814 ) | ( n16813 & n16814 ) ;
  assign n16816 = n3941 & n8859 ;
  assign n16817 = x62 & n16816 ;
  assign n16818 = x103 & n8866 ;
  assign n16819 = x102 & n8863 ;
  assign n16820 = n16818 | n16819 ;
  assign n16821 = x101 & n9125 ;
  assign n16822 = n16820 | n16821 ;
  assign n16823 = ( ~x62 & n16816 ) | ( ~x62 & n16822 ) | ( n16816 & n16822 ) ;
  assign n16824 = x62 & ~n16822 ;
  assign n16825 = ( ~n16817 & n16823 ) | ( ~n16817 & n16824 ) | ( n16823 & n16824 ) ;
  assign n16826 = ( x62 & x63 ) | ( x62 & x100 ) | ( x63 & x100 ) ;
  assign n16827 = ( x62 & x99 ) | ( x62 & ~n9394 ) | ( x99 & ~n9394 ) ;
  assign n16828 = ( x99 & n16826 ) | ( x99 & ~n16827 ) | ( n16826 & ~n16827 ) ;
  assign n16829 = ( x35 & n16706 ) | ( x35 & n16828 ) | ( n16706 & n16828 ) ;
  assign n16830 = ( ~x35 & n16706 ) | ( ~x35 & n16828 ) | ( n16706 & n16828 ) ;
  assign n16831 = ( x35 & ~n16829 ) | ( x35 & n16830 ) | ( ~n16829 & n16830 ) ;
  assign n16832 = ( n16708 & n16825 ) | ( n16708 & ~n16831 ) | ( n16825 & ~n16831 ) ;
  assign n16833 = ( ~n16708 & n16825 ) | ( ~n16708 & n16831 ) | ( n16825 & n16831 ) ;
  assign n16834 = ( ~n16825 & n16832 ) | ( ~n16825 & n16833 ) | ( n16832 & n16833 ) ;
  assign n16835 = ( n16711 & n16815 ) | ( n16711 & ~n16834 ) | ( n16815 & ~n16834 ) ;
  assign n16836 = ( n16711 & ~n16815 ) | ( n16711 & n16834 ) | ( ~n16815 & n16834 ) ;
  assign n16837 = ( ~n16711 & n16835 ) | ( ~n16711 & n16836 ) | ( n16835 & n16836 ) ;
  assign n16838 = ( n16713 & ~n16805 ) | ( n16713 & n16837 ) | ( ~n16805 & n16837 ) ;
  assign n16839 = ( n16713 & n16805 ) | ( n16713 & ~n16837 ) | ( n16805 & ~n16837 ) ;
  assign n16840 = ( ~n16713 & n16838 ) | ( ~n16713 & n16839 ) | ( n16838 & n16839 ) ;
  assign n16841 = ( n16716 & n16795 ) | ( n16716 & ~n16840 ) | ( n16795 & ~n16840 ) ;
  assign n16842 = ( n16716 & ~n16795 ) | ( n16716 & n16840 ) | ( ~n16795 & n16840 ) ;
  assign n16843 = ( ~n16716 & n16841 ) | ( ~n16716 & n16842 ) | ( n16841 & n16842 ) ;
  assign n16844 = ( n16719 & n16785 ) | ( n16719 & ~n16843 ) | ( n16785 & ~n16843 ) ;
  assign n16845 = ( n16719 & ~n16785 ) | ( n16719 & n16843 ) | ( ~n16785 & n16843 ) ;
  assign n16846 = ( ~n16719 & n16844 ) | ( ~n16719 & n16845 ) | ( n16844 & n16845 ) ;
  assign n16847 = ( n16722 & n16775 ) | ( n16722 & ~n16846 ) | ( n16775 & ~n16846 ) ;
  assign n16848 = ( n16722 & ~n16775 ) | ( n16722 & n16846 ) | ( ~n16775 & n16846 ) ;
  assign n16849 = ( ~n16722 & n16847 ) | ( ~n16722 & n16848 ) | ( n16847 & n16848 ) ;
  assign n16850 = ( n16725 & ~n16765 ) | ( n16725 & n16849 ) | ( ~n16765 & n16849 ) ;
  assign n16851 = ( n16725 & n16765 ) | ( n16725 & ~n16849 ) | ( n16765 & ~n16849 ) ;
  assign n16852 = ( ~n16725 & n16850 ) | ( ~n16725 & n16851 ) | ( n16850 & n16851 ) ;
  assign n16853 = ( n16728 & ~n16755 ) | ( n16728 & n16852 ) | ( ~n16755 & n16852 ) ;
  assign n16854 = ( n16728 & n16755 ) | ( n16728 & ~n16852 ) | ( n16755 & ~n16852 ) ;
  assign n16855 = ( ~n16728 & n16853 ) | ( ~n16728 & n16854 ) | ( n16853 & n16854 ) ;
  assign n16856 = n3492 & n9576 ;
  assign n16857 = x38 & n16856 ;
  assign n16858 = x127 & n3499 ;
  assign n16859 = x126 & n3496 ;
  assign n16860 = n16858 | n16859 ;
  assign n16861 = x125 & n3662 ;
  assign n16862 = n16860 | n16861 ;
  assign n16863 = ( ~x38 & n16856 ) | ( ~x38 & n16862 ) | ( n16856 & n16862 ) ;
  assign n16864 = x38 & ~n16862 ;
  assign n16865 = ( ~n16857 & n16863 ) | ( ~n16857 & n16864 ) | ( n16863 & n16864 ) ;
  assign n16866 = ( n16731 & ~n16855 ) | ( n16731 & n16865 ) | ( ~n16855 & n16865 ) ;
  assign n16867 = ( n16731 & n16855 ) | ( n16731 & ~n16865 ) | ( n16855 & ~n16865 ) ;
  assign n16868 = ( ~n16731 & n16866 ) | ( ~n16731 & n16867 ) | ( n16866 & n16867 ) ;
  assign n16869 = ( ~n16740 & n16743 ) | ( ~n16740 & n16868 ) | ( n16743 & n16868 ) ;
  assign n16870 = ( n16740 & n16743 ) | ( n16740 & ~n16868 ) | ( n16743 & ~n16868 ) ;
  assign n16871 = ( ~n16743 & n16869 ) | ( ~n16743 & n16870 ) | ( n16869 & n16870 ) ;
  assign n16872 = x127 & n3496 ;
  assign n16873 = n3492 | n16872 ;
  assign n16874 = ( n9867 & n16872 ) | ( n9867 & n16873 ) | ( n16872 & n16873 ) ;
  assign n16875 = x126 & n3662 ;
  assign n16876 = ( ~x38 & n16874 ) | ( ~x38 & n16875 ) | ( n16874 & n16875 ) ;
  assign n16877 = ( x38 & ~n16874 ) | ( x38 & n16875 ) | ( ~n16874 & n16875 ) ;
  assign n16878 = ~n16875 & n16877 ;
  assign n16879 = n16876 | n16878 ;
  assign n16880 = n4020 & n9009 ;
  assign n16881 = x41 & n16880 ;
  assign n16882 = x125 & n4027 ;
  assign n16883 = x124 & n4024 ;
  assign n16884 = n16882 | n16883 ;
  assign n16885 = x123 & n4223 ;
  assign n16886 = n16884 | n16885 ;
  assign n16887 = ( ~x41 & n16880 ) | ( ~x41 & n16886 ) | ( n16880 & n16886 ) ;
  assign n16888 = x41 & ~n16886 ;
  assign n16889 = ( ~n16881 & n16887 ) | ( ~n16881 & n16888 ) | ( n16887 & n16888 ) ;
  assign n16890 = n4625 & n8207 ;
  assign n16891 = x44 & n16890 ;
  assign n16892 = x122 & n4791 ;
  assign n16893 = x121 & n4621 ;
  assign n16894 = n16892 | n16893 ;
  assign n16895 = x120 & n4795 ;
  assign n16896 = n16894 | n16895 ;
  assign n16897 = ( ~x44 & n16890 ) | ( ~x44 & n16896 ) | ( n16890 & n16896 ) ;
  assign n16898 = x44 & ~n16896 ;
  assign n16899 = ( ~n16891 & n16897 ) | ( ~n16891 & n16898 ) | ( n16897 & n16898 ) ;
  assign n16900 = n5223 & n7181 ;
  assign n16901 = x47 & n16900 ;
  assign n16902 = x119 & n5230 ;
  assign n16903 = x118 & n5227 ;
  assign n16904 = n16902 | n16903 ;
  assign n16905 = x117 & n5434 ;
  assign n16906 = n16904 | n16905 ;
  assign n16907 = ( ~x47 & n16900 ) | ( ~x47 & n16906 ) | ( n16900 & n16906 ) ;
  assign n16908 = x47 & ~n16906 ;
  assign n16909 = ( ~n16901 & n16907 ) | ( ~n16901 & n16908 ) | ( n16907 & n16908 ) ;
  assign n16910 = n5858 & n6462 ;
  assign n16911 = x50 & n16910 ;
  assign n16912 = x116 & n5865 ;
  assign n16913 = x115 & n5862 ;
  assign n16914 = n16912 | n16913 ;
  assign n16915 = x114 & n6092 ;
  assign n16916 = n16914 | n16915 ;
  assign n16917 = ( ~x50 & n16910 ) | ( ~x50 & n16916 ) | ( n16910 & n16916 ) ;
  assign n16918 = x50 & ~n16916 ;
  assign n16919 = ( ~n16911 & n16917 ) | ( ~n16911 & n16918 ) | ( n16917 & n16918 ) ;
  assign n16920 = n5774 & n6546 ;
  assign n16921 = x53 & n16920 ;
  assign n16922 = x113 & n6553 ;
  assign n16923 = x112 & n6550 ;
  assign n16924 = n16922 | n16923 ;
  assign n16925 = x111 & n6787 ;
  assign n16926 = n16924 | n16925 ;
  assign n16927 = ( ~x53 & n16920 ) | ( ~x53 & n16926 ) | ( n16920 & n16926 ) ;
  assign n16928 = x53 & ~n16926 ;
  assign n16929 = ( ~n16921 & n16927 ) | ( ~n16921 & n16928 ) | ( n16927 & n16928 ) ;
  assign n16930 = n5331 & n7277 ;
  assign n16931 = x56 & n16930 ;
  assign n16932 = x110 & n7545 ;
  assign n16933 = x109 & n7273 ;
  assign n16934 = n16932 | n16933 ;
  assign n16935 = x108 & n7552 ;
  assign n16936 = n16934 | n16935 ;
  assign n16937 = ( ~x56 & n16930 ) | ( ~x56 & n16936 ) | ( n16930 & n16936 ) ;
  assign n16938 = x56 & ~n16936 ;
  assign n16939 = ( ~n16931 & n16937 ) | ( ~n16931 & n16938 ) | ( n16937 & n16938 ) ;
  assign n16940 = n4523 & n8067 ;
  assign n16941 = x59 & n16940 ;
  assign n16942 = x107 & n8074 ;
  assign n16943 = x106 & n8071 ;
  assign n16944 = n16942 | n16943 ;
  assign n16945 = x105 & n8298 ;
  assign n16946 = n16944 | n16945 ;
  assign n16947 = ( ~x59 & n16940 ) | ( ~x59 & n16946 ) | ( n16940 & n16946 ) ;
  assign n16948 = x59 & ~n16946 ;
  assign n16949 = ( ~n16941 & n16947 ) | ( ~n16941 & n16948 ) | ( n16947 & n16948 ) ;
  assign n16950 = ( x62 & x63 ) | ( x62 & x101 ) | ( x63 & x101 ) ;
  assign n16951 = ( x62 & x100 ) | ( x62 & ~n9394 ) | ( x100 & ~n9394 ) ;
  assign n16952 = ( x100 & n16950 ) | ( x100 & ~n16951 ) | ( n16950 & ~n16951 ) ;
  assign n16953 = x103 & n8863 ;
  assign n16954 = x102 | n16953 ;
  assign n16955 = ( n9125 & n16953 ) | ( n9125 & n16954 ) | ( n16953 & n16954 ) ;
  assign n16956 = n3957 & n8859 ;
  assign n16957 = n16955 | n16956 ;
  assign n16958 = x104 & n8866 ;
  assign n16959 = ( ~x62 & n16957 ) | ( ~x62 & n16958 ) | ( n16957 & n16958 ) ;
  assign n16960 = ( x62 & ~n16957 ) | ( x62 & n16958 ) | ( ~n16957 & n16958 ) ;
  assign n16961 = ~n16958 & n16960 ;
  assign n16962 = n16959 | n16961 ;
  assign n16963 = ( ~n16830 & n16952 ) | ( ~n16830 & n16962 ) | ( n16952 & n16962 ) ;
  assign n16964 = ( n16830 & n16952 ) | ( n16830 & ~n16962 ) | ( n16952 & ~n16962 ) ;
  assign n16965 = ( ~n16952 & n16963 ) | ( ~n16952 & n16964 ) | ( n16963 & n16964 ) ;
  assign n16966 = ( n16832 & n16949 ) | ( n16832 & ~n16965 ) | ( n16949 & ~n16965 ) ;
  assign n16967 = ( ~n16832 & n16949 ) | ( ~n16832 & n16965 ) | ( n16949 & n16965 ) ;
  assign n16968 = ( ~n16949 & n16966 ) | ( ~n16949 & n16967 ) | ( n16966 & n16967 ) ;
  assign n16969 = ( n16835 & n16939 ) | ( n16835 & ~n16968 ) | ( n16939 & ~n16968 ) ;
  assign n16970 = ( ~n16835 & n16939 ) | ( ~n16835 & n16968 ) | ( n16939 & n16968 ) ;
  assign n16971 = ( ~n16939 & n16969 ) | ( ~n16939 & n16970 ) | ( n16969 & n16970 ) ;
  assign n16972 = ( n16839 & n16929 ) | ( n16839 & ~n16971 ) | ( n16929 & ~n16971 ) ;
  assign n16973 = ( ~n16839 & n16929 ) | ( ~n16839 & n16971 ) | ( n16929 & n16971 ) ;
  assign n16974 = ( ~n16929 & n16972 ) | ( ~n16929 & n16973 ) | ( n16972 & n16973 ) ;
  assign n16975 = ( n16841 & n16919 ) | ( n16841 & ~n16974 ) | ( n16919 & ~n16974 ) ;
  assign n16976 = ( ~n16841 & n16919 ) | ( ~n16841 & n16974 ) | ( n16919 & n16974 ) ;
  assign n16977 = ( ~n16919 & n16975 ) | ( ~n16919 & n16976 ) | ( n16975 & n16976 ) ;
  assign n16978 = ( n16844 & n16909 ) | ( n16844 & ~n16977 ) | ( n16909 & ~n16977 ) ;
  assign n16979 = ( ~n16844 & n16909 ) | ( ~n16844 & n16977 ) | ( n16909 & n16977 ) ;
  assign n16980 = ( ~n16909 & n16978 ) | ( ~n16909 & n16979 ) | ( n16978 & n16979 ) ;
  assign n16981 = ( n16847 & n16899 ) | ( n16847 & ~n16980 ) | ( n16899 & ~n16980 ) ;
  assign n16982 = ( ~n16847 & n16899 ) | ( ~n16847 & n16980 ) | ( n16899 & n16980 ) ;
  assign n16983 = ( ~n16899 & n16981 ) | ( ~n16899 & n16982 ) | ( n16981 & n16982 ) ;
  assign n16984 = ( n16851 & n16889 ) | ( n16851 & ~n16983 ) | ( n16889 & ~n16983 ) ;
  assign n16985 = ( ~n16851 & n16889 ) | ( ~n16851 & n16983 ) | ( n16889 & n16983 ) ;
  assign n16986 = ( ~n16889 & n16984 ) | ( ~n16889 & n16985 ) | ( n16984 & n16985 ) ;
  assign n16987 = ( ~n16854 & n16879 ) | ( ~n16854 & n16986 ) | ( n16879 & n16986 ) ;
  assign n16988 = ( n16854 & n16879 ) | ( n16854 & ~n16986 ) | ( n16879 & ~n16986 ) ;
  assign n16989 = ( ~n16879 & n16987 ) | ( ~n16879 & n16988 ) | ( n16987 & n16988 ) ;
  assign n16990 = ( n16866 & n16869 ) | ( n16866 & ~n16989 ) | ( n16869 & ~n16989 ) ;
  assign n16991 = ( ~n16866 & n16869 ) | ( ~n16866 & n16989 ) | ( n16869 & n16989 ) ;
  assign n16992 = ( ~n16869 & n16990 ) | ( ~n16869 & n16991 ) | ( n16990 & n16991 ) ;
  assign n16993 = n4020 & n9038 ;
  assign n16994 = x41 & n16993 ;
  assign n16995 = x126 & n4027 ;
  assign n16996 = x125 & n4024 ;
  assign n16997 = n16995 | n16996 ;
  assign n16998 = x124 & n4223 ;
  assign n16999 = n16997 | n16998 ;
  assign n17000 = ( ~x41 & n16993 ) | ( ~x41 & n16999 ) | ( n16993 & n16999 ) ;
  assign n17001 = x41 & ~n16999 ;
  assign n17002 = ( ~n16994 & n17000 ) | ( ~n16994 & n17001 ) | ( n17000 & n17001 ) ;
  assign n17003 = n4625 & n8461 ;
  assign n17004 = x44 & n17003 ;
  assign n17005 = x123 & n4791 ;
  assign n17006 = x122 & n4621 ;
  assign n17007 = n17005 | n17006 ;
  assign n17008 = x121 & n4795 ;
  assign n17009 = n17007 | n17008 ;
  assign n17010 = ( ~x44 & n17003 ) | ( ~x44 & n17009 ) | ( n17003 & n17009 ) ;
  assign n17011 = x44 & ~n17009 ;
  assign n17012 = ( ~n17004 & n17010 ) | ( ~n17004 & n17011 ) | ( n17010 & n17011 ) ;
  assign n17013 = n5223 & n7444 ;
  assign n17014 = x47 & n17013 ;
  assign n17015 = x120 & n5230 ;
  assign n17016 = x119 & n5227 ;
  assign n17017 = n17015 | n17016 ;
  assign n17018 = x118 & n5434 ;
  assign n17019 = n17017 | n17018 ;
  assign n17020 = ( ~x47 & n17013 ) | ( ~x47 & n17019 ) | ( n17013 & n17019 ) ;
  assign n17021 = x47 & ~n17019 ;
  assign n17022 = ( ~n17014 & n17020 ) | ( ~n17014 & n17021 ) | ( n17020 & n17021 ) ;
  assign n17023 = n5858 & n6924 ;
  assign n17024 = x50 & n17023 ;
  assign n17025 = x117 & n5865 ;
  assign n17026 = x116 & n5862 ;
  assign n17027 = n17025 | n17026 ;
  assign n17028 = x115 & n6092 ;
  assign n17029 = n17027 | n17028 ;
  assign n17030 = ( ~x50 & n17023 ) | ( ~x50 & n17029 ) | ( n17023 & n17029 ) ;
  assign n17031 = x50 & ~n17029 ;
  assign n17032 = ( ~n17024 & n17030 ) | ( ~n17024 & n17031 ) | ( n17030 & n17031 ) ;
  assign n17033 = n6002 & n6546 ;
  assign n17034 = x53 & n17033 ;
  assign n17035 = x114 & n6553 ;
  assign n17036 = x113 & n6550 ;
  assign n17037 = n17035 | n17036 ;
  assign n17038 = x112 & n6787 ;
  assign n17039 = n17037 | n17038 ;
  assign n17040 = ( ~x53 & n17033 ) | ( ~x53 & n17039 ) | ( n17033 & n17039 ) ;
  assign n17041 = x53 & ~n17039 ;
  assign n17042 = ( ~n17034 & n17040 ) | ( ~n17034 & n17041 ) | ( n17040 & n17041 ) ;
  assign n17043 = n5347 & n7277 ;
  assign n17044 = x56 & n17043 ;
  assign n17045 = x111 & n7545 ;
  assign n17046 = x110 & n7273 ;
  assign n17047 = n17045 | n17046 ;
  assign n17048 = x109 & n7552 ;
  assign n17049 = n17047 | n17048 ;
  assign n17050 = ( ~x56 & n17043 ) | ( ~x56 & n17049 ) | ( n17043 & n17049 ) ;
  assign n17051 = x56 & ~n17049 ;
  assign n17052 = ( ~n17044 & n17050 ) | ( ~n17044 & n17051 ) | ( n17050 & n17051 ) ;
  assign n17053 = n4914 & n8067 ;
  assign n17054 = x59 & n17053 ;
  assign n17055 = x108 & n8074 ;
  assign n17056 = x107 & n8071 ;
  assign n17057 = n17055 | n17056 ;
  assign n17058 = x106 & n8298 ;
  assign n17059 = n17057 | n17058 ;
  assign n17060 = ( ~x59 & n17053 ) | ( ~x59 & n17059 ) | ( n17053 & n17059 ) ;
  assign n17061 = x59 & ~n17059 ;
  assign n17062 = ( ~n17054 & n17060 ) | ( ~n17054 & n17061 ) | ( n17060 & n17061 ) ;
  assign n17063 = n4145 & n8859 ;
  assign n17064 = x62 & n17063 ;
  assign n17065 = x105 & n8866 ;
  assign n17066 = x104 & n8863 ;
  assign n17067 = n17065 | n17066 ;
  assign n17068 = x103 & n9125 ;
  assign n17069 = n17067 | n17068 ;
  assign n17070 = ( ~x62 & n17063 ) | ( ~x62 & n17069 ) | ( n17063 & n17069 ) ;
  assign n17071 = x62 & ~n17069 ;
  assign n17072 = ( ~n17064 & n17070 ) | ( ~n17064 & n17071 ) | ( n17070 & n17071 ) ;
  assign n17073 = ( x62 & x63 ) | ( x62 & x102 ) | ( x63 & x102 ) ;
  assign n17074 = ( x62 & x101 ) | ( x62 & ~n9394 ) | ( x101 & ~n9394 ) ;
  assign n17075 = ( x101 & n17073 ) | ( x101 & ~n17074 ) | ( n17073 & ~n17074 ) ;
  assign n17076 = ( ~n16830 & n16962 ) | ( ~n16830 & n17075 ) | ( n16962 & n17075 ) ;
  assign n17077 = ( n16830 & ~n16952 ) | ( n16830 & n17076 ) | ( ~n16952 & n17076 ) ;
  assign n17078 = ( n16830 & n16963 ) | ( n16830 & n17075 ) | ( n16963 & n17075 ) ;
  assign n17079 = ( n16952 & n17077 ) | ( n16952 & ~n17078 ) | ( n17077 & ~n17078 ) ;
  assign n17080 = ( n17062 & n17072 ) | ( n17062 & ~n17079 ) | ( n17072 & ~n17079 ) ;
  assign n17081 = ( n17062 & ~n17072 ) | ( n17062 & n17079 ) | ( ~n17072 & n17079 ) ;
  assign n17082 = ( ~n17062 & n17080 ) | ( ~n17062 & n17081 ) | ( n17080 & n17081 ) ;
  assign n17083 = ( n16966 & n17052 ) | ( n16966 & ~n17082 ) | ( n17052 & ~n17082 ) ;
  assign n17084 = ( ~n16966 & n17052 ) | ( ~n16966 & n17082 ) | ( n17052 & n17082 ) ;
  assign n17085 = ( ~n17052 & n17083 ) | ( ~n17052 & n17084 ) | ( n17083 & n17084 ) ;
  assign n17086 = ( n16969 & n17042 ) | ( n16969 & ~n17085 ) | ( n17042 & ~n17085 ) ;
  assign n17087 = ( ~n16969 & n17042 ) | ( ~n16969 & n17085 ) | ( n17042 & n17085 ) ;
  assign n17088 = ( ~n17042 & n17086 ) | ( ~n17042 & n17087 ) | ( n17086 & n17087 ) ;
  assign n17089 = ( n16972 & n17032 ) | ( n16972 & ~n17088 ) | ( n17032 & ~n17088 ) ;
  assign n17090 = ( ~n16972 & n17032 ) | ( ~n16972 & n17088 ) | ( n17032 & n17088 ) ;
  assign n17091 = ( ~n17032 & n17089 ) | ( ~n17032 & n17090 ) | ( n17089 & n17090 ) ;
  assign n17092 = ( n16975 & n17022 ) | ( n16975 & ~n17091 ) | ( n17022 & ~n17091 ) ;
  assign n17093 = ( ~n16975 & n17022 ) | ( ~n16975 & n17091 ) | ( n17022 & n17091 ) ;
  assign n17094 = ( ~n17022 & n17092 ) | ( ~n17022 & n17093 ) | ( n17092 & n17093 ) ;
  assign n17095 = ( n16978 & n17012 ) | ( n16978 & ~n17094 ) | ( n17012 & ~n17094 ) ;
  assign n17096 = ( ~n16978 & n17012 ) | ( ~n16978 & n17094 ) | ( n17012 & n17094 ) ;
  assign n17097 = ( ~n17012 & n17095 ) | ( ~n17012 & n17096 ) | ( n17095 & n17096 ) ;
  assign n17098 = ( n16981 & n17002 ) | ( n16981 & ~n17097 ) | ( n17002 & ~n17097 ) ;
  assign n17099 = ( ~n16981 & n17002 ) | ( ~n16981 & n17097 ) | ( n17002 & n17097 ) ;
  assign n17100 = ( ~n17002 & n17098 ) | ( ~n17002 & n17099 ) | ( n17098 & n17099 ) ;
  assign n17101 = x127 & n3662 ;
  assign n17102 = n3492 | n17101 ;
  assign n17103 = ( n9865 & n17101 ) | ( n9865 & n17102 ) | ( n17101 & n17102 ) ;
  assign n17104 = x38 & ~n17103 ;
  assign n17105 = ~x38 & n17103 ;
  assign n17106 = n17104 | n17105 ;
  assign n17107 = ( n16984 & ~n17100 ) | ( n16984 & n17106 ) | ( ~n17100 & n17106 ) ;
  assign n17108 = ( n16984 & n17100 ) | ( n16984 & n17106 ) | ( n17100 & n17106 ) ;
  assign n17109 = ( n17100 & n17107 ) | ( n17100 & ~n17108 ) | ( n17107 & ~n17108 ) ;
  assign n17110 = ( ~n16988 & n16991 ) | ( ~n16988 & n17109 ) | ( n16991 & n17109 ) ;
  assign n17111 = ( n16988 & n16991 ) | ( n16988 & ~n17109 ) | ( n16991 & ~n17109 ) ;
  assign n17112 = ( ~n16991 & n17110 ) | ( ~n16991 & n17111 ) | ( n17110 & n17111 ) ;
  assign n17113 = n4625 & n8729 ;
  assign n17114 = x44 & n17113 ;
  assign n17115 = x124 & n4791 ;
  assign n17116 = x123 & n4621 ;
  assign n17117 = n17115 | n17116 ;
  assign n17118 = x122 & n4795 ;
  assign n17119 = n17117 | n17118 ;
  assign n17120 = ( ~x44 & n17113 ) | ( ~x44 & n17119 ) | ( n17113 & n17119 ) ;
  assign n17121 = x44 & ~n17119 ;
  assign n17122 = ( ~n17114 & n17120 ) | ( ~n17114 & n17121 ) | ( n17120 & n17121 ) ;
  assign n17123 = n5223 & n7696 ;
  assign n17124 = x47 & n17123 ;
  assign n17125 = x121 & n5230 ;
  assign n17126 = x120 & n5227 ;
  assign n17127 = n17125 | n17126 ;
  assign n17128 = x119 & n5434 ;
  assign n17129 = n17127 | n17128 ;
  assign n17130 = ( ~x47 & n17123 ) | ( ~x47 & n17129 ) | ( n17123 & n17129 ) ;
  assign n17131 = x47 & ~n17129 ;
  assign n17132 = ( ~n17124 & n17130 ) | ( ~n17124 & n17131 ) | ( n17130 & n17131 ) ;
  assign n17133 = n5858 & n6940 ;
  assign n17134 = x50 & n17133 ;
  assign n17135 = x118 & n5865 ;
  assign n17136 = x117 & n5862 ;
  assign n17137 = n17135 | n17136 ;
  assign n17138 = x116 & n6092 ;
  assign n17139 = n17137 | n17138 ;
  assign n17140 = ( ~x50 & n17133 ) | ( ~x50 & n17139 ) | ( n17133 & n17139 ) ;
  assign n17141 = x50 & ~n17139 ;
  assign n17142 = ( ~n17134 & n17140 ) | ( ~n17134 & n17141 ) | ( n17140 & n17141 ) ;
  assign n17143 = n6446 & n6546 ;
  assign n17144 = x53 & n17143 ;
  assign n17145 = x115 & n6553 ;
  assign n17146 = x114 & n6550 ;
  assign n17147 = n17145 | n17146 ;
  assign n17148 = x113 & n6787 ;
  assign n17149 = n17147 | n17148 ;
  assign n17150 = ( ~x53 & n17143 ) | ( ~x53 & n17149 ) | ( n17143 & n17149 ) ;
  assign n17151 = x53 & ~n17149 ;
  assign n17152 = ( ~n17144 & n17150 ) | ( ~n17144 & n17151 ) | ( n17150 & n17151 ) ;
  assign n17153 = n5558 & n7277 ;
  assign n17154 = x56 & n17153 ;
  assign n17155 = x112 & n7545 ;
  assign n17156 = x111 & n7273 ;
  assign n17157 = n17155 | n17156 ;
  assign n17158 = x110 & n7552 ;
  assign n17159 = n17157 | n17158 ;
  assign n17160 = ( ~x56 & n17153 ) | ( ~x56 & n17159 ) | ( n17153 & n17159 ) ;
  assign n17161 = x56 & ~n17159 ;
  assign n17162 = ( ~n17154 & n17160 ) | ( ~n17154 & n17161 ) | ( n17160 & n17161 ) ;
  assign n17163 = n4930 & n8067 ;
  assign n17164 = x59 & n17163 ;
  assign n17165 = x109 & n8074 ;
  assign n17166 = x108 & n8071 ;
  assign n17167 = n17165 | n17166 ;
  assign n17168 = x107 & n8298 ;
  assign n17169 = n17167 | n17168 ;
  assign n17170 = ( ~x59 & n17163 ) | ( ~x59 & n17169 ) | ( n17163 & n17169 ) ;
  assign n17171 = x59 & ~n17169 ;
  assign n17172 = ( ~n17164 & n17170 ) | ( ~n17164 & n17171 ) | ( n17170 & n17171 ) ;
  assign n17173 = n4331 & n8859 ;
  assign n17174 = x62 & n17173 ;
  assign n17175 = x106 & n8866 ;
  assign n17176 = x105 & n8863 ;
  assign n17177 = n17175 | n17176 ;
  assign n17178 = x104 & n9125 ;
  assign n17179 = n17177 | n17178 ;
  assign n17180 = ( ~x62 & n17173 ) | ( ~x62 & n17179 ) | ( n17173 & n17179 ) ;
  assign n17181 = x62 & ~n17179 ;
  assign n17182 = ( ~n17174 & n17180 ) | ( ~n17174 & n17181 ) | ( n17180 & n17181 ) ;
  assign n17183 = ( x62 & x63 ) | ( x62 & x103 ) | ( x63 & x103 ) ;
  assign n17184 = ( x62 & x102 ) | ( x62 & ~n9394 ) | ( x102 & ~n9394 ) ;
  assign n17185 = ( x102 & n17183 ) | ( x102 & ~n17184 ) | ( n17183 & ~n17184 ) ;
  assign n17186 = ( x38 & n16952 ) | ( x38 & n17185 ) | ( n16952 & n17185 ) ;
  assign n17187 = ( ~x38 & n16952 ) | ( ~x38 & n17185 ) | ( n16952 & n17185 ) ;
  assign n17188 = ( x38 & ~n17186 ) | ( x38 & n17187 ) | ( ~n17186 & n17187 ) ;
  assign n17189 = ( n17077 & n17182 ) | ( n17077 & ~n17188 ) | ( n17182 & ~n17188 ) ;
  assign n17190 = ( n17077 & ~n17182 ) | ( n17077 & n17188 ) | ( ~n17182 & n17188 ) ;
  assign n17191 = ( ~n17077 & n17189 ) | ( ~n17077 & n17190 ) | ( n17189 & n17190 ) ;
  assign n17192 = ( n17080 & n17172 ) | ( n17080 & ~n17191 ) | ( n17172 & ~n17191 ) ;
  assign n17193 = ( n17080 & ~n17172 ) | ( n17080 & n17191 ) | ( ~n17172 & n17191 ) ;
  assign n17194 = ( ~n17080 & n17192 ) | ( ~n17080 & n17193 ) | ( n17192 & n17193 ) ;
  assign n17195 = ( n17083 & n17162 ) | ( n17083 & ~n17194 ) | ( n17162 & ~n17194 ) ;
  assign n17196 = ( n17083 & ~n17162 ) | ( n17083 & n17194 ) | ( ~n17162 & n17194 ) ;
  assign n17197 = ( ~n17083 & n17195 ) | ( ~n17083 & n17196 ) | ( n17195 & n17196 ) ;
  assign n17198 = ( n17086 & n17152 ) | ( n17086 & ~n17197 ) | ( n17152 & ~n17197 ) ;
  assign n17199 = ( n17086 & ~n17152 ) | ( n17086 & n17197 ) | ( ~n17152 & n17197 ) ;
  assign n17200 = ( ~n17086 & n17198 ) | ( ~n17086 & n17199 ) | ( n17198 & n17199 ) ;
  assign n17201 = ( n17089 & n17142 ) | ( n17089 & ~n17200 ) | ( n17142 & ~n17200 ) ;
  assign n17202 = ( n17089 & ~n17142 ) | ( n17089 & n17200 ) | ( ~n17142 & n17200 ) ;
  assign n17203 = ( ~n17089 & n17201 ) | ( ~n17089 & n17202 ) | ( n17201 & n17202 ) ;
  assign n17204 = ( n17092 & n17132 ) | ( n17092 & ~n17203 ) | ( n17132 & ~n17203 ) ;
  assign n17205 = ( n17092 & ~n17132 ) | ( n17092 & n17203 ) | ( ~n17132 & n17203 ) ;
  assign n17206 = ( ~n17092 & n17204 ) | ( ~n17092 & n17205 ) | ( n17204 & n17205 ) ;
  assign n17207 = ( n17095 & n17122 ) | ( n17095 & ~n17206 ) | ( n17122 & ~n17206 ) ;
  assign n17208 = ( n17095 & ~n17122 ) | ( n17095 & n17206 ) | ( ~n17122 & n17206 ) ;
  assign n17209 = ( ~n17095 & n17207 ) | ( ~n17095 & n17208 ) | ( n17207 & n17208 ) ;
  assign n17210 = n4020 & n9576 ;
  assign n17211 = x41 & n17210 ;
  assign n17212 = x127 & n4027 ;
  assign n17213 = x126 & n4024 ;
  assign n17214 = n17212 | n17213 ;
  assign n17215 = x125 & n4223 ;
  assign n17216 = n17214 | n17215 ;
  assign n17217 = ( ~x41 & n17210 ) | ( ~x41 & n17216 ) | ( n17210 & n17216 ) ;
  assign n17218 = x41 & ~n17216 ;
  assign n17219 = ( ~n17211 & n17217 ) | ( ~n17211 & n17218 ) | ( n17217 & n17218 ) ;
  assign n17220 = ( n17098 & ~n17209 ) | ( n17098 & n17219 ) | ( ~n17209 & n17219 ) ;
  assign n17221 = ( n17098 & n17209 ) | ( n17098 & ~n17219 ) | ( n17209 & ~n17219 ) ;
  assign n17222 = ( ~n17098 & n17220 ) | ( ~n17098 & n17221 ) | ( n17220 & n17221 ) ;
  assign n17223 = ( ~n17107 & n17110 ) | ( ~n17107 & n17222 ) | ( n17110 & n17222 ) ;
  assign n17224 = ( n17107 & n17110 ) | ( n17107 & ~n17222 ) | ( n17110 & ~n17222 ) ;
  assign n17225 = ( ~n17110 & n17223 ) | ( ~n17110 & n17224 ) | ( n17223 & n17224 ) ;
  assign n17226 = x126 & n4223 ;
  assign n17227 = x41 & n17226 ;
  assign n17228 = x127 & n4024 ;
  assign n17229 = n4020 | n17228 ;
  assign n17230 = ( n9867 & n17228 ) | ( n9867 & n17229 ) | ( n17228 & n17229 ) ;
  assign n17231 = ( ~x41 & n17226 ) | ( ~x41 & n17230 ) | ( n17226 & n17230 ) ;
  assign n17232 = x41 & ~n17230 ;
  assign n17233 = ( ~n17227 & n17231 ) | ( ~n17227 & n17232 ) | ( n17231 & n17232 ) ;
  assign n17234 = n4625 & n9009 ;
  assign n17235 = x44 & n17234 ;
  assign n17236 = x125 & n4791 ;
  assign n17237 = x124 & n4621 ;
  assign n17238 = n17236 | n17237 ;
  assign n17239 = x123 & n4795 ;
  assign n17240 = n17238 | n17239 ;
  assign n17241 = ( ~x44 & n17234 ) | ( ~x44 & n17240 ) | ( n17234 & n17240 ) ;
  assign n17242 = x44 & ~n17240 ;
  assign n17243 = ( ~n17235 & n17241 ) | ( ~n17235 & n17242 ) | ( n17241 & n17242 ) ;
  assign n17244 = n5223 & n8207 ;
  assign n17245 = x47 & n17244 ;
  assign n17246 = x122 & n5230 ;
  assign n17247 = x121 & n5227 ;
  assign n17248 = n17246 | n17247 ;
  assign n17249 = x120 & n5434 ;
  assign n17250 = n17248 | n17249 ;
  assign n17251 = ( ~x47 & n17244 ) | ( ~x47 & n17250 ) | ( n17244 & n17250 ) ;
  assign n17252 = x47 & ~n17250 ;
  assign n17253 = ( ~n17245 & n17251 ) | ( ~n17245 & n17252 ) | ( n17251 & n17252 ) ;
  assign n17254 = n5858 & n7181 ;
  assign n17255 = x50 & n17254 ;
  assign n17256 = x119 & n5865 ;
  assign n17257 = x118 & n5862 ;
  assign n17258 = n17256 | n17257 ;
  assign n17259 = x117 & n6092 ;
  assign n17260 = n17258 | n17259 ;
  assign n17261 = ( ~x50 & n17254 ) | ( ~x50 & n17260 ) | ( n17254 & n17260 ) ;
  assign n17262 = x50 & ~n17260 ;
  assign n17263 = ( ~n17255 & n17261 ) | ( ~n17255 & n17262 ) | ( n17261 & n17262 ) ;
  assign n17264 = n6462 & n6546 ;
  assign n17265 = x53 & n17264 ;
  assign n17266 = x116 & n6553 ;
  assign n17267 = x115 & n6550 ;
  assign n17268 = n17266 | n17267 ;
  assign n17269 = x114 & n6787 ;
  assign n17270 = n17268 | n17269 ;
  assign n17271 = ( ~x53 & n17264 ) | ( ~x53 & n17270 ) | ( n17264 & n17270 ) ;
  assign n17272 = x53 & ~n17270 ;
  assign n17273 = ( ~n17265 & n17271 ) | ( ~n17265 & n17272 ) | ( n17271 & n17272 ) ;
  assign n17274 = n5774 & n7277 ;
  assign n17275 = x56 & n17274 ;
  assign n17276 = x113 & n7545 ;
  assign n17277 = x112 & n7273 ;
  assign n17278 = n17276 | n17277 ;
  assign n17279 = x111 & n7552 ;
  assign n17280 = n17278 | n17279 ;
  assign n17281 = ( ~x56 & n17274 ) | ( ~x56 & n17280 ) | ( n17274 & n17280 ) ;
  assign n17282 = x56 & ~n17280 ;
  assign n17283 = ( ~n17275 & n17281 ) | ( ~n17275 & n17282 ) | ( n17281 & n17282 ) ;
  assign n17284 = n5331 & n8067 ;
  assign n17285 = x59 & n17284 ;
  assign n17286 = x110 & n8074 ;
  assign n17287 = x109 & n8071 ;
  assign n17288 = n17286 | n17287 ;
  assign n17289 = x108 & n8298 ;
  assign n17290 = n17288 | n17289 ;
  assign n17291 = ( ~x59 & n17284 ) | ( ~x59 & n17290 ) | ( n17284 & n17290 ) ;
  assign n17292 = x59 & ~n17290 ;
  assign n17293 = ( ~n17285 & n17291 ) | ( ~n17285 & n17292 ) | ( n17291 & n17292 ) ;
  assign n17294 = ( x62 & x63 ) | ( x62 & x104 ) | ( x63 & x104 ) ;
  assign n17295 = ( x62 & x103 ) | ( x62 & ~n9394 ) | ( x103 & ~n9394 ) ;
  assign n17296 = ( x103 & n17294 ) | ( x103 & ~n17295 ) | ( n17294 & ~n17295 ) ;
  assign n17297 = n4523 & n8859 ;
  assign n17298 = x62 & n17297 ;
  assign n17299 = x107 & n8866 ;
  assign n17300 = x106 & n8863 ;
  assign n17301 = n17299 | n17300 ;
  assign n17302 = x105 & n9125 ;
  assign n17303 = n17301 | n17302 ;
  assign n17304 = ( ~x62 & n17297 ) | ( ~x62 & n17303 ) | ( n17297 & n17303 ) ;
  assign n17305 = x62 & ~n17303 ;
  assign n17306 = ( ~n17298 & n17304 ) | ( ~n17298 & n17305 ) | ( n17304 & n17305 ) ;
  assign n17307 = ( ~n17187 & n17296 ) | ( ~n17187 & n17306 ) | ( n17296 & n17306 ) ;
  assign n17308 = ( n17187 & n17296 ) | ( n17187 & ~n17306 ) | ( n17296 & ~n17306 ) ;
  assign n17309 = ( ~n17296 & n17307 ) | ( ~n17296 & n17308 ) | ( n17307 & n17308 ) ;
  assign n17310 = ( n17189 & n17293 ) | ( n17189 & ~n17309 ) | ( n17293 & ~n17309 ) ;
  assign n17311 = ( ~n17189 & n17293 ) | ( ~n17189 & n17309 ) | ( n17293 & n17309 ) ;
  assign n17312 = ( ~n17293 & n17310 ) | ( ~n17293 & n17311 ) | ( n17310 & n17311 ) ;
  assign n17313 = ( n17192 & n17283 ) | ( n17192 & ~n17312 ) | ( n17283 & ~n17312 ) ;
  assign n17314 = ( ~n17192 & n17283 ) | ( ~n17192 & n17312 ) | ( n17283 & n17312 ) ;
  assign n17315 = ( ~n17283 & n17313 ) | ( ~n17283 & n17314 ) | ( n17313 & n17314 ) ;
  assign n17316 = ( n17195 & n17273 ) | ( n17195 & ~n17315 ) | ( n17273 & ~n17315 ) ;
  assign n17317 = ( ~n17195 & n17273 ) | ( ~n17195 & n17315 ) | ( n17273 & n17315 ) ;
  assign n17318 = ( ~n17273 & n17316 ) | ( ~n17273 & n17317 ) | ( n17316 & n17317 ) ;
  assign n17319 = ( n17198 & n17263 ) | ( n17198 & ~n17318 ) | ( n17263 & ~n17318 ) ;
  assign n17320 = ( ~n17198 & n17263 ) | ( ~n17198 & n17318 ) | ( n17263 & n17318 ) ;
  assign n17321 = ( ~n17263 & n17319 ) | ( ~n17263 & n17320 ) | ( n17319 & n17320 ) ;
  assign n17322 = ( n17201 & n17253 ) | ( n17201 & ~n17321 ) | ( n17253 & ~n17321 ) ;
  assign n17323 = ( ~n17201 & n17253 ) | ( ~n17201 & n17321 ) | ( n17253 & n17321 ) ;
  assign n17324 = ( ~n17253 & n17322 ) | ( ~n17253 & n17323 ) | ( n17322 & n17323 ) ;
  assign n17325 = ( ~n17204 & n17243 ) | ( ~n17204 & n17324 ) | ( n17243 & n17324 ) ;
  assign n17326 = ( n17204 & n17243 ) | ( n17204 & ~n17324 ) | ( n17243 & ~n17324 ) ;
  assign n17327 = ( ~n17243 & n17325 ) | ( ~n17243 & n17326 ) | ( n17325 & n17326 ) ;
  assign n17328 = ( ~n17207 & n17233 ) | ( ~n17207 & n17327 ) | ( n17233 & n17327 ) ;
  assign n17329 = ( n17207 & n17233 ) | ( n17207 & ~n17327 ) | ( n17233 & ~n17327 ) ;
  assign n17330 = ( ~n17233 & n17328 ) | ( ~n17233 & n17329 ) | ( n17328 & n17329 ) ;
  assign n17331 = ( ~n17220 & n17223 ) | ( ~n17220 & n17330 ) | ( n17223 & n17330 ) ;
  assign n17332 = ( n17220 & n17223 ) | ( n17220 & ~n17330 ) | ( n17223 & ~n17330 ) ;
  assign n17333 = ( ~n17223 & n17331 ) | ( ~n17223 & n17332 ) | ( n17331 & n17332 ) ;
  assign n17334 = n4625 & n9038 ;
  assign n17335 = x44 & n17334 ;
  assign n17336 = x126 & n4791 ;
  assign n17337 = x125 & n4621 ;
  assign n17338 = n17336 | n17337 ;
  assign n17339 = x124 & n4795 ;
  assign n17340 = n17338 | n17339 ;
  assign n17341 = ( ~x44 & n17334 ) | ( ~x44 & n17340 ) | ( n17334 & n17340 ) ;
  assign n17342 = x44 & ~n17340 ;
  assign n17343 = ( ~n17335 & n17341 ) | ( ~n17335 & n17342 ) | ( n17341 & n17342 ) ;
  assign n17344 = n5223 & n8461 ;
  assign n17345 = x47 & n17344 ;
  assign n17346 = x123 & n5230 ;
  assign n17347 = x122 & n5227 ;
  assign n17348 = n17346 | n17347 ;
  assign n17349 = x121 & n5434 ;
  assign n17350 = n17348 | n17349 ;
  assign n17351 = ( ~x47 & n17344 ) | ( ~x47 & n17350 ) | ( n17344 & n17350 ) ;
  assign n17352 = x47 & ~n17350 ;
  assign n17353 = ( ~n17345 & n17351 ) | ( ~n17345 & n17352 ) | ( n17351 & n17352 ) ;
  assign n17354 = n5858 & n7444 ;
  assign n17355 = x50 & n17354 ;
  assign n17356 = x120 & n5865 ;
  assign n17357 = x119 & n5862 ;
  assign n17358 = n17356 | n17357 ;
  assign n17359 = x118 & n6092 ;
  assign n17360 = n17358 | n17359 ;
  assign n17361 = ( ~x50 & n17354 ) | ( ~x50 & n17360 ) | ( n17354 & n17360 ) ;
  assign n17362 = x50 & ~n17360 ;
  assign n17363 = ( ~n17355 & n17361 ) | ( ~n17355 & n17362 ) | ( n17361 & n17362 ) ;
  assign n17364 = n6546 & n6924 ;
  assign n17365 = x53 & n17364 ;
  assign n17366 = x117 & n6553 ;
  assign n17367 = x116 & n6550 ;
  assign n17368 = n17366 | n17367 ;
  assign n17369 = x115 & n6787 ;
  assign n17370 = n17368 | n17369 ;
  assign n17371 = ( ~x53 & n17364 ) | ( ~x53 & n17370 ) | ( n17364 & n17370 ) ;
  assign n17372 = x53 & ~n17370 ;
  assign n17373 = ( ~n17365 & n17371 ) | ( ~n17365 & n17372 ) | ( n17371 & n17372 ) ;
  assign n17374 = n6002 & n7277 ;
  assign n17375 = x56 & n17374 ;
  assign n17376 = x114 & n7545 ;
  assign n17377 = x113 & n7273 ;
  assign n17378 = n17376 | n17377 ;
  assign n17379 = x112 & n7552 ;
  assign n17380 = n17378 | n17379 ;
  assign n17381 = ( ~x56 & n17374 ) | ( ~x56 & n17380 ) | ( n17374 & n17380 ) ;
  assign n17382 = x56 & ~n17380 ;
  assign n17383 = ( ~n17375 & n17381 ) | ( ~n17375 & n17382 ) | ( n17381 & n17382 ) ;
  assign n17384 = n5347 & n8067 ;
  assign n17385 = x59 & n17384 ;
  assign n17386 = x111 & n8074 ;
  assign n17387 = x110 & n8071 ;
  assign n17388 = n17386 | n17387 ;
  assign n17389 = x109 & n8298 ;
  assign n17390 = n17388 | n17389 ;
  assign n17391 = ( ~x59 & n17384 ) | ( ~x59 & n17390 ) | ( n17384 & n17390 ) ;
  assign n17392 = x59 & ~n17390 ;
  assign n17393 = ( ~n17385 & n17391 ) | ( ~n17385 & n17392 ) | ( n17391 & n17392 ) ;
  assign n17394 = n4914 & n8859 ;
  assign n17395 = x62 & n17394 ;
  assign n17396 = x108 & n8866 ;
  assign n17397 = x107 & n8863 ;
  assign n17398 = n17396 | n17397 ;
  assign n17399 = x106 & n9125 ;
  assign n17400 = n17398 | n17399 ;
  assign n17401 = ( ~x62 & n17394 ) | ( ~x62 & n17400 ) | ( n17394 & n17400 ) ;
  assign n17402 = x62 & ~n17400 ;
  assign n17403 = ( ~n17395 & n17401 ) | ( ~n17395 & n17402 ) | ( n17401 & n17402 ) ;
  assign n17404 = ( x62 & x63 ) | ( x62 & x105 ) | ( x63 & x105 ) ;
  assign n17405 = ( x62 & x104 ) | ( x62 & ~n9394 ) | ( x104 & ~n9394 ) ;
  assign n17406 = ( x104 & n17404 ) | ( x104 & ~n17405 ) | ( n17404 & ~n17405 ) ;
  assign n17407 = ( ~n17187 & n17306 ) | ( ~n17187 & n17406 ) | ( n17306 & n17406 ) ;
  assign n17408 = ( n17187 & ~n17296 ) | ( n17187 & n17407 ) | ( ~n17296 & n17407 ) ;
  assign n17409 = ( n17187 & n17307 ) | ( n17187 & n17406 ) | ( n17307 & n17406 ) ;
  assign n17410 = ( n17296 & n17408 ) | ( n17296 & ~n17409 ) | ( n17408 & ~n17409 ) ;
  assign n17411 = ( n17393 & n17403 ) | ( n17393 & ~n17410 ) | ( n17403 & ~n17410 ) ;
  assign n17412 = ( n17393 & ~n17403 ) | ( n17393 & n17410 ) | ( ~n17403 & n17410 ) ;
  assign n17413 = ( ~n17393 & n17411 ) | ( ~n17393 & n17412 ) | ( n17411 & n17412 ) ;
  assign n17414 = ( n17310 & n17383 ) | ( n17310 & ~n17413 ) | ( n17383 & ~n17413 ) ;
  assign n17415 = ( ~n17310 & n17383 ) | ( ~n17310 & n17413 ) | ( n17383 & n17413 ) ;
  assign n17416 = ( ~n17383 & n17414 ) | ( ~n17383 & n17415 ) | ( n17414 & n17415 ) ;
  assign n17417 = ( ~n17313 & n17373 ) | ( ~n17313 & n17416 ) | ( n17373 & n17416 ) ;
  assign n17418 = ( n17313 & n17373 ) | ( n17313 & ~n17416 ) | ( n17373 & ~n17416 ) ;
  assign n17419 = ( ~n17373 & n17417 ) | ( ~n17373 & n17418 ) | ( n17417 & n17418 ) ;
  assign n17420 = ( n17316 & n17363 ) | ( n17316 & ~n17419 ) | ( n17363 & ~n17419 ) ;
  assign n17421 = ( ~n17316 & n17363 ) | ( ~n17316 & n17419 ) | ( n17363 & n17419 ) ;
  assign n17422 = ( ~n17363 & n17420 ) | ( ~n17363 & n17421 ) | ( n17420 & n17421 ) ;
  assign n17423 = ( n17319 & n17353 ) | ( n17319 & ~n17422 ) | ( n17353 & ~n17422 ) ;
  assign n17424 = ( ~n17319 & n17353 ) | ( ~n17319 & n17422 ) | ( n17353 & n17422 ) ;
  assign n17425 = ( ~n17353 & n17423 ) | ( ~n17353 & n17424 ) | ( n17423 & n17424 ) ;
  assign n17426 = ( n17322 & n17343 ) | ( n17322 & ~n17425 ) | ( n17343 & ~n17425 ) ;
  assign n17427 = ( ~n17322 & n17343 ) | ( ~n17322 & n17425 ) | ( n17343 & n17425 ) ;
  assign n17428 = ( ~n17343 & n17426 ) | ( ~n17343 & n17427 ) | ( n17426 & n17427 ) ;
  assign n17429 = x127 & n4223 ;
  assign n17430 = n4020 | n17429 ;
  assign n17431 = ( n9865 & n17429 ) | ( n9865 & n17430 ) | ( n17429 & n17430 ) ;
  assign n17432 = x41 & ~n17431 ;
  assign n17433 = ~x41 & n17431 ;
  assign n17434 = n17432 | n17433 ;
  assign n17435 = ( n17326 & ~n17428 ) | ( n17326 & n17434 ) | ( ~n17428 & n17434 ) ;
  assign n17436 = ( n17326 & n17428 ) | ( n17326 & n17434 ) | ( n17428 & n17434 ) ;
  assign n17437 = ( n17428 & n17435 ) | ( n17428 & ~n17436 ) | ( n17435 & ~n17436 ) ;
  assign n17438 = ( n17329 & n17331 ) | ( n17329 & ~n17437 ) | ( n17331 & ~n17437 ) ;
  assign n17439 = ( ~n17329 & n17331 ) | ( ~n17329 & n17437 ) | ( n17331 & n17437 ) ;
  assign n17440 = ( ~n17331 & n17438 ) | ( ~n17331 & n17439 ) | ( n17438 & n17439 ) ;
  assign n17441 = n5223 & n8729 ;
  assign n17442 = x47 & n17441 ;
  assign n17443 = x124 & n5230 ;
  assign n17444 = x123 & n5227 ;
  assign n17445 = n17443 | n17444 ;
  assign n17446 = x122 & n5434 ;
  assign n17447 = n17445 | n17446 ;
  assign n17448 = ( ~x47 & n17441 ) | ( ~x47 & n17447 ) | ( n17441 & n17447 ) ;
  assign n17449 = x47 & ~n17447 ;
  assign n17450 = ( ~n17442 & n17448 ) | ( ~n17442 & n17449 ) | ( n17448 & n17449 ) ;
  assign n17451 = n5858 & n7696 ;
  assign n17452 = x50 & n17451 ;
  assign n17453 = x121 & n5865 ;
  assign n17454 = x120 & n5862 ;
  assign n17455 = n17453 | n17454 ;
  assign n17456 = x119 & n6092 ;
  assign n17457 = n17455 | n17456 ;
  assign n17458 = ( ~x50 & n17451 ) | ( ~x50 & n17457 ) | ( n17451 & n17457 ) ;
  assign n17459 = x50 & ~n17457 ;
  assign n17460 = ( ~n17452 & n17458 ) | ( ~n17452 & n17459 ) | ( n17458 & n17459 ) ;
  assign n17461 = n6546 & n6940 ;
  assign n17462 = x53 & n17461 ;
  assign n17463 = x118 & n6553 ;
  assign n17464 = x117 & n6550 ;
  assign n17465 = n17463 | n17464 ;
  assign n17466 = x116 & n6787 ;
  assign n17467 = n17465 | n17466 ;
  assign n17468 = ( ~x53 & n17461 ) | ( ~x53 & n17467 ) | ( n17461 & n17467 ) ;
  assign n17469 = x53 & ~n17467 ;
  assign n17470 = ( ~n17462 & n17468 ) | ( ~n17462 & n17469 ) | ( n17468 & n17469 ) ;
  assign n17471 = n6446 & n7277 ;
  assign n17472 = x56 & n17471 ;
  assign n17473 = x115 & n7545 ;
  assign n17474 = x114 & n7273 ;
  assign n17475 = n17473 | n17474 ;
  assign n17476 = x113 & n7552 ;
  assign n17477 = n17475 | n17476 ;
  assign n17478 = ( ~x56 & n17471 ) | ( ~x56 & n17477 ) | ( n17471 & n17477 ) ;
  assign n17479 = x56 & ~n17477 ;
  assign n17480 = ( ~n17472 & n17478 ) | ( ~n17472 & n17479 ) | ( n17478 & n17479 ) ;
  assign n17481 = n5558 & n8067 ;
  assign n17482 = x59 & n17481 ;
  assign n17483 = x112 & n8074 ;
  assign n17484 = x111 & n8071 ;
  assign n17485 = n17483 | n17484 ;
  assign n17486 = x110 & n8298 ;
  assign n17487 = n17485 | n17486 ;
  assign n17488 = ( ~x59 & n17481 ) | ( ~x59 & n17487 ) | ( n17481 & n17487 ) ;
  assign n17489 = x59 & ~n17487 ;
  assign n17490 = ( ~n17482 & n17488 ) | ( ~n17482 & n17489 ) | ( n17488 & n17489 ) ;
  assign n17491 = n4930 & n8859 ;
  assign n17492 = x62 & n17491 ;
  assign n17493 = x109 & n8866 ;
  assign n17494 = x108 & n8863 ;
  assign n17495 = n17493 | n17494 ;
  assign n17496 = x107 & n9125 ;
  assign n17497 = n17495 | n17496 ;
  assign n17498 = ( ~x62 & n17491 ) | ( ~x62 & n17497 ) | ( n17491 & n17497 ) ;
  assign n17499 = x62 & ~n17497 ;
  assign n17500 = ( ~n17492 & n17498 ) | ( ~n17492 & n17499 ) | ( n17498 & n17499 ) ;
  assign n17501 = ( x62 & x63 ) | ( x62 & x106 ) | ( x63 & x106 ) ;
  assign n17502 = ( x62 & x105 ) | ( x62 & ~n9394 ) | ( x105 & ~n9394 ) ;
  assign n17503 = ( x105 & n17501 ) | ( x105 & ~n17502 ) | ( n17501 & ~n17502 ) ;
  assign n17504 = ( x41 & n17296 ) | ( x41 & n17503 ) | ( n17296 & n17503 ) ;
  assign n17505 = ( ~x41 & n17296 ) | ( ~x41 & n17503 ) | ( n17296 & n17503 ) ;
  assign n17506 = ( x41 & ~n17504 ) | ( x41 & n17505 ) | ( ~n17504 & n17505 ) ;
  assign n17507 = ( n17408 & n17500 ) | ( n17408 & ~n17506 ) | ( n17500 & ~n17506 ) ;
  assign n17508 = ( ~n17408 & n17500 ) | ( ~n17408 & n17506 ) | ( n17500 & n17506 ) ;
  assign n17509 = ( ~n17500 & n17507 ) | ( ~n17500 & n17508 ) | ( n17507 & n17508 ) ;
  assign n17510 = ( n17411 & n17490 ) | ( n17411 & ~n17509 ) | ( n17490 & ~n17509 ) ;
  assign n17511 = ( n17411 & ~n17490 ) | ( n17411 & n17509 ) | ( ~n17490 & n17509 ) ;
  assign n17512 = ( ~n17411 & n17510 ) | ( ~n17411 & n17511 ) | ( n17510 & n17511 ) ;
  assign n17513 = ( n17414 & n17480 ) | ( n17414 & ~n17512 ) | ( n17480 & ~n17512 ) ;
  assign n17514 = ( n17414 & ~n17480 ) | ( n17414 & n17512 ) | ( ~n17480 & n17512 ) ;
  assign n17515 = ( ~n17414 & n17513 ) | ( ~n17414 & n17514 ) | ( n17513 & n17514 ) ;
  assign n17516 = ( n17418 & ~n17470 ) | ( n17418 & n17515 ) | ( ~n17470 & n17515 ) ;
  assign n17517 = ( n17418 & n17470 ) | ( n17418 & ~n17515 ) | ( n17470 & ~n17515 ) ;
  assign n17518 = ( ~n17418 & n17516 ) | ( ~n17418 & n17517 ) | ( n17516 & n17517 ) ;
  assign n17519 = ( n17420 & n17460 ) | ( n17420 & ~n17518 ) | ( n17460 & ~n17518 ) ;
  assign n17520 = ( ~n17420 & n17460 ) | ( ~n17420 & n17518 ) | ( n17460 & n17518 ) ;
  assign n17521 = ( ~n17460 & n17519 ) | ( ~n17460 & n17520 ) | ( n17519 & n17520 ) ;
  assign n17522 = ( n17423 & n17450 ) | ( n17423 & ~n17521 ) | ( n17450 & ~n17521 ) ;
  assign n17523 = ( n17423 & ~n17450 ) | ( n17423 & n17521 ) | ( ~n17450 & n17521 ) ;
  assign n17524 = ( ~n17423 & n17522 ) | ( ~n17423 & n17523 ) | ( n17522 & n17523 ) ;
  assign n17525 = n4625 & n9576 ;
  assign n17526 = x44 & n17525 ;
  assign n17527 = x127 & n4791 ;
  assign n17528 = x126 & n4621 ;
  assign n17529 = n17527 | n17528 ;
  assign n17530 = x125 & n4795 ;
  assign n17531 = n17529 | n17530 ;
  assign n17532 = ( ~x44 & n17525 ) | ( ~x44 & n17531 ) | ( n17525 & n17531 ) ;
  assign n17533 = x44 & ~n17531 ;
  assign n17534 = ( ~n17526 & n17532 ) | ( ~n17526 & n17533 ) | ( n17532 & n17533 ) ;
  assign n17535 = ( n17426 & ~n17524 ) | ( n17426 & n17534 ) | ( ~n17524 & n17534 ) ;
  assign n17536 = ( n17426 & n17524 ) | ( n17426 & ~n17534 ) | ( n17524 & ~n17534 ) ;
  assign n17537 = ( ~n17426 & n17535 ) | ( ~n17426 & n17536 ) | ( n17535 & n17536 ) ;
  assign n17538 = ( ~n17435 & n17439 ) | ( ~n17435 & n17537 ) | ( n17439 & n17537 ) ;
  assign n17539 = ( n17435 & n17439 ) | ( n17435 & ~n17537 ) | ( n17439 & ~n17537 ) ;
  assign n17540 = ( ~n17439 & n17538 ) | ( ~n17439 & n17539 ) | ( n17538 & n17539 ) ;
  assign n17541 = x126 & n4795 ;
  assign n17542 = n4625 | n17541 ;
  assign n17543 = ( n9867 & n17541 ) | ( n9867 & n17542 ) | ( n17541 & n17542 ) ;
  assign n17544 = x127 & n4621 ;
  assign n17545 = ( ~x44 & n17543 ) | ( ~x44 & n17544 ) | ( n17543 & n17544 ) ;
  assign n17546 = ( x44 & ~n17543 ) | ( x44 & n17544 ) | ( ~n17543 & n17544 ) ;
  assign n17547 = ~n17544 & n17546 ;
  assign n17548 = n17545 | n17547 ;
  assign n17549 = n5223 & n9009 ;
  assign n17550 = x47 & n17549 ;
  assign n17551 = x125 & n5230 ;
  assign n17552 = x124 & n5227 ;
  assign n17553 = n17551 | n17552 ;
  assign n17554 = x123 & n5434 ;
  assign n17555 = n17553 | n17554 ;
  assign n17556 = ( ~x47 & n17549 ) | ( ~x47 & n17555 ) | ( n17549 & n17555 ) ;
  assign n17557 = x47 & ~n17555 ;
  assign n17558 = ( ~n17550 & n17556 ) | ( ~n17550 & n17557 ) | ( n17556 & n17557 ) ;
  assign n17559 = n5858 & n8207 ;
  assign n17560 = x50 & n17559 ;
  assign n17561 = x122 & n5865 ;
  assign n17562 = x121 & n5862 ;
  assign n17563 = n17561 | n17562 ;
  assign n17564 = x120 & n6092 ;
  assign n17565 = n17563 | n17564 ;
  assign n17566 = ( ~x50 & n17559 ) | ( ~x50 & n17565 ) | ( n17559 & n17565 ) ;
  assign n17567 = x50 & ~n17565 ;
  assign n17568 = ( ~n17560 & n17566 ) | ( ~n17560 & n17567 ) | ( n17566 & n17567 ) ;
  assign n17569 = n6546 & n7181 ;
  assign n17570 = x53 & n17569 ;
  assign n17571 = x119 & n6553 ;
  assign n17572 = x118 & n6550 ;
  assign n17573 = n17571 | n17572 ;
  assign n17574 = x117 & n6787 ;
  assign n17575 = n17573 | n17574 ;
  assign n17576 = ( ~x53 & n17569 ) | ( ~x53 & n17575 ) | ( n17569 & n17575 ) ;
  assign n17577 = x53 & ~n17575 ;
  assign n17578 = ( ~n17570 & n17576 ) | ( ~n17570 & n17577 ) | ( n17576 & n17577 ) ;
  assign n17579 = n6462 & n7277 ;
  assign n17580 = x56 & n17579 ;
  assign n17581 = x116 & n7545 ;
  assign n17582 = x115 & n7273 ;
  assign n17583 = n17581 | n17582 ;
  assign n17584 = x114 & n7552 ;
  assign n17585 = n17583 | n17584 ;
  assign n17586 = ( ~x56 & n17579 ) | ( ~x56 & n17585 ) | ( n17579 & n17585 ) ;
  assign n17587 = x56 & ~n17585 ;
  assign n17588 = ( ~n17580 & n17586 ) | ( ~n17580 & n17587 ) | ( n17586 & n17587 ) ;
  assign n17589 = n5774 & n8067 ;
  assign n17590 = x59 & n17589 ;
  assign n17591 = x113 & n8074 ;
  assign n17592 = x112 & n8071 ;
  assign n17593 = n17591 | n17592 ;
  assign n17594 = x111 & n8298 ;
  assign n17595 = n17593 | n17594 ;
  assign n17596 = ( ~x59 & n17589 ) | ( ~x59 & n17595 ) | ( n17589 & n17595 ) ;
  assign n17597 = x59 & ~n17595 ;
  assign n17598 = ( ~n17590 & n17596 ) | ( ~n17590 & n17597 ) | ( n17596 & n17597 ) ;
  assign n17599 = n5331 & n8859 ;
  assign n17600 = x62 & n17599 ;
  assign n17601 = x110 & n8866 ;
  assign n17602 = x109 & n8863 ;
  assign n17603 = n17601 | n17602 ;
  assign n17604 = x108 & n9125 ;
  assign n17605 = n17603 | n17604 ;
  assign n17606 = ( ~x62 & n17599 ) | ( ~x62 & n17605 ) | ( n17599 & n17605 ) ;
  assign n17607 = x62 & ~n17605 ;
  assign n17608 = ( ~n17600 & n17606 ) | ( ~n17600 & n17607 ) | ( n17606 & n17607 ) ;
  assign n17609 = ( x62 & x63 ) | ( x62 & x107 ) | ( x63 & x107 ) ;
  assign n17610 = ( x62 & x106 ) | ( x62 & ~n9394 ) | ( x106 & ~n9394 ) ;
  assign n17611 = ( x106 & n17609 ) | ( x106 & ~n17610 ) | ( n17609 & ~n17610 ) ;
  assign n17612 = ( n17505 & n17608 ) | ( n17505 & ~n17611 ) | ( n17608 & ~n17611 ) ;
  assign n17613 = ( ~n17505 & n17608 ) | ( ~n17505 & n17611 ) | ( n17608 & n17611 ) ;
  assign n17614 = ( ~n17608 & n17612 ) | ( ~n17608 & n17613 ) | ( n17612 & n17613 ) ;
  assign n17615 = ( n17507 & n17598 ) | ( n17507 & ~n17614 ) | ( n17598 & ~n17614 ) ;
  assign n17616 = ( ~n17507 & n17598 ) | ( ~n17507 & n17614 ) | ( n17598 & n17614 ) ;
  assign n17617 = ( ~n17598 & n17615 ) | ( ~n17598 & n17616 ) | ( n17615 & n17616 ) ;
  assign n17618 = ( n17510 & n17588 ) | ( n17510 & ~n17617 ) | ( n17588 & ~n17617 ) ;
  assign n17619 = ( ~n17510 & n17588 ) | ( ~n17510 & n17617 ) | ( n17588 & n17617 ) ;
  assign n17620 = ( ~n17588 & n17618 ) | ( ~n17588 & n17619 ) | ( n17618 & n17619 ) ;
  assign n17621 = ( n17513 & n17578 ) | ( n17513 & ~n17620 ) | ( n17578 & ~n17620 ) ;
  assign n17622 = ( ~n17513 & n17578 ) | ( ~n17513 & n17620 ) | ( n17578 & n17620 ) ;
  assign n17623 = ( ~n17578 & n17621 ) | ( ~n17578 & n17622 ) | ( n17621 & n17622 ) ;
  assign n17624 = ( n17517 & n17568 ) | ( n17517 & ~n17623 ) | ( n17568 & ~n17623 ) ;
  assign n17625 = ( ~n17517 & n17568 ) | ( ~n17517 & n17623 ) | ( n17568 & n17623 ) ;
  assign n17626 = ( ~n17568 & n17624 ) | ( ~n17568 & n17625 ) | ( n17624 & n17625 ) ;
  assign n17627 = ( n17519 & n17558 ) | ( n17519 & ~n17626 ) | ( n17558 & ~n17626 ) ;
  assign n17628 = ( ~n17519 & n17558 ) | ( ~n17519 & n17626 ) | ( n17558 & n17626 ) ;
  assign n17629 = ( ~n17558 & n17627 ) | ( ~n17558 & n17628 ) | ( n17627 & n17628 ) ;
  assign n17630 = ( n17522 & n17548 ) | ( n17522 & ~n17629 ) | ( n17548 & ~n17629 ) ;
  assign n17631 = ( ~n17522 & n17548 ) | ( ~n17522 & n17629 ) | ( n17548 & n17629 ) ;
  assign n17632 = ( ~n17548 & n17630 ) | ( ~n17548 & n17631 ) | ( n17630 & n17631 ) ;
  assign n17633 = ( ~n17535 & n17538 ) | ( ~n17535 & n17632 ) | ( n17538 & n17632 ) ;
  assign n17634 = ( n17535 & n17538 ) | ( n17535 & ~n17632 ) | ( n17538 & ~n17632 ) ;
  assign n17635 = ( ~n17538 & n17633 ) | ( ~n17538 & n17634 ) | ( n17633 & n17634 ) ;
  assign n17636 = x43 & ~n4621 ;
  assign n17637 = ( x127 & n4794 ) | ( x127 & n9865 ) | ( n4794 & n9865 ) ;
  assign n17638 = ~n17636 & n17637 ;
  assign n17639 = ( n4621 & n17636 ) | ( n4621 & n17637 ) | ( n17636 & n17637 ) ;
  assign n17640 = ( x44 & ~n17638 ) | ( x44 & n17639 ) | ( ~n17638 & n17639 ) ;
  assign n17641 = n5223 & n9038 ;
  assign n17642 = x47 & n17641 ;
  assign n17643 = x126 & n5230 ;
  assign n17644 = x125 & n5227 ;
  assign n17645 = n17643 | n17644 ;
  assign n17646 = x124 & n5434 ;
  assign n17647 = n17645 | n17646 ;
  assign n17648 = ( ~x47 & n17641 ) | ( ~x47 & n17647 ) | ( n17641 & n17647 ) ;
  assign n17649 = x47 & ~n17647 ;
  assign n17650 = ( ~n17642 & n17648 ) | ( ~n17642 & n17649 ) | ( n17648 & n17649 ) ;
  assign n17651 = n5858 & n8461 ;
  assign n17652 = x50 & n17651 ;
  assign n17653 = x123 & n5865 ;
  assign n17654 = x122 & n5862 ;
  assign n17655 = n17653 | n17654 ;
  assign n17656 = x121 & n6092 ;
  assign n17657 = n17655 | n17656 ;
  assign n17658 = ( ~x50 & n17651 ) | ( ~x50 & n17657 ) | ( n17651 & n17657 ) ;
  assign n17659 = x50 & ~n17657 ;
  assign n17660 = ( ~n17652 & n17658 ) | ( ~n17652 & n17659 ) | ( n17658 & n17659 ) ;
  assign n17661 = n6546 & n7444 ;
  assign n17662 = x53 & n17661 ;
  assign n17663 = x120 & n6553 ;
  assign n17664 = x119 & n6550 ;
  assign n17665 = n17663 | n17664 ;
  assign n17666 = x118 & n6787 ;
  assign n17667 = n17665 | n17666 ;
  assign n17668 = ( ~x53 & n17661 ) | ( ~x53 & n17667 ) | ( n17661 & n17667 ) ;
  assign n17669 = x53 & ~n17667 ;
  assign n17670 = ( ~n17662 & n17668 ) | ( ~n17662 & n17669 ) | ( n17668 & n17669 ) ;
  assign n17671 = n6924 & n7277 ;
  assign n17672 = x56 & n17671 ;
  assign n17673 = x117 & n7545 ;
  assign n17674 = x116 & n7273 ;
  assign n17675 = n17673 | n17674 ;
  assign n17676 = x115 & n7552 ;
  assign n17677 = n17675 | n17676 ;
  assign n17678 = ( ~x56 & n17671 ) | ( ~x56 & n17677 ) | ( n17671 & n17677 ) ;
  assign n17679 = x56 & ~n17677 ;
  assign n17680 = ( ~n17672 & n17678 ) | ( ~n17672 & n17679 ) | ( n17678 & n17679 ) ;
  assign n17681 = n6002 & n8067 ;
  assign n17682 = x59 & n17681 ;
  assign n17683 = x114 & n8074 ;
  assign n17684 = x113 & n8071 ;
  assign n17685 = n17683 | n17684 ;
  assign n17686 = x112 & n8298 ;
  assign n17687 = n17685 | n17686 ;
  assign n17688 = ( ~x59 & n17681 ) | ( ~x59 & n17687 ) | ( n17681 & n17687 ) ;
  assign n17689 = x59 & ~n17687 ;
  assign n17690 = ( ~n17682 & n17688 ) | ( ~n17682 & n17689 ) | ( n17688 & n17689 ) ;
  assign n17691 = n5347 & n8859 ;
  assign n17692 = x62 & n17691 ;
  assign n17693 = x111 & n8866 ;
  assign n17694 = x110 & n8863 ;
  assign n17695 = n17693 | n17694 ;
  assign n17696 = x109 & n9125 ;
  assign n17697 = n17695 | n17696 ;
  assign n17698 = ( ~x62 & n17691 ) | ( ~x62 & n17697 ) | ( n17691 & n17697 ) ;
  assign n17699 = x62 & ~n17697 ;
  assign n17700 = ( ~n17692 & n17698 ) | ( ~n17692 & n17699 ) | ( n17698 & n17699 ) ;
  assign n17701 = ( x62 & x63 ) | ( x62 & x108 ) | ( x63 & x108 ) ;
  assign n17702 = ( x62 & x107 ) | ( x62 & ~n9394 ) | ( x107 & ~n9394 ) ;
  assign n17703 = ( x107 & n17701 ) | ( x107 & ~n17702 ) | ( n17701 & ~n17702 ) ;
  assign n17704 = ( ~n17611 & n17700 ) | ( ~n17611 & n17703 ) | ( n17700 & n17703 ) ;
  assign n17705 = ( n17611 & n17700 ) | ( n17611 & n17703 ) | ( n17700 & n17703 ) ;
  assign n17706 = ( n17611 & n17704 ) | ( n17611 & ~n17705 ) | ( n17704 & ~n17705 ) ;
  assign n17707 = ( ~n17612 & n17690 ) | ( ~n17612 & n17706 ) | ( n17690 & n17706 ) ;
  assign n17708 = ( n17612 & n17690 ) | ( n17612 & ~n17706 ) | ( n17690 & ~n17706 ) ;
  assign n17709 = ( ~n17690 & n17707 ) | ( ~n17690 & n17708 ) | ( n17707 & n17708 ) ;
  assign n17710 = ( n17615 & n17680 ) | ( n17615 & ~n17709 ) | ( n17680 & ~n17709 ) ;
  assign n17711 = ( ~n17615 & n17680 ) | ( ~n17615 & n17709 ) | ( n17680 & n17709 ) ;
  assign n17712 = ( ~n17680 & n17710 ) | ( ~n17680 & n17711 ) | ( n17710 & n17711 ) ;
  assign n17713 = ( n17618 & n17670 ) | ( n17618 & ~n17712 ) | ( n17670 & ~n17712 ) ;
  assign n17714 = ( ~n17618 & n17670 ) | ( ~n17618 & n17712 ) | ( n17670 & n17712 ) ;
  assign n17715 = ( ~n17670 & n17713 ) | ( ~n17670 & n17714 ) | ( n17713 & n17714 ) ;
  assign n17716 = ( n17621 & n17660 ) | ( n17621 & ~n17715 ) | ( n17660 & ~n17715 ) ;
  assign n17717 = ( ~n17621 & n17660 ) | ( ~n17621 & n17715 ) | ( n17660 & n17715 ) ;
  assign n17718 = ( ~n17660 & n17716 ) | ( ~n17660 & n17717 ) | ( n17716 & n17717 ) ;
  assign n17719 = ( ~n17624 & n17650 ) | ( ~n17624 & n17718 ) | ( n17650 & n17718 ) ;
  assign n17720 = ( n17624 & n17650 ) | ( n17624 & ~n17718 ) | ( n17650 & ~n17718 ) ;
  assign n17721 = ( ~n17650 & n17719 ) | ( ~n17650 & n17720 ) | ( n17719 & n17720 ) ;
  assign n17722 = ( ~n17627 & n17640 ) | ( ~n17627 & n17721 ) | ( n17640 & n17721 ) ;
  assign n17723 = ( n17627 & n17640 ) | ( n17627 & ~n17721 ) | ( n17640 & ~n17721 ) ;
  assign n17724 = ( ~n17640 & n17722 ) | ( ~n17640 & n17723 ) | ( n17722 & n17723 ) ;
  assign n17725 = ( ~n17630 & n17633 ) | ( ~n17630 & n17724 ) | ( n17633 & n17724 ) ;
  assign n17726 = ( n17630 & n17633 ) | ( n17630 & ~n17724 ) | ( n17633 & ~n17724 ) ;
  assign n17727 = ( ~n17633 & n17725 ) | ( ~n17633 & n17726 ) | ( n17725 & n17726 ) ;
  assign n17728 = n5858 & n8729 ;
  assign n17729 = x50 & n17728 ;
  assign n17730 = x124 & n5865 ;
  assign n17731 = x123 & n5862 ;
  assign n17732 = n17730 | n17731 ;
  assign n17733 = x122 & n6092 ;
  assign n17734 = n17732 | n17733 ;
  assign n17735 = ( ~x50 & n17728 ) | ( ~x50 & n17734 ) | ( n17728 & n17734 ) ;
  assign n17736 = x50 & ~n17734 ;
  assign n17737 = ( ~n17729 & n17735 ) | ( ~n17729 & n17736 ) | ( n17735 & n17736 ) ;
  assign n17738 = n6546 & n7696 ;
  assign n17739 = x53 & n17738 ;
  assign n17740 = x121 & n6553 ;
  assign n17741 = x120 & n6550 ;
  assign n17742 = n17740 | n17741 ;
  assign n17743 = x119 & n6787 ;
  assign n17744 = n17742 | n17743 ;
  assign n17745 = ( ~x53 & n17738 ) | ( ~x53 & n17744 ) | ( n17738 & n17744 ) ;
  assign n17746 = x53 & ~n17744 ;
  assign n17747 = ( ~n17739 & n17745 ) | ( ~n17739 & n17746 ) | ( n17745 & n17746 ) ;
  assign n17748 = n6940 & n7277 ;
  assign n17749 = x56 & n17748 ;
  assign n17750 = x118 & n7545 ;
  assign n17751 = x117 & n7273 ;
  assign n17752 = n17750 | n17751 ;
  assign n17753 = x116 & n7552 ;
  assign n17754 = n17752 | n17753 ;
  assign n17755 = ( ~x56 & n17748 ) | ( ~x56 & n17754 ) | ( n17748 & n17754 ) ;
  assign n17756 = x56 & ~n17754 ;
  assign n17757 = ( ~n17749 & n17755 ) | ( ~n17749 & n17756 ) | ( n17755 & n17756 ) ;
  assign n17758 = n6446 & n8067 ;
  assign n17759 = x59 & n17758 ;
  assign n17760 = x115 & n8074 ;
  assign n17761 = x114 & n8071 ;
  assign n17762 = n17760 | n17761 ;
  assign n17763 = x113 & n8298 ;
  assign n17764 = n17762 | n17763 ;
  assign n17765 = ( ~x59 & n17758 ) | ( ~x59 & n17764 ) | ( n17758 & n17764 ) ;
  assign n17766 = x59 & ~n17764 ;
  assign n17767 = ( ~n17759 & n17765 ) | ( ~n17759 & n17766 ) | ( n17765 & n17766 ) ;
  assign n17768 = n5558 & n8859 ;
  assign n17769 = x62 & n17768 ;
  assign n17770 = x112 & n8866 ;
  assign n17771 = x111 & n8863 ;
  assign n17772 = n17770 | n17771 ;
  assign n17773 = x110 & n9125 ;
  assign n17774 = n17772 | n17773 ;
  assign n17775 = ( ~x62 & n17768 ) | ( ~x62 & n17774 ) | ( n17768 & n17774 ) ;
  assign n17776 = x62 & ~n17774 ;
  assign n17777 = ( ~n17769 & n17775 ) | ( ~n17769 & n17776 ) | ( n17775 & n17776 ) ;
  assign n17778 = ( x62 & x63 ) | ( x62 & x109 ) | ( x63 & x109 ) ;
  assign n17779 = ( x62 & x108 ) | ( x62 & ~n9394 ) | ( x108 & ~n9394 ) ;
  assign n17780 = ( x108 & n17778 ) | ( x108 & ~n17779 ) | ( n17778 & ~n17779 ) ;
  assign n17781 = ( x44 & n17611 ) | ( x44 & n17780 ) | ( n17611 & n17780 ) ;
  assign n17782 = ( ~x44 & n17611 ) | ( ~x44 & n17780 ) | ( n17611 & n17780 ) ;
  assign n17783 = ( x44 & ~n17781 ) | ( x44 & n17782 ) | ( ~n17781 & n17782 ) ;
  assign n17784 = ( n17704 & n17777 ) | ( n17704 & ~n17783 ) | ( n17777 & ~n17783 ) ;
  assign n17785 = ( n17704 & ~n17777 ) | ( n17704 & n17783 ) | ( ~n17777 & n17783 ) ;
  assign n17786 = ( ~n17704 & n17784 ) | ( ~n17704 & n17785 ) | ( n17784 & n17785 ) ;
  assign n17787 = ( n17708 & n17767 ) | ( n17708 & ~n17786 ) | ( n17767 & ~n17786 ) ;
  assign n17788 = ( n17708 & ~n17767 ) | ( n17708 & n17786 ) | ( ~n17767 & n17786 ) ;
  assign n17789 = ( ~n17708 & n17787 ) | ( ~n17708 & n17788 ) | ( n17787 & n17788 ) ;
  assign n17790 = ( n17710 & n17757 ) | ( n17710 & ~n17789 ) | ( n17757 & ~n17789 ) ;
  assign n17791 = ( n17710 & ~n17757 ) | ( n17710 & n17789 ) | ( ~n17757 & n17789 ) ;
  assign n17792 = ( ~n17710 & n17790 ) | ( ~n17710 & n17791 ) | ( n17790 & n17791 ) ;
  assign n17793 = ( n17713 & n17747 ) | ( n17713 & ~n17792 ) | ( n17747 & ~n17792 ) ;
  assign n17794 = ( n17713 & ~n17747 ) | ( n17713 & n17792 ) | ( ~n17747 & n17792 ) ;
  assign n17795 = ( ~n17713 & n17793 ) | ( ~n17713 & n17794 ) | ( n17793 & n17794 ) ;
  assign n17796 = ( n17716 & ~n17737 ) | ( n17716 & n17795 ) | ( ~n17737 & n17795 ) ;
  assign n17797 = ( n17716 & n17737 ) | ( n17716 & ~n17795 ) | ( n17737 & ~n17795 ) ;
  assign n17798 = ( ~n17716 & n17796 ) | ( ~n17716 & n17797 ) | ( n17796 & n17797 ) ;
  assign n17799 = n5223 & n9576 ;
  assign n17800 = x47 & n17799 ;
  assign n17801 = x127 & n5230 ;
  assign n17802 = x126 & n5227 ;
  assign n17803 = n17801 | n17802 ;
  assign n17804 = x125 & n5434 ;
  assign n17805 = n17803 | n17804 ;
  assign n17806 = ( ~x47 & n17799 ) | ( ~x47 & n17805 ) | ( n17799 & n17805 ) ;
  assign n17807 = x47 & ~n17805 ;
  assign n17808 = ( ~n17800 & n17806 ) | ( ~n17800 & n17807 ) | ( n17806 & n17807 ) ;
  assign n17809 = ( n17720 & ~n17798 ) | ( n17720 & n17808 ) | ( ~n17798 & n17808 ) ;
  assign n17810 = ( n17720 & n17798 ) | ( n17720 & ~n17808 ) | ( n17798 & ~n17808 ) ;
  assign n17811 = ( ~n17720 & n17809 ) | ( ~n17720 & n17810 ) | ( n17809 & n17810 ) ;
  assign n17812 = ( n17723 & n17725 ) | ( n17723 & ~n17811 ) | ( n17725 & ~n17811 ) ;
  assign n17813 = ( ~n17723 & n17725 ) | ( ~n17723 & n17811 ) | ( n17725 & n17811 ) ;
  assign n17814 = ( ~n17725 & n17812 ) | ( ~n17725 & n17813 ) | ( n17812 & n17813 ) ;
  assign n17815 = x127 & n5227 ;
  assign n17816 = n5223 | n17815 ;
  assign n17817 = ( n9867 & n17815 ) | ( n9867 & n17816 ) | ( n17815 & n17816 ) ;
  assign n17818 = x126 & n5434 ;
  assign n17819 = ( ~x47 & n17817 ) | ( ~x47 & n17818 ) | ( n17817 & n17818 ) ;
  assign n17820 = ( x47 & ~n17817 ) | ( x47 & n17818 ) | ( ~n17817 & n17818 ) ;
  assign n17821 = ~n17818 & n17820 ;
  assign n17822 = n17819 | n17821 ;
  assign n17823 = n5858 & n9009 ;
  assign n17824 = x50 & n17823 ;
  assign n17825 = x125 & n5865 ;
  assign n17826 = x124 & n5862 ;
  assign n17827 = n17825 | n17826 ;
  assign n17828 = x123 & n6092 ;
  assign n17829 = n17827 | n17828 ;
  assign n17830 = ( ~x50 & n17823 ) | ( ~x50 & n17829 ) | ( n17823 & n17829 ) ;
  assign n17831 = x50 & ~n17829 ;
  assign n17832 = ( ~n17824 & n17830 ) | ( ~n17824 & n17831 ) | ( n17830 & n17831 ) ;
  assign n17833 = n6546 & n8207 ;
  assign n17834 = x53 & n17833 ;
  assign n17835 = x122 & n6553 ;
  assign n17836 = x121 & n6550 ;
  assign n17837 = n17835 | n17836 ;
  assign n17838 = x120 & n6787 ;
  assign n17839 = n17837 | n17838 ;
  assign n17840 = ( ~x53 & n17833 ) | ( ~x53 & n17839 ) | ( n17833 & n17839 ) ;
  assign n17841 = x53 & ~n17839 ;
  assign n17842 = ( ~n17834 & n17840 ) | ( ~n17834 & n17841 ) | ( n17840 & n17841 ) ;
  assign n17843 = n7181 & n7277 ;
  assign n17844 = x56 & n17843 ;
  assign n17845 = x119 & n7545 ;
  assign n17846 = x118 & n7273 ;
  assign n17847 = n17845 | n17846 ;
  assign n17848 = x117 & n7552 ;
  assign n17849 = n17847 | n17848 ;
  assign n17850 = ( ~x56 & n17843 ) | ( ~x56 & n17849 ) | ( n17843 & n17849 ) ;
  assign n17851 = x56 & ~n17849 ;
  assign n17852 = ( ~n17844 & n17850 ) | ( ~n17844 & n17851 ) | ( n17850 & n17851 ) ;
  assign n17853 = n6462 & n8067 ;
  assign n17854 = x59 & n17853 ;
  assign n17855 = x116 & n8074 ;
  assign n17856 = x115 & n8071 ;
  assign n17857 = n17855 | n17856 ;
  assign n17858 = x114 & n8298 ;
  assign n17859 = n17857 | n17858 ;
  assign n17860 = ( ~x59 & n17853 ) | ( ~x59 & n17859 ) | ( n17853 & n17859 ) ;
  assign n17861 = x59 & ~n17859 ;
  assign n17862 = ( ~n17854 & n17860 ) | ( ~n17854 & n17861 ) | ( n17860 & n17861 ) ;
  assign n17863 = ( x62 & x63 ) | ( x62 & x110 ) | ( x63 & x110 ) ;
  assign n17864 = ( x62 & x109 ) | ( x62 & ~n9394 ) | ( x109 & ~n9394 ) ;
  assign n17865 = ( x109 & n17863 ) | ( x109 & ~n17864 ) | ( n17863 & ~n17864 ) ;
  assign n17866 = n5774 & n8859 ;
  assign n17867 = x62 & n17866 ;
  assign n17868 = x113 & n8866 ;
  assign n17869 = x112 & n8863 ;
  assign n17870 = n17868 | n17869 ;
  assign n17871 = x111 & n9125 ;
  assign n17872 = n17870 | n17871 ;
  assign n17873 = ( ~x62 & n17866 ) | ( ~x62 & n17872 ) | ( n17866 & n17872 ) ;
  assign n17874 = x62 & ~n17872 ;
  assign n17875 = ( ~n17867 & n17873 ) | ( ~n17867 & n17874 ) | ( n17873 & n17874 ) ;
  assign n17876 = ( ~n17782 & n17865 ) | ( ~n17782 & n17875 ) | ( n17865 & n17875 ) ;
  assign n17877 = ( n17782 & n17865 ) | ( n17782 & ~n17875 ) | ( n17865 & ~n17875 ) ;
  assign n17878 = ( ~n17865 & n17876 ) | ( ~n17865 & n17877 ) | ( n17876 & n17877 ) ;
  assign n17879 = ( ~n17784 & n17862 ) | ( ~n17784 & n17878 ) | ( n17862 & n17878 ) ;
  assign n17880 = ( n17784 & n17862 ) | ( n17784 & ~n17878 ) | ( n17862 & ~n17878 ) ;
  assign n17881 = ( ~n17862 & n17879 ) | ( ~n17862 & n17880 ) | ( n17879 & n17880 ) ;
  assign n17882 = ( n17787 & n17852 ) | ( n17787 & ~n17881 ) | ( n17852 & ~n17881 ) ;
  assign n17883 = ( ~n17787 & n17852 ) | ( ~n17787 & n17881 ) | ( n17852 & n17881 ) ;
  assign n17884 = ( ~n17852 & n17882 ) | ( ~n17852 & n17883 ) | ( n17882 & n17883 ) ;
  assign n17885 = ( n17790 & n17842 ) | ( n17790 & ~n17884 ) | ( n17842 & ~n17884 ) ;
  assign n17886 = ( ~n17790 & n17842 ) | ( ~n17790 & n17884 ) | ( n17842 & n17884 ) ;
  assign n17887 = ( ~n17842 & n17885 ) | ( ~n17842 & n17886 ) | ( n17885 & n17886 ) ;
  assign n17888 = ( ~n17793 & n17832 ) | ( ~n17793 & n17887 ) | ( n17832 & n17887 ) ;
  assign n17889 = ( n17793 & n17832 ) | ( n17793 & ~n17887 ) | ( n17832 & ~n17887 ) ;
  assign n17890 = ( ~n17832 & n17888 ) | ( ~n17832 & n17889 ) | ( n17888 & n17889 ) ;
  assign n17891 = ( n17797 & n17822 ) | ( n17797 & ~n17890 ) | ( n17822 & ~n17890 ) ;
  assign n17892 = ( ~n17797 & n17822 ) | ( ~n17797 & n17890 ) | ( n17822 & n17890 ) ;
  assign n17893 = ( ~n17822 & n17891 ) | ( ~n17822 & n17892 ) | ( n17891 & n17892 ) ;
  assign n17894 = ( n17809 & n17813 ) | ( n17809 & ~n17893 ) | ( n17813 & ~n17893 ) ;
  assign n17895 = ( ~n17809 & n17813 ) | ( ~n17809 & n17893 ) | ( n17813 & n17893 ) ;
  assign n17896 = ( ~n17813 & n17894 ) | ( ~n17813 & n17895 ) | ( n17894 & n17895 ) ;
  assign n17897 = n5858 & n9038 ;
  assign n17898 = x50 & n17897 ;
  assign n17899 = x126 & n5865 ;
  assign n17900 = x125 & n5862 ;
  assign n17901 = n17899 | n17900 ;
  assign n17902 = x124 & n6092 ;
  assign n17903 = n17901 | n17902 ;
  assign n17904 = ( ~x50 & n17897 ) | ( ~x50 & n17903 ) | ( n17897 & n17903 ) ;
  assign n17905 = x50 & ~n17903 ;
  assign n17906 = ( ~n17898 & n17904 ) | ( ~n17898 & n17905 ) | ( n17904 & n17905 ) ;
  assign n17907 = n6546 & n8461 ;
  assign n17908 = x53 & n17907 ;
  assign n17909 = x123 & n6553 ;
  assign n17910 = x122 & n6550 ;
  assign n17911 = n17909 | n17910 ;
  assign n17912 = x121 & n6787 ;
  assign n17913 = n17911 | n17912 ;
  assign n17914 = ( ~x53 & n17907 ) | ( ~x53 & n17913 ) | ( n17907 & n17913 ) ;
  assign n17915 = x53 & ~n17913 ;
  assign n17916 = ( ~n17908 & n17914 ) | ( ~n17908 & n17915 ) | ( n17914 & n17915 ) ;
  assign n17917 = n7277 & n7444 ;
  assign n17918 = x56 & n17917 ;
  assign n17919 = x120 & n7545 ;
  assign n17920 = x119 & n7273 ;
  assign n17921 = n17919 | n17920 ;
  assign n17922 = x118 & n7552 ;
  assign n17923 = n17921 | n17922 ;
  assign n17924 = ( ~x56 & n17917 ) | ( ~x56 & n17923 ) | ( n17917 & n17923 ) ;
  assign n17925 = x56 & ~n17923 ;
  assign n17926 = ( ~n17918 & n17924 ) | ( ~n17918 & n17925 ) | ( n17924 & n17925 ) ;
  assign n17927 = n6924 & n8067 ;
  assign n17928 = x59 & n17927 ;
  assign n17929 = x117 & n8074 ;
  assign n17930 = x116 & n8071 ;
  assign n17931 = n17929 | n17930 ;
  assign n17932 = x115 & n8298 ;
  assign n17933 = n17931 | n17932 ;
  assign n17934 = ( ~x59 & n17927 ) | ( ~x59 & n17933 ) | ( n17927 & n17933 ) ;
  assign n17935 = x59 & ~n17933 ;
  assign n17936 = ( ~n17928 & n17934 ) | ( ~n17928 & n17935 ) | ( n17934 & n17935 ) ;
  assign n17937 = n6002 & n8859 ;
  assign n17938 = x62 & n17937 ;
  assign n17939 = x114 & n8866 ;
  assign n17940 = x113 & n8863 ;
  assign n17941 = n17939 | n17940 ;
  assign n17942 = x112 & n9125 ;
  assign n17943 = n17941 | n17942 ;
  assign n17944 = ( ~x62 & n17937 ) | ( ~x62 & n17943 ) | ( n17937 & n17943 ) ;
  assign n17945 = x62 & ~n17943 ;
  assign n17946 = ( ~n17938 & n17944 ) | ( ~n17938 & n17945 ) | ( n17944 & n17945 ) ;
  assign n17947 = ( x62 & x63 ) | ( x62 & x111 ) | ( x63 & x111 ) ;
  assign n17948 = ( x62 & x110 ) | ( x62 & ~n9394 ) | ( x110 & ~n9394 ) ;
  assign n17949 = ( x110 & n17947 ) | ( x110 & ~n17948 ) | ( n17947 & ~n17948 ) ;
  assign n17950 = ( n17875 & ~n17877 ) | ( n17875 & n17949 ) | ( ~n17877 & n17949 ) ;
  assign n17951 = ( n17782 & n17876 ) | ( n17782 & ~n17949 ) | ( n17876 & ~n17949 ) ;
  assign n17952 = ( ~n17875 & n17950 ) | ( ~n17875 & n17951 ) | ( n17950 & n17951 ) ;
  assign n17953 = ( n17936 & n17946 ) | ( n17936 & ~n17952 ) | ( n17946 & ~n17952 ) ;
  assign n17954 = ( n17936 & ~n17946 ) | ( n17936 & n17952 ) | ( ~n17946 & n17952 ) ;
  assign n17955 = ( ~n17936 & n17953 ) | ( ~n17936 & n17954 ) | ( n17953 & n17954 ) ;
  assign n17956 = ( n17880 & n17926 ) | ( n17880 & ~n17955 ) | ( n17926 & ~n17955 ) ;
  assign n17957 = ( ~n17880 & n17926 ) | ( ~n17880 & n17955 ) | ( n17926 & n17955 ) ;
  assign n17958 = ( ~n17926 & n17956 ) | ( ~n17926 & n17957 ) | ( n17956 & n17957 ) ;
  assign n17959 = ( n17882 & n17916 ) | ( n17882 & ~n17958 ) | ( n17916 & ~n17958 ) ;
  assign n17960 = ( ~n17882 & n17916 ) | ( ~n17882 & n17958 ) | ( n17916 & n17958 ) ;
  assign n17961 = ( ~n17916 & n17959 ) | ( ~n17916 & n17960 ) | ( n17959 & n17960 ) ;
  assign n17962 = ( ~n17885 & n17906 ) | ( ~n17885 & n17961 ) | ( n17906 & n17961 ) ;
  assign n17963 = ( n17885 & n17906 ) | ( n17885 & ~n17961 ) | ( n17906 & ~n17961 ) ;
  assign n17964 = ( ~n17906 & n17962 ) | ( ~n17906 & n17963 ) | ( n17962 & n17963 ) ;
  assign n17965 = n5433 | n9864 ;
  assign n17966 = x127 & ~n5227 ;
  assign n17967 = n17965 & n17966 ;
  assign n17968 = x47 | n17967 ;
  assign n17969 = ~x46 & n17967 ;
  assign n17970 = n17968 & ~n17969 ;
  assign n17971 = ( n17889 & ~n17964 ) | ( n17889 & n17970 ) | ( ~n17964 & n17970 ) ;
  assign n17972 = ( n17889 & n17964 ) | ( n17889 & n17970 ) | ( n17964 & n17970 ) ;
  assign n17973 = ( n17964 & n17971 ) | ( n17964 & ~n17972 ) | ( n17971 & ~n17972 ) ;
  assign n17974 = ( ~n17891 & n17895 ) | ( ~n17891 & n17973 ) | ( n17895 & n17973 ) ;
  assign n17975 = ( n17891 & n17895 ) | ( n17891 & ~n17973 ) | ( n17895 & ~n17973 ) ;
  assign n17976 = ( ~n17895 & n17974 ) | ( ~n17895 & n17975 ) | ( n17974 & n17975 ) ;
  assign n17977 = n5858 & n9576 ;
  assign n17978 = x50 & n17977 ;
  assign n17979 = x127 & n5865 ;
  assign n17980 = x126 & n5862 ;
  assign n17981 = n17979 | n17980 ;
  assign n17982 = x125 & n6092 ;
  assign n17983 = n17981 | n17982 ;
  assign n17984 = ( ~x50 & n17977 ) | ( ~x50 & n17983 ) | ( n17977 & n17983 ) ;
  assign n17985 = x50 & ~n17983 ;
  assign n17986 = ( ~n17978 & n17984 ) | ( ~n17978 & n17985 ) | ( n17984 & n17985 ) ;
  assign n17987 = n6546 & n8729 ;
  assign n17988 = x53 & n17987 ;
  assign n17989 = x124 & n6553 ;
  assign n17990 = x123 & n6550 ;
  assign n17991 = n17989 | n17990 ;
  assign n17992 = x122 & n6787 ;
  assign n17993 = n17991 | n17992 ;
  assign n17994 = ( ~x53 & n17987 ) | ( ~x53 & n17993 ) | ( n17987 & n17993 ) ;
  assign n17995 = x53 & ~n17993 ;
  assign n17996 = ( ~n17988 & n17994 ) | ( ~n17988 & n17995 ) | ( n17994 & n17995 ) ;
  assign n17997 = n7277 & n7696 ;
  assign n17998 = x56 & n17997 ;
  assign n17999 = x121 & n7545 ;
  assign n18000 = x120 & n7273 ;
  assign n18001 = n17999 | n18000 ;
  assign n18002 = x119 & n7552 ;
  assign n18003 = n18001 | n18002 ;
  assign n18004 = ( ~x56 & n17997 ) | ( ~x56 & n18003 ) | ( n17997 & n18003 ) ;
  assign n18005 = x56 & ~n18003 ;
  assign n18006 = ( ~n17998 & n18004 ) | ( ~n17998 & n18005 ) | ( n18004 & n18005 ) ;
  assign n18007 = n6940 & n8067 ;
  assign n18008 = x59 & n18007 ;
  assign n18009 = x118 & n8074 ;
  assign n18010 = x117 & n8071 ;
  assign n18011 = n18009 | n18010 ;
  assign n18012 = x116 & n8298 ;
  assign n18013 = n18011 | n18012 ;
  assign n18014 = ( ~x59 & n18007 ) | ( ~x59 & n18013 ) | ( n18007 & n18013 ) ;
  assign n18015 = x59 & ~n18013 ;
  assign n18016 = ( ~n18008 & n18014 ) | ( ~n18008 & n18015 ) | ( n18014 & n18015 ) ;
  assign n18017 = n6446 & n8859 ;
  assign n18018 = x62 & n18017 ;
  assign n18019 = x115 & n8866 ;
  assign n18020 = x114 & n8863 ;
  assign n18021 = n18019 | n18020 ;
  assign n18022 = x113 & n9125 ;
  assign n18023 = n18021 | n18022 ;
  assign n18024 = ( ~x62 & n18017 ) | ( ~x62 & n18023 ) | ( n18017 & n18023 ) ;
  assign n18025 = x62 & ~n18023 ;
  assign n18026 = ( ~n18018 & n18024 ) | ( ~n18018 & n18025 ) | ( n18024 & n18025 ) ;
  assign n18027 = ( x62 & x63 ) | ( x62 & x112 ) | ( x63 & x112 ) ;
  assign n18028 = ( x62 & x111 ) | ( x62 & ~n9394 ) | ( x111 & ~n9394 ) ;
  assign n18029 = ( x111 & n18027 ) | ( x111 & ~n18028 ) | ( n18027 & ~n18028 ) ;
  assign n18030 = ( x47 & n17949 ) | ( x47 & n18029 ) | ( n17949 & n18029 ) ;
  assign n18031 = ( ~x47 & n17949 ) | ( ~x47 & n18029 ) | ( n17949 & n18029 ) ;
  assign n18032 = ( x47 & ~n18030 ) | ( x47 & n18031 ) | ( ~n18030 & n18031 ) ;
  assign n18033 = ( n17951 & n18026 ) | ( n17951 & ~n18032 ) | ( n18026 & ~n18032 ) ;
  assign n18034 = ( ~n17951 & n18026 ) | ( ~n17951 & n18032 ) | ( n18026 & n18032 ) ;
  assign n18035 = ( ~n18026 & n18033 ) | ( ~n18026 & n18034 ) | ( n18033 & n18034 ) ;
  assign n18036 = ( n17953 & n18016 ) | ( n17953 & ~n18035 ) | ( n18016 & ~n18035 ) ;
  assign n18037 = ( n17953 & ~n18016 ) | ( n17953 & n18035 ) | ( ~n18016 & n18035 ) ;
  assign n18038 = ( ~n17953 & n18036 ) | ( ~n17953 & n18037 ) | ( n18036 & n18037 ) ;
  assign n18039 = ( n17956 & n18006 ) | ( n17956 & ~n18038 ) | ( n18006 & ~n18038 ) ;
  assign n18040 = ( n17956 & ~n18006 ) | ( n17956 & n18038 ) | ( ~n18006 & n18038 ) ;
  assign n18041 = ( ~n17956 & n18039 ) | ( ~n17956 & n18040 ) | ( n18039 & n18040 ) ;
  assign n18042 = ( n17959 & n17996 ) | ( n17959 & ~n18041 ) | ( n17996 & ~n18041 ) ;
  assign n18043 = ( n17959 & ~n17996 ) | ( n17959 & n18041 ) | ( ~n17996 & n18041 ) ;
  assign n18044 = ( ~n17959 & n18042 ) | ( ~n17959 & n18043 ) | ( n18042 & n18043 ) ;
  assign n18045 = ( n17963 & n17986 ) | ( n17963 & ~n18044 ) | ( n17986 & ~n18044 ) ;
  assign n18046 = ( n17963 & ~n17986 ) | ( n17963 & n18044 ) | ( ~n17986 & n18044 ) ;
  assign n18047 = ( ~n17963 & n18045 ) | ( ~n17963 & n18046 ) | ( n18045 & n18046 ) ;
  assign n18048 = ( n17971 & n17974 ) | ( n17971 & ~n18047 ) | ( n17974 & ~n18047 ) ;
  assign n18049 = ( ~n17971 & n17974 ) | ( ~n17971 & n18047 ) | ( n17974 & n18047 ) ;
  assign n18050 = ( ~n17974 & n18048 ) | ( ~n17974 & n18049 ) | ( n18048 & n18049 ) ;
  assign n18051 = x127 & n5862 ;
  assign n18052 = n5858 | n18051 ;
  assign n18053 = ( n9867 & n18051 ) | ( n9867 & n18052 ) | ( n18051 & n18052 ) ;
  assign n18054 = x126 & n6092 ;
  assign n18055 = ( ~x50 & n18053 ) | ( ~x50 & n18054 ) | ( n18053 & n18054 ) ;
  assign n18056 = ( x50 & ~n18053 ) | ( x50 & n18054 ) | ( ~n18053 & n18054 ) ;
  assign n18057 = ~n18054 & n18056 ;
  assign n18058 = n18055 | n18057 ;
  assign n18059 = n6546 & n9009 ;
  assign n18060 = x53 & n18059 ;
  assign n18061 = x125 & n6553 ;
  assign n18062 = x124 & n6550 ;
  assign n18063 = n18061 | n18062 ;
  assign n18064 = x123 & n6787 ;
  assign n18065 = n18063 | n18064 ;
  assign n18066 = ( ~x53 & n18059 ) | ( ~x53 & n18065 ) | ( n18059 & n18065 ) ;
  assign n18067 = x53 & ~n18065 ;
  assign n18068 = ( ~n18060 & n18066 ) | ( ~n18060 & n18067 ) | ( n18066 & n18067 ) ;
  assign n18069 = n7277 & n8207 ;
  assign n18070 = x56 & n18069 ;
  assign n18071 = x122 & n7545 ;
  assign n18072 = x121 & n7273 ;
  assign n18073 = n18071 | n18072 ;
  assign n18074 = x120 & n7552 ;
  assign n18075 = n18073 | n18074 ;
  assign n18076 = ( ~x56 & n18069 ) | ( ~x56 & n18075 ) | ( n18069 & n18075 ) ;
  assign n18077 = x56 & ~n18075 ;
  assign n18078 = ( ~n18070 & n18076 ) | ( ~n18070 & n18077 ) | ( n18076 & n18077 ) ;
  assign n18079 = n7181 & n8067 ;
  assign n18080 = x59 & n18079 ;
  assign n18081 = x119 & n8074 ;
  assign n18082 = x118 & n8071 ;
  assign n18083 = n18081 | n18082 ;
  assign n18084 = x117 & n8298 ;
  assign n18085 = n18083 | n18084 ;
  assign n18086 = ( ~x59 & n18079 ) | ( ~x59 & n18085 ) | ( n18079 & n18085 ) ;
  assign n18087 = x59 & ~n18085 ;
  assign n18088 = ( ~n18080 & n18086 ) | ( ~n18080 & n18087 ) | ( n18086 & n18087 ) ;
  assign n18089 = n6462 & n8859 ;
  assign n18090 = x62 & n18089 ;
  assign n18091 = x116 & n8866 ;
  assign n18092 = x115 & n8863 ;
  assign n18093 = n18091 | n18092 ;
  assign n18094 = x114 & n9125 ;
  assign n18095 = n18093 | n18094 ;
  assign n18096 = ( ~x62 & n18089 ) | ( ~x62 & n18095 ) | ( n18089 & n18095 ) ;
  assign n18097 = x62 & ~n18095 ;
  assign n18098 = ( ~n18090 & n18096 ) | ( ~n18090 & n18097 ) | ( n18096 & n18097 ) ;
  assign n18099 = ( x62 & x63 ) | ( x62 & x113 ) | ( x63 & x113 ) ;
  assign n18100 = ( x62 & x112 ) | ( x62 & ~n9394 ) | ( x112 & ~n9394 ) ;
  assign n18101 = ( x112 & n18099 ) | ( x112 & ~n18100 ) | ( n18099 & ~n18100 ) ;
  assign n18102 = ( n18031 & n18098 ) | ( n18031 & ~n18101 ) | ( n18098 & ~n18101 ) ;
  assign n18103 = ( ~n18031 & n18098 ) | ( ~n18031 & n18101 ) | ( n18098 & n18101 ) ;
  assign n18104 = ( ~n18098 & n18102 ) | ( ~n18098 & n18103 ) | ( n18102 & n18103 ) ;
  assign n18105 = ( n18033 & n18088 ) | ( n18033 & ~n18104 ) | ( n18088 & ~n18104 ) ;
  assign n18106 = ( ~n18033 & n18088 ) | ( ~n18033 & n18104 ) | ( n18088 & n18104 ) ;
  assign n18107 = ( ~n18088 & n18105 ) | ( ~n18088 & n18106 ) | ( n18105 & n18106 ) ;
  assign n18108 = ( n18036 & n18078 ) | ( n18036 & ~n18107 ) | ( n18078 & ~n18107 ) ;
  assign n18109 = ( ~n18036 & n18078 ) | ( ~n18036 & n18107 ) | ( n18078 & n18107 ) ;
  assign n18110 = ( ~n18078 & n18108 ) | ( ~n18078 & n18109 ) | ( n18108 & n18109 ) ;
  assign n18111 = ( n18039 & n18068 ) | ( n18039 & ~n18110 ) | ( n18068 & ~n18110 ) ;
  assign n18112 = ( ~n18039 & n18068 ) | ( ~n18039 & n18110 ) | ( n18068 & n18110 ) ;
  assign n18113 = ( ~n18068 & n18111 ) | ( ~n18068 & n18112 ) | ( n18111 & n18112 ) ;
  assign n18114 = ( ~n18042 & n18058 ) | ( ~n18042 & n18113 ) | ( n18058 & n18113 ) ;
  assign n18115 = ( n18042 & n18058 ) | ( n18042 & ~n18113 ) | ( n18058 & ~n18113 ) ;
  assign n18116 = ( ~n18058 & n18114 ) | ( ~n18058 & n18115 ) | ( n18114 & n18115 ) ;
  assign n18117 = ( ~n18045 & n18049 ) | ( ~n18045 & n18116 ) | ( n18049 & n18116 ) ;
  assign n18118 = ( n18045 & n18049 ) | ( n18045 & ~n18116 ) | ( n18049 & ~n18116 ) ;
  assign n18119 = ( ~n18049 & n18117 ) | ( ~n18049 & n18118 ) | ( n18117 & n18118 ) ;
  assign n18120 = n6546 & n9038 ;
  assign n18121 = x53 & n18120 ;
  assign n18122 = x126 & n6553 ;
  assign n18123 = x125 & n6550 ;
  assign n18124 = n18122 | n18123 ;
  assign n18125 = x124 & n6787 ;
  assign n18126 = n18124 | n18125 ;
  assign n18127 = ( ~x53 & n18120 ) | ( ~x53 & n18126 ) | ( n18120 & n18126 ) ;
  assign n18128 = x53 & ~n18126 ;
  assign n18129 = ( ~n18121 & n18127 ) | ( ~n18121 & n18128 ) | ( n18127 & n18128 ) ;
  assign n18130 = n7277 & n8461 ;
  assign n18131 = x56 & n18130 ;
  assign n18132 = x123 & n7545 ;
  assign n18133 = x122 & n7273 ;
  assign n18134 = n18132 | n18133 ;
  assign n18135 = x121 & n7552 ;
  assign n18136 = n18134 | n18135 ;
  assign n18137 = ( ~x56 & n18130 ) | ( ~x56 & n18136 ) | ( n18130 & n18136 ) ;
  assign n18138 = x56 & ~n18136 ;
  assign n18139 = ( ~n18131 & n18137 ) | ( ~n18131 & n18138 ) | ( n18137 & n18138 ) ;
  assign n18140 = n7444 & n8067 ;
  assign n18141 = x59 & n18140 ;
  assign n18142 = x120 & n8074 ;
  assign n18143 = x119 & n8071 ;
  assign n18144 = n18142 | n18143 ;
  assign n18145 = x118 & n8298 ;
  assign n18146 = n18144 | n18145 ;
  assign n18147 = ( ~x59 & n18140 ) | ( ~x59 & n18146 ) | ( n18140 & n18146 ) ;
  assign n18148 = x59 & ~n18146 ;
  assign n18149 = ( ~n18141 & n18147 ) | ( ~n18141 & n18148 ) | ( n18147 & n18148 ) ;
  assign n18150 = n6924 & n8859 ;
  assign n18151 = x62 & n18150 ;
  assign n18152 = x117 & n8866 ;
  assign n18153 = x116 & n8863 ;
  assign n18154 = n18152 | n18153 ;
  assign n18155 = x115 & n9125 ;
  assign n18156 = n18154 | n18155 ;
  assign n18157 = ( ~x62 & n18150 ) | ( ~x62 & n18156 ) | ( n18150 & n18156 ) ;
  assign n18158 = x62 & ~n18156 ;
  assign n18159 = ( ~n18151 & n18157 ) | ( ~n18151 & n18158 ) | ( n18157 & n18158 ) ;
  assign n18160 = ( x62 & x63 ) | ( x62 & x114 ) | ( x63 & x114 ) ;
  assign n18161 = ( x62 & x113 ) | ( x62 & ~n9394 ) | ( x113 & ~n9394 ) ;
  assign n18162 = ( x113 & n18160 ) | ( x113 & ~n18161 ) | ( n18160 & ~n18161 ) ;
  assign n18163 = ( ~n18101 & n18159 ) | ( ~n18101 & n18162 ) | ( n18159 & n18162 ) ;
  assign n18164 = ( n18101 & n18159 ) | ( n18101 & n18162 ) | ( n18159 & n18162 ) ;
  assign n18165 = ( n18101 & n18163 ) | ( n18101 & ~n18164 ) | ( n18163 & ~n18164 ) ;
  assign n18166 = ( n18102 & ~n18149 ) | ( n18102 & n18165 ) | ( ~n18149 & n18165 ) ;
  assign n18167 = ( n18102 & n18149 ) | ( n18102 & ~n18165 ) | ( n18149 & ~n18165 ) ;
  assign n18168 = ( ~n18102 & n18166 ) | ( ~n18102 & n18167 ) | ( n18166 & n18167 ) ;
  assign n18169 = ( n18105 & n18139 ) | ( n18105 & ~n18168 ) | ( n18139 & ~n18168 ) ;
  assign n18170 = ( ~n18105 & n18139 ) | ( ~n18105 & n18168 ) | ( n18139 & n18168 ) ;
  assign n18171 = ( ~n18139 & n18169 ) | ( ~n18139 & n18170 ) | ( n18169 & n18170 ) ;
  assign n18172 = ( n18108 & n18129 ) | ( n18108 & ~n18171 ) | ( n18129 & ~n18171 ) ;
  assign n18173 = ( ~n18108 & n18129 ) | ( ~n18108 & n18171 ) | ( n18129 & n18171 ) ;
  assign n18174 = ( ~n18129 & n18172 ) | ( ~n18129 & n18173 ) | ( n18172 & n18173 ) ;
  assign n18175 = n6091 | n9864 ;
  assign n18176 = x127 & ~n5862 ;
  assign n18177 = n18175 & n18176 ;
  assign n18178 = x50 | n18177 ;
  assign n18179 = ~x49 & n18177 ;
  assign n18180 = n18178 & ~n18179 ;
  assign n18181 = ( n18111 & ~n18174 ) | ( n18111 & n18180 ) | ( ~n18174 & n18180 ) ;
  assign n18182 = ( n18111 & n18174 ) | ( n18111 & n18180 ) | ( n18174 & n18180 ) ;
  assign n18183 = ( n18174 & n18181 ) | ( n18174 & ~n18182 ) | ( n18181 & ~n18182 ) ;
  assign n18184 = ( ~n18115 & n18117 ) | ( ~n18115 & n18183 ) | ( n18117 & n18183 ) ;
  assign n18185 = ( n18115 & n18117 ) | ( n18115 & ~n18183 ) | ( n18117 & ~n18183 ) ;
  assign n18186 = ( ~n18117 & n18184 ) | ( ~n18117 & n18185 ) | ( n18184 & n18185 ) ;
  assign n18187 = n6546 & n9576 ;
  assign n18188 = x53 & n18187 ;
  assign n18189 = x127 & n6553 ;
  assign n18190 = x126 & n6550 ;
  assign n18191 = n18189 | n18190 ;
  assign n18192 = x125 & n6787 ;
  assign n18193 = n18191 | n18192 ;
  assign n18194 = ( ~x53 & n18187 ) | ( ~x53 & n18193 ) | ( n18187 & n18193 ) ;
  assign n18195 = x53 & ~n18193 ;
  assign n18196 = ( ~n18188 & n18194 ) | ( ~n18188 & n18195 ) | ( n18194 & n18195 ) ;
  assign n18197 = n7277 & n8729 ;
  assign n18198 = x56 & n18197 ;
  assign n18199 = x124 & n7545 ;
  assign n18200 = x123 & n7273 ;
  assign n18201 = n18199 | n18200 ;
  assign n18202 = x122 & n7552 ;
  assign n18203 = n18201 | n18202 ;
  assign n18204 = ( ~x56 & n18197 ) | ( ~x56 & n18203 ) | ( n18197 & n18203 ) ;
  assign n18205 = x56 & ~n18203 ;
  assign n18206 = ( ~n18198 & n18204 ) | ( ~n18198 & n18205 ) | ( n18204 & n18205 ) ;
  assign n18207 = n7696 & n8067 ;
  assign n18208 = x59 & n18207 ;
  assign n18209 = x121 & n8074 ;
  assign n18210 = x120 & n8071 ;
  assign n18211 = n18209 | n18210 ;
  assign n18212 = x119 & n8298 ;
  assign n18213 = n18211 | n18212 ;
  assign n18214 = ( ~x59 & n18207 ) | ( ~x59 & n18213 ) | ( n18207 & n18213 ) ;
  assign n18215 = x59 & ~n18213 ;
  assign n18216 = ( ~n18208 & n18214 ) | ( ~n18208 & n18215 ) | ( n18214 & n18215 ) ;
  assign n18217 = n6940 & n8859 ;
  assign n18218 = x62 & n18217 ;
  assign n18219 = x118 & n8866 ;
  assign n18220 = x117 & n8863 ;
  assign n18221 = n18219 | n18220 ;
  assign n18222 = x116 & n9125 ;
  assign n18223 = n18221 | n18222 ;
  assign n18224 = ( ~x62 & n18217 ) | ( ~x62 & n18223 ) | ( n18217 & n18223 ) ;
  assign n18225 = x62 & ~n18223 ;
  assign n18226 = ( ~n18218 & n18224 ) | ( ~n18218 & n18225 ) | ( n18224 & n18225 ) ;
  assign n18227 = ( x62 & x63 ) | ( x62 & x115 ) | ( x63 & x115 ) ;
  assign n18228 = ( x62 & x114 ) | ( x62 & ~n9394 ) | ( x114 & ~n9394 ) ;
  assign n18229 = ( x114 & n18227 ) | ( x114 & ~n18228 ) | ( n18227 & ~n18228 ) ;
  assign n18230 = ( x50 & n18101 ) | ( x50 & n18229 ) | ( n18101 & n18229 ) ;
  assign n18231 = ( ~x50 & n18101 ) | ( ~x50 & n18229 ) | ( n18101 & n18229 ) ;
  assign n18232 = ( x50 & ~n18230 ) | ( x50 & n18231 ) | ( ~n18230 & n18231 ) ;
  assign n18233 = ( n18163 & n18226 ) | ( n18163 & ~n18232 ) | ( n18226 & ~n18232 ) ;
  assign n18234 = ( n18163 & ~n18226 ) | ( n18163 & n18232 ) | ( ~n18226 & n18232 ) ;
  assign n18235 = ( ~n18163 & n18233 ) | ( ~n18163 & n18234 ) | ( n18233 & n18234 ) ;
  assign n18236 = ( n18167 & n18216 ) | ( n18167 & ~n18235 ) | ( n18216 & ~n18235 ) ;
  assign n18237 = ( n18167 & ~n18216 ) | ( n18167 & n18235 ) | ( ~n18216 & n18235 ) ;
  assign n18238 = ( ~n18167 & n18236 ) | ( ~n18167 & n18237 ) | ( n18236 & n18237 ) ;
  assign n18239 = ( n18169 & n18206 ) | ( n18169 & ~n18238 ) | ( n18206 & ~n18238 ) ;
  assign n18240 = ( n18169 & ~n18206 ) | ( n18169 & n18238 ) | ( ~n18206 & n18238 ) ;
  assign n18241 = ( ~n18169 & n18239 ) | ( ~n18169 & n18240 ) | ( n18239 & n18240 ) ;
  assign n18242 = ( n18172 & n18196 ) | ( n18172 & ~n18241 ) | ( n18196 & ~n18241 ) ;
  assign n18243 = ( n18172 & ~n18196 ) | ( n18172 & n18241 ) | ( ~n18196 & n18241 ) ;
  assign n18244 = ( ~n18172 & n18242 ) | ( ~n18172 & n18243 ) | ( n18242 & n18243 ) ;
  assign n18245 = ( ~n18181 & n18184 ) | ( ~n18181 & n18244 ) | ( n18184 & n18244 ) ;
  assign n18246 = ( n18181 & n18184 ) | ( n18181 & ~n18244 ) | ( n18184 & ~n18244 ) ;
  assign n18247 = ( ~n18184 & n18245 ) | ( ~n18184 & n18246 ) | ( n18245 & n18246 ) ;
  assign n18248 = x127 & n6550 ;
  assign n18249 = n6546 | n18248 ;
  assign n18250 = ( n9867 & n18248 ) | ( n9867 & n18249 ) | ( n18248 & n18249 ) ;
  assign n18251 = x126 & n6787 ;
  assign n18252 = ( ~x53 & n18250 ) | ( ~x53 & n18251 ) | ( n18250 & n18251 ) ;
  assign n18253 = ( x53 & ~n18250 ) | ( x53 & n18251 ) | ( ~n18250 & n18251 ) ;
  assign n18254 = ~n18251 & n18253 ;
  assign n18255 = n18252 | n18254 ;
  assign n18256 = n7277 & n9009 ;
  assign n18257 = x56 & n18256 ;
  assign n18258 = x125 & n7545 ;
  assign n18259 = x124 & n7273 ;
  assign n18260 = n18258 | n18259 ;
  assign n18261 = x123 & n7552 ;
  assign n18262 = n18260 | n18261 ;
  assign n18263 = ( ~x56 & n18256 ) | ( ~x56 & n18262 ) | ( n18256 & n18262 ) ;
  assign n18264 = x56 & ~n18262 ;
  assign n18265 = ( ~n18257 & n18263 ) | ( ~n18257 & n18264 ) | ( n18263 & n18264 ) ;
  assign n18266 = n8067 & n8207 ;
  assign n18267 = x59 & n18266 ;
  assign n18268 = x122 & n8074 ;
  assign n18269 = x121 & n8071 ;
  assign n18270 = n18268 | n18269 ;
  assign n18271 = x120 & n8298 ;
  assign n18272 = n18270 | n18271 ;
  assign n18273 = ( ~x59 & n18266 ) | ( ~x59 & n18272 ) | ( n18266 & n18272 ) ;
  assign n18274 = x59 & ~n18272 ;
  assign n18275 = ( ~n18267 & n18273 ) | ( ~n18267 & n18274 ) | ( n18273 & n18274 ) ;
  assign n18276 = ( x62 & x63 ) | ( x62 & x116 ) | ( x63 & x116 ) ;
  assign n18277 = ( x62 & x115 ) | ( x62 & ~n9394 ) | ( x115 & ~n9394 ) ;
  assign n18278 = ( x115 & n18276 ) | ( x115 & ~n18277 ) | ( n18276 & ~n18277 ) ;
  assign n18279 = n7181 & n8859 ;
  assign n18280 = x62 & n18279 ;
  assign n18281 = x119 & n8866 ;
  assign n18282 = x118 & n8863 ;
  assign n18283 = n18281 | n18282 ;
  assign n18284 = x117 & n9125 ;
  assign n18285 = n18283 | n18284 ;
  assign n18286 = ( ~x62 & n18279 ) | ( ~x62 & n18285 ) | ( n18279 & n18285 ) ;
  assign n18287 = x62 & ~n18285 ;
  assign n18288 = ( ~n18280 & n18286 ) | ( ~n18280 & n18287 ) | ( n18286 & n18287 ) ;
  assign n18289 = ( ~n18231 & n18278 ) | ( ~n18231 & n18288 ) | ( n18278 & n18288 ) ;
  assign n18290 = ( n18231 & n18278 ) | ( n18231 & ~n18288 ) | ( n18278 & ~n18288 ) ;
  assign n18291 = ( ~n18278 & n18289 ) | ( ~n18278 & n18290 ) | ( n18289 & n18290 ) ;
  assign n18292 = ( ~n18233 & n18275 ) | ( ~n18233 & n18291 ) | ( n18275 & n18291 ) ;
  assign n18293 = ( n18233 & n18275 ) | ( n18233 & ~n18291 ) | ( n18275 & ~n18291 ) ;
  assign n18294 = ( ~n18275 & n18292 ) | ( ~n18275 & n18293 ) | ( n18292 & n18293 ) ;
  assign n18295 = ( n18236 & n18265 ) | ( n18236 & ~n18294 ) | ( n18265 & ~n18294 ) ;
  assign n18296 = ( ~n18236 & n18265 ) | ( ~n18236 & n18294 ) | ( n18265 & n18294 ) ;
  assign n18297 = ( ~n18265 & n18295 ) | ( ~n18265 & n18296 ) | ( n18295 & n18296 ) ;
  assign n18298 = ( n18239 & n18255 ) | ( n18239 & ~n18297 ) | ( n18255 & ~n18297 ) ;
  assign n18299 = ( ~n18239 & n18255 ) | ( ~n18239 & n18297 ) | ( n18255 & n18297 ) ;
  assign n18300 = ( ~n18255 & n18298 ) | ( ~n18255 & n18299 ) | ( n18298 & n18299 ) ;
  assign n18301 = ( n18242 & n18245 ) | ( n18242 & ~n18300 ) | ( n18245 & ~n18300 ) ;
  assign n18302 = ( ~n18242 & n18245 ) | ( ~n18242 & n18300 ) | ( n18245 & n18300 ) ;
  assign n18303 = ( ~n18245 & n18301 ) | ( ~n18245 & n18302 ) | ( n18301 & n18302 ) ;
  assign n18304 = n6786 | n9864 ;
  assign n18305 = x127 & ~n6550 ;
  assign n18306 = n18304 & n18305 ;
  assign n18307 = x53 | n18306 ;
  assign n18308 = ~x52 & n18306 ;
  assign n18309 = n18307 & ~n18308 ;
  assign n18310 = n7277 & n9038 ;
  assign n18311 = x56 & n18310 ;
  assign n18312 = x126 & n7545 ;
  assign n18313 = x125 & n7273 ;
  assign n18314 = n18312 | n18313 ;
  assign n18315 = x124 & n7552 ;
  assign n18316 = n18314 | n18315 ;
  assign n18317 = ( ~x56 & n18310 ) | ( ~x56 & n18316 ) | ( n18310 & n18316 ) ;
  assign n18318 = x56 & ~n18316 ;
  assign n18319 = ( ~n18311 & n18317 ) | ( ~n18311 & n18318 ) | ( n18317 & n18318 ) ;
  assign n18320 = n8067 & n8461 ;
  assign n18321 = x59 & n18320 ;
  assign n18322 = x123 & n8074 ;
  assign n18323 = x122 & n8071 ;
  assign n18324 = n18322 | n18323 ;
  assign n18325 = x121 & n8298 ;
  assign n18326 = n18324 | n18325 ;
  assign n18327 = ( ~x59 & n18320 ) | ( ~x59 & n18326 ) | ( n18320 & n18326 ) ;
  assign n18328 = x59 & ~n18326 ;
  assign n18329 = ( ~n18321 & n18327 ) | ( ~n18321 & n18328 ) | ( n18327 & n18328 ) ;
  assign n18330 = n7444 & n8859 ;
  assign n18331 = x62 & n18330 ;
  assign n18332 = x120 & n8866 ;
  assign n18333 = x119 & n8863 ;
  assign n18334 = n18332 | n18333 ;
  assign n18335 = x118 & n9125 ;
  assign n18336 = n18334 | n18335 ;
  assign n18337 = ( ~x62 & n18330 ) | ( ~x62 & n18336 ) | ( n18330 & n18336 ) ;
  assign n18338 = x62 & ~n18336 ;
  assign n18339 = ( ~n18331 & n18337 ) | ( ~n18331 & n18338 ) | ( n18337 & n18338 ) ;
  assign n18340 = ( x62 & x63 ) | ( x62 & x117 ) | ( x63 & x117 ) ;
  assign n18341 = ( x62 & x116 ) | ( x62 & ~n9394 ) | ( x116 & ~n9394 ) ;
  assign n18342 = ( x116 & n18340 ) | ( x116 & ~n18341 ) | ( n18340 & ~n18341 ) ;
  assign n18343 = ( n18288 & ~n18290 ) | ( n18288 & n18342 ) | ( ~n18290 & n18342 ) ;
  assign n18344 = ( n18231 & n18289 ) | ( n18231 & ~n18342 ) | ( n18289 & ~n18342 ) ;
  assign n18345 = ( ~n18288 & n18343 ) | ( ~n18288 & n18344 ) | ( n18343 & n18344 ) ;
  assign n18346 = ( n18329 & n18339 ) | ( n18329 & ~n18345 ) | ( n18339 & ~n18345 ) ;
  assign n18347 = ( n18329 & ~n18339 ) | ( n18329 & n18345 ) | ( ~n18339 & n18345 ) ;
  assign n18348 = ( ~n18329 & n18346 ) | ( ~n18329 & n18347 ) | ( n18346 & n18347 ) ;
  assign n18349 = ( n18293 & n18319 ) | ( n18293 & ~n18348 ) | ( n18319 & ~n18348 ) ;
  assign n18350 = ( ~n18293 & n18319 ) | ( ~n18293 & n18348 ) | ( n18319 & n18348 ) ;
  assign n18351 = ( ~n18319 & n18349 ) | ( ~n18319 & n18350 ) | ( n18349 & n18350 ) ;
  assign n18352 = ( n18295 & ~n18309 ) | ( n18295 & n18351 ) | ( ~n18309 & n18351 ) ;
  assign n18353 = ( n18295 & n18309 ) | ( n18295 & ~n18351 ) | ( n18309 & ~n18351 ) ;
  assign n18354 = ( ~n18295 & n18352 ) | ( ~n18295 & n18353 ) | ( n18352 & n18353 ) ;
  assign n18355 = ( ~n18298 & n18302 ) | ( ~n18298 & n18354 ) | ( n18302 & n18354 ) ;
  assign n18356 = ( n18298 & n18302 ) | ( n18298 & ~n18354 ) | ( n18302 & ~n18354 ) ;
  assign n18357 = ( ~n18302 & n18355 ) | ( ~n18302 & n18356 ) | ( n18355 & n18356 ) ;
  assign n18358 = n7277 & n9576 ;
  assign n18359 = x56 & n18358 ;
  assign n18360 = x127 & n7545 ;
  assign n18361 = x126 & n7273 ;
  assign n18362 = n18360 | n18361 ;
  assign n18363 = x125 & n7552 ;
  assign n18364 = n18362 | n18363 ;
  assign n18365 = ( ~x56 & n18358 ) | ( ~x56 & n18364 ) | ( n18358 & n18364 ) ;
  assign n18366 = x56 & ~n18364 ;
  assign n18367 = ( ~n18359 & n18365 ) | ( ~n18359 & n18366 ) | ( n18365 & n18366 ) ;
  assign n18368 = n8067 & n8729 ;
  assign n18369 = x59 & n18368 ;
  assign n18370 = x124 & n8074 ;
  assign n18371 = x123 & n8071 ;
  assign n18372 = n18370 | n18371 ;
  assign n18373 = x122 & n8298 ;
  assign n18374 = n18372 | n18373 ;
  assign n18375 = ( ~x59 & n18368 ) | ( ~x59 & n18374 ) | ( n18368 & n18374 ) ;
  assign n18376 = x59 & ~n18374 ;
  assign n18377 = ( ~n18369 & n18375 ) | ( ~n18369 & n18376 ) | ( n18375 & n18376 ) ;
  assign n18378 = n7696 & n8859 ;
  assign n18379 = x62 & n18378 ;
  assign n18380 = x121 & n8866 ;
  assign n18381 = x120 & n8863 ;
  assign n18382 = n18380 | n18381 ;
  assign n18383 = x119 & n9125 ;
  assign n18384 = n18382 | n18383 ;
  assign n18385 = ( ~x62 & n18378 ) | ( ~x62 & n18384 ) | ( n18378 & n18384 ) ;
  assign n18386 = x62 & ~n18384 ;
  assign n18387 = ( ~n18379 & n18385 ) | ( ~n18379 & n18386 ) | ( n18385 & n18386 ) ;
  assign n18388 = ( x62 & x63 ) | ( x62 & x118 ) | ( x63 & x118 ) ;
  assign n18389 = ( x62 & x117 ) | ( x62 & ~n9394 ) | ( x117 & ~n9394 ) ;
  assign n18390 = ( x117 & n18388 ) | ( x117 & ~n18389 ) | ( n18388 & ~n18389 ) ;
  assign n18391 = ( x53 & n18342 ) | ( x53 & n18390 ) | ( n18342 & n18390 ) ;
  assign n18392 = ( ~x53 & n18342 ) | ( ~x53 & n18390 ) | ( n18342 & n18390 ) ;
  assign n18393 = ( x53 & ~n18391 ) | ( x53 & n18392 ) | ( ~n18391 & n18392 ) ;
  assign n18394 = ( n18344 & n18387 ) | ( n18344 & ~n18393 ) | ( n18387 & ~n18393 ) ;
  assign n18395 = ( ~n18344 & n18387 ) | ( ~n18344 & n18393 ) | ( n18387 & n18393 ) ;
  assign n18396 = ( ~n18387 & n18394 ) | ( ~n18387 & n18395 ) | ( n18394 & n18395 ) ;
  assign n18397 = ( n18346 & n18377 ) | ( n18346 & ~n18396 ) | ( n18377 & ~n18396 ) ;
  assign n18398 = ( n18346 & ~n18377 ) | ( n18346 & n18396 ) | ( ~n18377 & n18396 ) ;
  assign n18399 = ( ~n18346 & n18397 ) | ( ~n18346 & n18398 ) | ( n18397 & n18398 ) ;
  assign n18400 = ( n18349 & n18367 ) | ( n18349 & ~n18399 ) | ( n18367 & ~n18399 ) ;
  assign n18401 = ( n18349 & ~n18367 ) | ( n18349 & n18399 ) | ( ~n18367 & n18399 ) ;
  assign n18402 = ( ~n18349 & n18400 ) | ( ~n18349 & n18401 ) | ( n18400 & n18401 ) ;
  assign n18403 = ( ~n18353 & n18355 ) | ( ~n18353 & n18402 ) | ( n18355 & n18402 ) ;
  assign n18404 = ( n18353 & n18355 ) | ( n18353 & ~n18402 ) | ( n18355 & ~n18402 ) ;
  assign n18405 = ( ~n18355 & n18403 ) | ( ~n18355 & n18404 ) | ( n18403 & n18404 ) ;
  assign n18406 = x127 & n7273 ;
  assign n18407 = n7277 | n18406 ;
  assign n18408 = ( n9867 & n18406 ) | ( n9867 & n18407 ) | ( n18406 & n18407 ) ;
  assign n18409 = x126 & n7552 ;
  assign n18410 = ( ~x56 & n18408 ) | ( ~x56 & n18409 ) | ( n18408 & n18409 ) ;
  assign n18411 = ( x56 & ~n18408 ) | ( x56 & n18409 ) | ( ~n18408 & n18409 ) ;
  assign n18412 = ~n18409 & n18411 ;
  assign n18413 = n18410 | n18412 ;
  assign n18414 = n8067 & n9009 ;
  assign n18415 = x59 & n18414 ;
  assign n18416 = x125 & n8074 ;
  assign n18417 = x124 & n8071 ;
  assign n18418 = n18416 | n18417 ;
  assign n18419 = x123 & n8298 ;
  assign n18420 = n18418 | n18419 ;
  assign n18421 = ( ~x59 & n18414 ) | ( ~x59 & n18420 ) | ( n18414 & n18420 ) ;
  assign n18422 = x59 & ~n18420 ;
  assign n18423 = ( ~n18415 & n18421 ) | ( ~n18415 & n18422 ) | ( n18421 & n18422 ) ;
  assign n18424 = n8207 & n8859 ;
  assign n18425 = x62 & n18424 ;
  assign n18426 = x122 & n8866 ;
  assign n18427 = x121 & n8863 ;
  assign n18428 = n18426 | n18427 ;
  assign n18429 = x120 & n9125 ;
  assign n18430 = n18428 | n18429 ;
  assign n18431 = ( ~x62 & n18424 ) | ( ~x62 & n18430 ) | ( n18424 & n18430 ) ;
  assign n18432 = x62 & ~n18430 ;
  assign n18433 = ( ~n18425 & n18431 ) | ( ~n18425 & n18432 ) | ( n18431 & n18432 ) ;
  assign n18434 = ( x62 & x63 ) | ( x62 & x119 ) | ( x63 & x119 ) ;
  assign n18435 = ( x62 & x118 ) | ( x62 & ~n9394 ) | ( x118 & ~n9394 ) ;
  assign n18436 = ( x118 & n18434 ) | ( x118 & ~n18435 ) | ( n18434 & ~n18435 ) ;
  assign n18437 = ( n18392 & n18433 ) | ( n18392 & ~n18436 ) | ( n18433 & ~n18436 ) ;
  assign n18438 = ( ~n18392 & n18433 ) | ( ~n18392 & n18436 ) | ( n18433 & n18436 ) ;
  assign n18439 = ( ~n18433 & n18437 ) | ( ~n18433 & n18438 ) | ( n18437 & n18438 ) ;
  assign n18440 = ( ~n18394 & n18423 ) | ( ~n18394 & n18439 ) | ( n18423 & n18439 ) ;
  assign n18441 = ( n18394 & n18423 ) | ( n18394 & ~n18439 ) | ( n18423 & ~n18439 ) ;
  assign n18442 = ( ~n18423 & n18440 ) | ( ~n18423 & n18441 ) | ( n18440 & n18441 ) ;
  assign n18443 = ( n18397 & n18413 ) | ( n18397 & ~n18442 ) | ( n18413 & ~n18442 ) ;
  assign n18444 = ( ~n18397 & n18413 ) | ( ~n18397 & n18442 ) | ( n18413 & n18442 ) ;
  assign n18445 = ( ~n18413 & n18443 ) | ( ~n18413 & n18444 ) | ( n18443 & n18444 ) ;
  assign n18446 = ( ~n18400 & n18403 ) | ( ~n18400 & n18445 ) | ( n18403 & n18445 ) ;
  assign n18447 = ( n18400 & n18403 ) | ( n18400 & ~n18445 ) | ( n18403 & ~n18445 ) ;
  assign n18448 = ( ~n18403 & n18446 ) | ( ~n18403 & n18447 ) | ( n18446 & n18447 ) ;
  assign n18449 = n8067 & n9038 ;
  assign n18450 = x59 & n18449 ;
  assign n18451 = x126 & n8074 ;
  assign n18452 = x125 & n8071 ;
  assign n18453 = n18451 | n18452 ;
  assign n18454 = x124 & n8298 ;
  assign n18455 = n18453 | n18454 ;
  assign n18456 = ( ~x59 & n18449 ) | ( ~x59 & n18455 ) | ( n18449 & n18455 ) ;
  assign n18457 = x59 & ~n18455 ;
  assign n18458 = ( ~n18450 & n18456 ) | ( ~n18450 & n18457 ) | ( n18456 & n18457 ) ;
  assign n18459 = n8461 & n8859 ;
  assign n18460 = x62 & n18459 ;
  assign n18461 = x123 & n8866 ;
  assign n18462 = x122 & n8863 ;
  assign n18463 = n18461 | n18462 ;
  assign n18464 = x121 & n9125 ;
  assign n18465 = n18463 | n18464 ;
  assign n18466 = ( ~x62 & n18459 ) | ( ~x62 & n18465 ) | ( n18459 & n18465 ) ;
  assign n18467 = x62 & ~n18465 ;
  assign n18468 = ( ~n18460 & n18466 ) | ( ~n18460 & n18467 ) | ( n18466 & n18467 ) ;
  assign n18469 = ( x62 & x63 ) | ( x62 & x120 ) | ( x63 & x120 ) ;
  assign n18470 = ( x62 & x119 ) | ( x62 & ~n9394 ) | ( x119 & ~n9394 ) ;
  assign n18471 = ( x119 & n18469 ) | ( x119 & ~n18470 ) | ( n18469 & ~n18470 ) ;
  assign n18472 = ( ~n18436 & n18468 ) | ( ~n18436 & n18471 ) | ( n18468 & n18471 ) ;
  assign n18473 = ( n18436 & n18468 ) | ( n18436 & n18471 ) | ( n18468 & n18471 ) ;
  assign n18474 = ( n18436 & n18472 ) | ( n18436 & ~n18473 ) | ( n18472 & ~n18473 ) ;
  assign n18475 = ( ~n18437 & n18458 ) | ( ~n18437 & n18474 ) | ( n18458 & n18474 ) ;
  assign n18476 = ( n18437 & n18458 ) | ( n18437 & ~n18474 ) | ( n18458 & ~n18474 ) ;
  assign n18477 = ( ~n18458 & n18475 ) | ( ~n18458 & n18476 ) | ( n18475 & n18476 ) ;
  assign n18478 = x55 & ~n7273 ;
  assign n18479 = ( x127 & n7551 ) | ( x127 & n9865 ) | ( n7551 & n9865 ) ;
  assign n18480 = ~n18478 & n18479 ;
  assign n18481 = ( n7273 & n18478 ) | ( n7273 & n18479 ) | ( n18478 & n18479 ) ;
  assign n18482 = ( x56 & ~n18480 ) | ( x56 & n18481 ) | ( ~n18480 & n18481 ) ;
  assign n18483 = ( n18441 & ~n18477 ) | ( n18441 & n18482 ) | ( ~n18477 & n18482 ) ;
  assign n18484 = ( n18441 & n18477 ) | ( n18441 & n18482 ) | ( n18477 & n18482 ) ;
  assign n18485 = ( n18477 & n18483 ) | ( n18477 & ~n18484 ) | ( n18483 & ~n18484 ) ;
  assign n18486 = ( ~n18443 & n18446 ) | ( ~n18443 & n18485 ) | ( n18446 & n18485 ) ;
  assign n18487 = ( n18443 & n18446 ) | ( n18443 & ~n18485 ) | ( n18446 & ~n18485 ) ;
  assign n18488 = ( ~n18446 & n18486 ) | ( ~n18446 & n18487 ) | ( n18486 & n18487 ) ;
  assign n18489 = x127 & n8074 ;
  assign n18490 = n8067 | n18489 ;
  assign n18491 = ( n9576 & n18489 ) | ( n9576 & n18490 ) | ( n18489 & n18490 ) ;
  assign n18492 = x125 & n8298 ;
  assign n18493 = n18491 | n18492 ;
  assign n18494 = x126 & n8071 ;
  assign n18495 = ( ~x59 & n18493 ) | ( ~x59 & n18494 ) | ( n18493 & n18494 ) ;
  assign n18496 = ( x59 & ~n18493 ) | ( x59 & n18494 ) | ( ~n18493 & n18494 ) ;
  assign n18497 = ~n18494 & n18496 ;
  assign n18498 = n18495 | n18497 ;
  assign n18499 = n8729 & n8859 ;
  assign n18500 = x62 & n18499 ;
  assign n18501 = x124 & n8866 ;
  assign n18502 = x123 & n8863 ;
  assign n18503 = n18501 | n18502 ;
  assign n18504 = x122 & n9125 ;
  assign n18505 = n18503 | n18504 ;
  assign n18506 = ( ~x62 & n18499 ) | ( ~x62 & n18505 ) | ( n18499 & n18505 ) ;
  assign n18507 = x62 & ~n18505 ;
  assign n18508 = ( ~n18500 & n18506 ) | ( ~n18500 & n18507 ) | ( n18506 & n18507 ) ;
  assign n18509 = ( x62 & x63 ) | ( x62 & x121 ) | ( x63 & x121 ) ;
  assign n18510 = ( x62 & x120 ) | ( x62 & ~n9394 ) | ( x120 & ~n9394 ) ;
  assign n18511 = ( x120 & n18509 ) | ( x120 & ~n18510 ) | ( n18509 & ~n18510 ) ;
  assign n18512 = ( x56 & n18436 ) | ( x56 & n18511 ) | ( n18436 & n18511 ) ;
  assign n18513 = ( ~x56 & n18436 ) | ( ~x56 & n18511 ) | ( n18436 & n18511 ) ;
  assign n18514 = ( x56 & ~n18512 ) | ( x56 & n18513 ) | ( ~n18512 & n18513 ) ;
  assign n18515 = ( n18472 & n18508 ) | ( n18472 & ~n18514 ) | ( n18508 & ~n18514 ) ;
  assign n18516 = ( n18472 & ~n18508 ) | ( n18472 & n18514 ) | ( ~n18508 & n18514 ) ;
  assign n18517 = ( ~n18472 & n18515 ) | ( ~n18472 & n18516 ) | ( n18515 & n18516 ) ;
  assign n18518 = ( n18476 & n18498 ) | ( n18476 & ~n18517 ) | ( n18498 & ~n18517 ) ;
  assign n18519 = ( ~n18476 & n18498 ) | ( ~n18476 & n18517 ) | ( n18498 & n18517 ) ;
  assign n18520 = ( ~n18498 & n18518 ) | ( ~n18498 & n18519 ) | ( n18518 & n18519 ) ;
  assign n18521 = ( ~n18483 & n18486 ) | ( ~n18483 & n18520 ) | ( n18486 & n18520 ) ;
  assign n18522 = ( n18483 & n18486 ) | ( n18483 & ~n18520 ) | ( n18486 & ~n18520 ) ;
  assign n18523 = ( ~n18486 & n18521 ) | ( ~n18486 & n18522 ) | ( n18521 & n18522 ) ;
  assign n18524 = x127 & n8071 ;
  assign n18525 = n8067 | n18524 ;
  assign n18526 = ( n9867 & n18524 ) | ( n9867 & n18525 ) | ( n18524 & n18525 ) ;
  assign n18527 = x126 & n8298 ;
  assign n18528 = ( ~x59 & n18526 ) | ( ~x59 & n18527 ) | ( n18526 & n18527 ) ;
  assign n18529 = ( x59 & ~n18526 ) | ( x59 & n18527 ) | ( ~n18526 & n18527 ) ;
  assign n18530 = ~n18527 & n18529 ;
  assign n18531 = n18528 | n18530 ;
  assign n18532 = ( x62 & x63 ) | ( x62 & x122 ) | ( x63 & x122 ) ;
  assign n18533 = ( x62 & x121 ) | ( x62 & ~n9394 ) | ( x121 & ~n9394 ) ;
  assign n18534 = ( x121 & n18532 ) | ( x121 & ~n18533 ) | ( n18532 & ~n18533 ) ;
  assign n18535 = n8859 & n9009 ;
  assign n18536 = x62 & n18535 ;
  assign n18537 = x125 & n8866 ;
  assign n18538 = x124 & n8863 ;
  assign n18539 = n18537 | n18538 ;
  assign n18540 = x123 & n9125 ;
  assign n18541 = n18539 | n18540 ;
  assign n18542 = ( ~x62 & n18535 ) | ( ~x62 & n18541 ) | ( n18535 & n18541 ) ;
  assign n18543 = x62 & ~n18541 ;
  assign n18544 = ( ~n18536 & n18542 ) | ( ~n18536 & n18543 ) | ( n18542 & n18543 ) ;
  assign n18545 = ( ~n18513 & n18534 ) | ( ~n18513 & n18544 ) | ( n18534 & n18544 ) ;
  assign n18546 = ( n18513 & n18534 ) | ( n18513 & ~n18544 ) | ( n18534 & ~n18544 ) ;
  assign n18547 = ( ~n18534 & n18545 ) | ( ~n18534 & n18546 ) | ( n18545 & n18546 ) ;
  assign n18548 = ( n18515 & n18531 ) | ( n18515 & ~n18547 ) | ( n18531 & ~n18547 ) ;
  assign n18549 = ( ~n18515 & n18531 ) | ( ~n18515 & n18547 ) | ( n18531 & n18547 ) ;
  assign n18550 = ( ~n18531 & n18548 ) | ( ~n18531 & n18549 ) | ( n18548 & n18549 ) ;
  assign n18551 = ( ~n18518 & n18521 ) | ( ~n18518 & n18550 ) | ( n18521 & n18550 ) ;
  assign n18552 = ( n18518 & n18521 ) | ( n18518 & ~n18550 ) | ( n18521 & ~n18550 ) ;
  assign n18553 = ( ~n18521 & n18551 ) | ( ~n18521 & n18552 ) | ( n18551 & n18552 ) ;
  assign n18554 = n8297 | n9864 ;
  assign n18555 = x127 & ~n8071 ;
  assign n18556 = n18554 & n18555 ;
  assign n18557 = x59 | n18556 ;
  assign n18558 = ~x58 & n18556 ;
  assign n18559 = n18557 & ~n18558 ;
  assign n18560 = ( x62 & x63 ) | ( x62 & x123 ) | ( x63 & x123 ) ;
  assign n18561 = ( x62 & x122 ) | ( x62 & ~n9394 ) | ( x122 & ~n9394 ) ;
  assign n18562 = ( x122 & n18560 ) | ( x122 & ~n18561 ) | ( n18560 & ~n18561 ) ;
  assign n18563 = ( n18544 & ~n18546 ) | ( n18544 & n18562 ) | ( ~n18546 & n18562 ) ;
  assign n18564 = ( n18513 & n18545 ) | ( n18513 & ~n18562 ) | ( n18545 & ~n18562 ) ;
  assign n18565 = ( ~n18544 & n18563 ) | ( ~n18544 & n18564 ) | ( n18563 & n18564 ) ;
  assign n18566 = n8859 & n9038 ;
  assign n18567 = x62 & n18566 ;
  assign n18568 = x126 & n8866 ;
  assign n18569 = x125 & n8863 ;
  assign n18570 = n18568 | n18569 ;
  assign n18571 = x124 & n9125 ;
  assign n18572 = n18570 | n18571 ;
  assign n18573 = ( ~x62 & n18566 ) | ( ~x62 & n18572 ) | ( n18566 & n18572 ) ;
  assign n18574 = x62 & ~n18572 ;
  assign n18575 = ( ~n18567 & n18573 ) | ( ~n18567 & n18574 ) | ( n18573 & n18574 ) ;
  assign n18576 = ( n18559 & ~n18565 ) | ( n18559 & n18575 ) | ( ~n18565 & n18575 ) ;
  assign n18577 = ( n18559 & n18565 ) | ( n18559 & ~n18575 ) | ( n18565 & ~n18575 ) ;
  assign n18578 = ( ~n18559 & n18576 ) | ( ~n18559 & n18577 ) | ( n18576 & n18577 ) ;
  assign n18579 = ( ~n18548 & n18551 ) | ( ~n18548 & n18578 ) | ( n18551 & n18578 ) ;
  assign n18580 = ( n18548 & n18551 ) | ( n18548 & ~n18578 ) | ( n18551 & ~n18578 ) ;
  assign n18581 = ( ~n18551 & n18579 ) | ( ~n18551 & n18580 ) | ( n18579 & n18580 ) ;
  assign n18582 = ~n18544 & n18562 ;
  assign n18583 = ( n18513 & n18534 ) | ( n18513 & ~n18562 ) | ( n18534 & ~n18562 ) ;
  assign n18584 = n18562 & n18583 ;
  assign n18585 = n18544 | n18583 ;
  assign n18586 = ( n18582 & ~n18584 ) | ( n18582 & n18585 ) | ( ~n18584 & n18585 ) ;
  assign n18587 = ( x62 & x63 ) | ( x62 & x124 ) | ( x63 & x124 ) ;
  assign n18588 = ( x62 & x123 ) | ( x62 & ~n9394 ) | ( x123 & ~n9394 ) ;
  assign n18589 = ( x123 & n18587 ) | ( x123 & ~n18588 ) | ( n18587 & ~n18588 ) ;
  assign n18590 = x62 & ~n18589 ;
  assign n18591 = x62 | x124 ;
  assign n18592 = ( n9395 & n18590 ) | ( n9395 & n18591 ) | ( n18590 & n18591 ) ;
  assign n18593 = ( ~x59 & n18586 ) | ( ~x59 & n18592 ) | ( n18586 & n18592 ) ;
  assign n18594 = ( x59 & n18586 ) | ( x59 & n18592 ) | ( n18586 & n18592 ) ;
  assign n18595 = ( x59 & n18593 ) | ( x59 & ~n18594 ) | ( n18593 & ~n18594 ) ;
  assign n18596 = x127 & n8866 ;
  assign n18597 = x125 & n9125 ;
  assign n18598 = n18596 | n18597 ;
  assign n18599 = n8859 | n18598 ;
  assign n18600 = ( n9576 & n18598 ) | ( n9576 & n18599 ) | ( n18598 & n18599 ) ;
  assign n18601 = x126 & n8863 ;
  assign n18602 = n18600 | n18601 ;
  assign n18603 = n18595 | n18602 ;
  assign n18604 = n18595 & n18602 ;
  assign n18605 = n18603 & ~n18604 ;
  assign n18606 = ( ~n18576 & n18579 ) | ( ~n18576 & n18605 ) | ( n18579 & n18605 ) ;
  assign n18607 = ( n18576 & n18579 ) | ( n18576 & ~n18605 ) | ( n18579 & ~n18605 ) ;
  assign n18608 = ( ~n18579 & n18606 ) | ( ~n18579 & n18607 ) | ( n18606 & n18607 ) ;
  assign n18609 = ( x62 & ~n18564 ) | ( x62 & n18595 ) | ( ~n18564 & n18595 ) ;
  assign n18610 = ( x62 & n18564 ) | ( x62 & n18595 ) | ( n18564 & n18595 ) ;
  assign n18611 = ( n18605 & ~n18609 ) | ( n18605 & n18610 ) | ( ~n18609 & n18610 ) ;
  assign n18612 = ( x62 & x63 ) | ( x62 & x125 ) | ( x63 & x125 ) ;
  assign n18613 = ( x62 & x124 ) | ( x62 & ~n9394 ) | ( x124 & ~n9394 ) ;
  assign n18614 = ( x124 & n18612 ) | ( x124 & ~n18613 ) | ( n18612 & ~n18613 ) ;
  assign n18615 = x127 & n8863 ;
  assign n18616 = n8859 | n18615 ;
  assign n18617 = ( n9867 & n18615 ) | ( n9867 & n18616 ) | ( n18615 & n18616 ) ;
  assign n18618 = x126 & n9125 ;
  assign n18619 = ( ~x62 & n18617 ) | ( ~x62 & n18618 ) | ( n18617 & n18618 ) ;
  assign n18620 = ( x62 & ~n18617 ) | ( x62 & n18618 ) | ( ~n18617 & n18618 ) ;
  assign n18621 = ~n18618 & n18620 ;
  assign n18622 = n18619 | n18621 ;
  assign n18623 = ( ~x59 & n18562 ) | ( ~x59 & n18589 ) | ( n18562 & n18589 ) ;
  assign n18624 = ( n18614 & n18622 ) | ( n18614 & n18623 ) | ( n18622 & n18623 ) ;
  assign n18625 = ( ~n18614 & n18622 ) | ( ~n18614 & n18623 ) | ( n18622 & n18623 ) ;
  assign n18626 = ( n18614 & ~n18624 ) | ( n18614 & n18625 ) | ( ~n18624 & n18625 ) ;
  assign n18627 = ( n18606 & n18611 ) | ( n18606 & ~n18626 ) | ( n18611 & ~n18626 ) ;
  assign n18628 = ( n18606 & ~n18611 ) | ( n18606 & n18626 ) | ( ~n18611 & n18626 ) ;
  assign n18629 = ( ~n18606 & n18627 ) | ( ~n18606 & n18628 ) | ( n18627 & n18628 ) ;
  assign n18630 = ( x62 & x63 ) | ( x62 & x126 ) | ( x63 & x126 ) ;
  assign n18631 = ( x62 & x125 ) | ( x62 & ~n9394 ) | ( x125 & ~n9394 ) ;
  assign n18632 = ( x125 & n18630 ) | ( x125 & ~n18631 ) | ( n18630 & ~n18631 ) ;
  assign n18633 = n9124 | n9864 ;
  assign n18634 = x127 & ~n8863 ;
  assign n18635 = n18633 & n18634 ;
  assign n18636 = x62 | n18635 ;
  assign n18637 = ~x61 & n18635 ;
  assign n18638 = n18636 & ~n18637 ;
  assign n18639 = ( n18614 & n18632 ) | ( n18614 & ~n18638 ) | ( n18632 & ~n18638 ) ;
  assign n18640 = ( ~n18614 & n18632 ) | ( ~n18614 & n18638 ) | ( n18632 & n18638 ) ;
  assign n18641 = ( ~n18632 & n18639 ) | ( ~n18632 & n18640 ) | ( n18639 & n18640 ) ;
  assign n18642 = ( ~n18625 & n18628 ) | ( ~n18625 & n18641 ) | ( n18628 & n18641 ) ;
  assign n18643 = ( n18625 & n18628 ) | ( n18625 & ~n18641 ) | ( n18628 & ~n18641 ) ;
  assign n18644 = ( ~n18628 & n18642 ) | ( ~n18628 & n18643 ) | ( n18642 & n18643 ) ;
  assign n18645 = ( x63 & ~x125 ) | ( x63 & x127 ) | ( ~x125 & x127 ) ;
  assign n18646 = ( x62 & x63 ) | ( x62 & ~n18645 ) | ( x63 & ~n18645 ) ;
  assign n18647 = x125 & n18645 ;
  assign n18648 = ( x127 & n18646 ) | ( x127 & ~n18647 ) | ( n18646 & ~n18647 ) ;
  assign n18649 = ( x63 & x126 ) | ( x63 & x127 ) | ( x126 & x127 ) ;
  assign n18650 = ( n9863 & n18614 ) | ( n9863 & n18649 ) | ( n18614 & n18649 ) ;
  assign n18651 = ( n9863 & ~n18614 ) | ( n9863 & n18649 ) | ( ~n18614 & n18649 ) ;
  assign n18652 = ( n18614 & ~n18650 ) | ( n18614 & n18651 ) | ( ~n18650 & n18651 ) ;
  assign n18653 = x125 | x127 ;
  assign n18654 = n9395 & n18653 ;
  assign n18655 = n18648 & n18654 ;
  assign n18656 = ( n18648 & ~n18652 ) | ( n18648 & n18655 ) | ( ~n18652 & n18655 ) ;
  assign n18657 = ( ~n18640 & n18642 ) | ( ~n18640 & n18656 ) | ( n18642 & n18656 ) ;
  assign n18658 = ( n18640 & n18642 ) | ( n18640 & ~n18656 ) | ( n18642 & ~n18656 ) ;
  assign n18659 = ( ~n18642 & n18657 ) | ( ~n18642 & n18658 ) | ( n18657 & n18658 ) ;
  assign n18660 = x63 & x126 ;
  assign n18661 = n18614 & n18660 ;
  assign n18662 = x127 & n18646 ;
  assign n18663 = ( n18654 & ~n18661 ) | ( n18654 & n18662 ) | ( ~n18661 & n18662 ) ;
  assign n18664 = ( n18654 & n18661 ) | ( n18654 & ~n18662 ) | ( n18661 & ~n18662 ) ;
  assign n18665 = n18663 | n18664 ;
  assign n18666 = ~n18657 & n18665 ;
  assign n18667 = n18657 & ~n18665 ;
  assign n18668 = n18666 | n18667 ;
  assign y0 = n129 ;
  assign y1 = n134 ;
  assign y2 = n158 ;
  assign y3 = n184 ;
  assign y4 = n218 ;
  assign y5 = n253 ;
  assign y6 = n289 ;
  assign y7 = n335 ;
  assign y8 = n385 ;
  assign y9 = n433 ;
  assign y10 = n491 ;
  assign y11 = n561 ;
  assign y12 = n623 ;
  assign y13 = n694 ;
  assign y14 = n763 ;
  assign y15 = n837 ;
  assign y16 = n922 ;
  assign y17 = n1003 ;
  assign y18 = n1090 ;
  assign y19 = n1187 ;
  assign y20 = n1282 ;
  assign y21 = n1381 ;
  assign y22 = n1491 ;
  assign y23 = n1599 ;
  assign y24 = n1711 ;
  assign y25 = n1835 ;
  assign y26 = n1956 ;
  assign y27 = n2080 ;
  assign y28 = n2217 ;
  assign y29 = n2351 ;
  assign y30 = n2489 ;
  assign y31 = n2638 ;
  assign y32 = n2785 ;
  assign y33 = n2936 ;
  assign y34 = n3098 ;
  assign y35 = n3261 ;
  assign y36 = n3429 ;
  assign y37 = n3604 ;
  assign y38 = n3777 ;
  assign y39 = n3954 ;
  assign y40 = n4142 ;
  assign y41 = n4328 ;
  assign y42 = n4520 ;
  assign y43 = n4727 ;
  assign y44 = n4927 ;
  assign y45 = n5129 ;
  assign y46 = n5344 ;
  assign y47 = n5555 ;
  assign y48 = n5771 ;
  assign y49 = n5999 ;
  assign y50 = n6226 ;
  assign y51 = n6459 ;
  assign y52 = n6700 ;
  assign y53 = n6937 ;
  assign y54 = n7178 ;
  assign y55 = n7441 ;
  assign y56 = n7693 ;
  assign y57 = n7949 ;
  assign y58 = n8220 ;
  assign y59 = n8487 ;
  assign y60 = n8755 ;
  assign y61 = n9035 ;
  assign y62 = n9311 ;
  assign y63 = n9592 ;
  assign y64 = n9877 ;
  assign y65 = n10148 ;
  assign y66 = n10414 ;
  assign y67 = n10678 ;
  assign y68 = n10940 ;
  assign y69 = n11196 ;
  assign y70 = n11447 ;
  assign y71 = n11696 ;
  assign y72 = n11939 ;
  assign y73 = n12177 ;
  assign y74 = n12414 ;
  assign y75 = n12644 ;
  assign y76 = n12869 ;
  assign y77 = n13092 ;
  assign y78 = n13309 ;
  assign y79 = n13521 ;
  assign y80 = n13731 ;
  assign y81 = n13935 ;
  assign y82 = n14134 ;
  assign y83 = n14331 ;
  assign y84 = n14522 ;
  assign y85 = n14708 ;
  assign y86 = n14892 ;
  assign y87 = n15070 ;
  assign y88 = n15243 ;
  assign y89 = n15413 ;
  assign y90 = n15578 ;
  assign y91 = n15738 ;
  assign y92 = n15896 ;
  assign y93 = n16048 ;
  assign y94 = n16195 ;
  assign y95 = n16340 ;
  assign y96 = n16479 ;
  assign y97 = n16613 ;
  assign y98 = n16745 ;
  assign y99 = n16871 ;
  assign y100 = n16992 ;
  assign y101 = n17112 ;
  assign y102 = n17225 ;
  assign y103 = n17333 ;
  assign y104 = n17440 ;
  assign y105 = n17540 ;
  assign y106 = n17635 ;
  assign y107 = n17727 ;
  assign y108 = n17814 ;
  assign y109 = n17896 ;
  assign y110 = n17976 ;
  assign y111 = n18050 ;
  assign y112 = n18119 ;
  assign y113 = n18186 ;
  assign y114 = n18247 ;
  assign y115 = n18303 ;
  assign y116 = n18357 ;
  assign y117 = n18405 ;
  assign y118 = n18448 ;
  assign y119 = n18488 ;
  assign y120 = n18523 ;
  assign y121 = n18553 ;
  assign y122 = n18581 ;
  assign y123 = n18608 ;
  assign y124 = n18629 ;
  assign y125 = n18644 ;
  assign y126 = n18659 ;
  assign y127 = n18668 ;
endmodule
