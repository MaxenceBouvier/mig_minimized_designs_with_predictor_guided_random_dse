module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 ;
  assign n12 = x6 & x7 ;
  assign n13 = x10 & n12 ;
  assign n14 = x8 & x9 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = x6 | x7 ;
  assign n17 = x10 & n16 ;
  assign n18 = x5 & x6 ;
  assign n19 = x9 & ~x10 ;
  assign n20 = ( x5 & x6 ) | ( x5 & n19 ) | ( x6 & n19 ) ;
  assign n21 = ( n17 & ~n18 ) | ( n17 & n20 ) | ( ~n18 & n20 ) ;
  assign n22 = ~n15 & n21 ;
  assign n23 = x4 & x5 ;
  assign n24 = ( x4 & x5 ) | ( x4 & x8 ) | ( x5 & x8 ) ;
  assign n25 = ( x2 & ~x3 ) | ( x2 & x6 ) | ( ~x3 & x6 ) ;
  assign n26 = ( x2 & ~x3 ) | ( x2 & x7 ) | ( ~x3 & x7 ) ;
  assign n27 = n25 & ~n26 ;
  assign n28 = x7 | x8 ;
  assign n29 = x3 & x4 ;
  assign n30 = x3 & ~x4 ;
  assign n31 = ( x4 & ~n29 ) | ( x4 & n30 ) | ( ~n29 & n30 ) ;
  assign n32 = ( x8 & n28 ) | ( x8 & ~n31 ) | ( n28 & ~n31 ) ;
  assign n33 = n27 | n32 ;
  assign n34 = ( n23 & ~n24 ) | ( n23 & n33 ) | ( ~n24 & n33 ) ;
  assign n35 = x1 & x4 ;
  assign n36 = ( x0 & ~x5 ) | ( x0 & n35 ) | ( ~x5 & n35 ) ;
  assign n37 = x0 & n35 ;
  assign n38 = x6 | x8 ;
  assign n39 = x7 | n38 ;
  assign n40 = ~x1 & x5 ;
  assign n41 = ( x2 & n39 ) | ( x2 & ~n40 ) | ( n39 & ~n40 ) ;
  assign n42 = ~n39 & n41 ;
  assign n43 = ( x1 & x2 ) | ( x1 & x5 ) | ( x2 & x5 ) ;
  assign n44 = ( n39 & ~n42 ) | ( n39 & n43 ) | ( ~n42 & n43 ) ;
  assign n45 = ( n36 & ~n37 ) | ( n36 & n44 ) | ( ~n37 & n44 ) ;
  assign n46 = ~n34 & n45 ;
  assign n47 = x9 | x10 ;
  assign n48 = ~n22 & n47 ;
  assign n49 = ( n22 & n46 ) | ( n22 & ~n48 ) | ( n46 & ~n48 ) ;
  assign n50 = ( ~x8 & x10 ) | ( ~x8 & n12 ) | ( x10 & n12 ) ;
  assign n51 = ( ~x8 & n12 ) | ( ~x8 & n14 ) | ( n12 & n14 ) ;
  assign n52 = n50 & ~n51 ;
  assign n53 = ( ~x7 & n18 ) | ( ~x7 & n19 ) | ( n18 & n19 ) ;
  assign n54 = ~x7 & n18 ;
  assign n55 = ( n52 & n53 ) | ( n52 & ~n54 ) | ( n53 & ~n54 ) ;
  assign n56 = x0 & x1 ;
  assign n57 = x3 & x5 ;
  assign n58 = ~x3 & x5 ;
  assign n59 = ( n56 & n57 ) | ( n56 & ~n58 ) | ( n57 & ~n58 ) ;
  assign n60 = x4 | x5 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n42 & ~n61 ;
  assign n63 = ~x8 & n29 ;
  assign n64 = x2 & n63 ;
  assign n65 = ( x6 & n12 ) | ( x6 & n64 ) | ( n12 & n64 ) ;
  assign n66 = n62 | n65 ;
  assign n67 = x4 & x6 ;
  assign n68 = ( ~n39 & n42 ) | ( ~n39 & n59 ) | ( n42 & n59 ) ;
  assign n69 = ( ~x8 & n67 ) | ( ~x8 & n68 ) | ( n67 & n68 ) ;
  assign n70 = ~n66 & n69 ;
  assign n71 = x7 & ~x8 ;
  assign n72 = ( x5 & n29 ) | ( x5 & ~n71 ) | ( n29 & ~n71 ) ;
  assign n73 = ( x5 & n29 ) | ( x5 & n71 ) | ( n29 & n71 ) ;
  assign n74 = ~n72 & n73 ;
  assign n75 = ( x6 & x8 ) | ( x6 & n23 ) | ( x8 & n23 ) ;
  assign n76 = x6 & n23 ;
  assign n77 = ( n74 & n75 ) | ( n74 & ~n76 ) | ( n75 & ~n76 ) ;
  assign n78 = n47 | n77 ;
  assign n79 = n27 & n30 ;
  assign n80 = n39 | n60 ;
  assign n81 = x1 & ~n80 ;
  assign n82 = ( ~n78 & n79 ) | ( ~n78 & n81 ) | ( n79 & n81 ) ;
  assign n83 = n78 | n82 ;
  assign n84 = ~n55 & n83 ;
  assign n85 = ( ~n55 & n70 ) | ( ~n55 & n84 ) | ( n70 & n84 ) ;
  assign n86 = x7 & ~x10 ;
  assign n87 = ~n18 & n86 ;
  assign n88 = ( x7 & x8 ) | ( x7 & n87 ) | ( x8 & n87 ) ;
  assign n89 = ( x10 & n28 ) | ( x10 & ~n88 ) | ( n28 & ~n88 ) ;
  assign n90 = x9 & n89 ;
  assign n91 = ( x8 & n13 ) | ( x8 & n87 ) | ( n13 & n87 ) ;
  assign n92 = n90 | n91 ;
  assign n93 = ( n54 & n63 ) | ( n54 & ~n67 ) | ( n63 & ~n67 ) ;
  assign n94 = ( n23 & ~n77 ) | ( n23 & n93 ) | ( ~n77 & n93 ) ;
  assign n95 = ( n47 & n66 ) | ( n47 & n94 ) | ( n66 & n94 ) ;
  assign n96 = n66 | n94 ;
  assign n97 = ( n92 & ~n95 ) | ( n92 & n96 ) | ( ~n95 & n96 ) ;
  assign n98 = n66 & n94 ;
  assign n99 = x2 & n80 ;
  assign n100 = ( n80 & ~n98 ) | ( n80 & n99 ) | ( ~n98 & n99 ) ;
  assign n101 = x3 | n47 ;
  assign n102 = n100 | n101 ;
  assign n103 = n98 & n102 ;
  assign n104 = ( x4 & ~n23 ) | ( x4 & n38 ) | ( ~n23 & n38 ) ;
  assign n105 = ~n71 & n104 ;
  assign n106 = ( n47 & n103 ) | ( n47 & ~n105 ) | ( n103 & ~n105 ) ;
  assign n107 = ~n103 & n105 ;
  assign n108 = ( ~x8 & n19 ) | ( ~x8 & n54 ) | ( n19 & n54 ) ;
  assign n109 = ( ~n18 & n19 ) | ( ~n18 & n108 ) | ( n19 & n108 ) ;
  assign n110 = ( n106 & n107 ) | ( n106 & ~n109 ) | ( n107 & ~n109 ) ;
  assign n111 = x6 & n98 ;
  assign n112 = x5 | x6 ;
  assign n113 = ~n28 & n112 ;
  assign n114 = n98 | n113 ;
  assign n115 = ~n111 & n114 ;
  assign n116 = x8 | n47 ;
  assign n117 = ( n47 & n103 ) | ( n47 & n116 ) | ( n103 & n116 ) ;
  assign n118 = n115 | n117 ;
  assign n119 = n28 | n47 ;
  assign n120 = n111 | n119 ;
  assign y0 = n49 ;
  assign y1 = n85 ;
  assign y2 = n97 ;
  assign y3 = n102 ;
  assign y4 = n110 ;
  assign y5 = n118 ;
  assign y6 = n120 ;
endmodule
