module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 ;
  assign n257 = x254 | x255 ;
  assign n258 = x253 | n257 ;
  assign n259 = x251 | x252 ;
  assign n260 = x249 | x250 ;
  assign n261 = n259 | n260 ;
  assign n262 = n258 | n261 ;
  assign n263 = x247 | x248 ;
  assign n264 = x245 | x246 ;
  assign n265 = x243 | x244 ;
  assign n266 = n264 | n265 ;
  assign n267 = n263 | n266 ;
  assign n268 = n262 | n267 ;
  assign n269 = x238 | x239 ;
  assign n270 = x237 | n269 ;
  assign n271 = x241 | x242 ;
  assign n272 = x240 | n271 ;
  assign n273 = n270 | n272 ;
  assign n274 = x106 & ~x234 ;
  assign n275 = x107 | n274 ;
  assign n276 = x235 | x236 ;
  assign n277 = n275 & ~n276 ;
  assign n278 = ( x108 & ~x236 ) | ( x108 & n277 ) | ( ~x236 & n277 ) ;
  assign n279 = x109 | n278 ;
  assign n280 = ~n273 & n279 ;
  assign n281 = x110 & ~n269 ;
  assign n282 = ( x111 & ~x239 ) | ( x111 & n281 ) | ( ~x239 & n281 ) ;
  assign n283 = x112 | n282 ;
  assign n284 = ~n272 & n283 ;
  assign n285 = x113 & ~n271 ;
  assign n286 = ( x114 & ~x242 ) | ( x114 & n285 ) | ( ~x242 & n285 ) ;
  assign n287 = x115 | n286 ;
  assign n288 = n284 | n287 ;
  assign n289 = x233 | x234 ;
  assign n290 = n276 | n289 ;
  assign n291 = n273 | n290 ;
  assign n292 = x231 | x232 ;
  assign n293 = x103 & ~n292 ;
  assign n294 = ( x104 & ~x232 ) | ( x104 & n293 ) | ( ~x232 & n293 ) ;
  assign n295 = x105 | n294 ;
  assign n296 = ~n291 & n295 ;
  assign n297 = n288 | n296 ;
  assign n298 = n280 | n297 ;
  assign n299 = x223 | x224 ;
  assign n300 = x225 | n299 ;
  assign n301 = x227 | x228 ;
  assign n302 = x226 | n301 ;
  assign n303 = x229 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = x219 | x220 ;
  assign n306 = x221 | x222 ;
  assign n307 = n305 | n306 ;
  assign n308 = x218 | n307 ;
  assign n309 = n304 | n308 ;
  assign n310 = x216 | x217 ;
  assign n311 = x88 & ~n310 ;
  assign n312 = ( x89 & ~x217 ) | ( x89 & n311 ) | ( ~x217 & n311 ) ;
  assign n313 = x90 | x102 ;
  assign n314 = n312 | n313 ;
  assign n315 = ( x102 & ~n309 ) | ( x102 & n314 ) | ( ~n309 & n314 ) ;
  assign n316 = x99 & ~n301 ;
  assign n317 = ( x100 & ~x228 ) | ( x100 & n316 ) | ( ~x228 & n316 ) ;
  assign n318 = x101 | n317 ;
  assign n319 = x96 & ~x224 ;
  assign n320 = x97 | n319 ;
  assign n321 = ~x225 & n320 ;
  assign n322 = x98 | n321 ;
  assign n323 = x92 & ~x220 ;
  assign n324 = x93 | n323 ;
  assign n325 = x91 & ~n305 ;
  assign n326 = n324 | n325 ;
  assign n327 = ~x94 & x221 ;
  assign n328 = ( x94 & n326 ) | ( x94 & ~n327 ) | ( n326 & ~n327 ) ;
  assign n329 = ~x222 & n328 ;
  assign n330 = x95 | n329 ;
  assign n331 = ~n304 & n330 ;
  assign n332 = ( ~n303 & n322 ) | ( ~n303 & n331 ) | ( n322 & n331 ) ;
  assign n333 = ( ~x229 & n318 ) | ( ~x229 & n332 ) | ( n318 & n332 ) ;
  assign n334 = n315 | n333 ;
  assign n335 = x215 | n310 ;
  assign n336 = n309 | n335 ;
  assign n337 = x86 & ~x214 ;
  assign n338 = x203 | x204 ;
  assign n339 = x202 | n338 ;
  assign n340 = x74 | x77 ;
  assign n341 = ( x77 & ~n339 ) | ( x77 & n340 ) | ( ~n339 & n340 ) ;
  assign n342 = x75 & ~n338 ;
  assign n343 = ( x76 & ~x204 ) | ( x76 & n342 ) | ( ~x204 & n342 ) ;
  assign n344 = n341 | n343 ;
  assign n345 = x207 | x208 ;
  assign n346 = x206 | n345 ;
  assign n347 = x205 | n346 ;
  assign n348 = n344 & ~n347 ;
  assign n349 = x79 | x81 ;
  assign n350 = ( x81 & ~n345 ) | ( x81 & n349 ) | ( ~n345 & n349 ) ;
  assign n351 = x78 & ~n346 ;
  assign n352 = ( x80 & ~x208 ) | ( x80 & n351 ) | ( ~x208 & n351 ) ;
  assign n353 = n350 | n352 ;
  assign n354 = n348 | n353 ;
  assign n355 = x83 & ~x211 ;
  assign n356 = x84 | n355 ;
  assign n357 = x210 | x211 ;
  assign n358 = ~n356 & n357 ;
  assign n359 = ( x82 & n356 ) | ( x82 & ~n358 ) | ( n356 & ~n358 ) ;
  assign n360 = ~x212 & n359 ;
  assign n361 = x85 | n360 ;
  assign n362 = x209 | x212 ;
  assign n363 = n357 | n362 ;
  assign n364 = ~n361 & n363 ;
  assign n365 = ( n354 & n361 ) | ( n354 & ~n364 ) | ( n361 & ~n364 ) ;
  assign n366 = x213 | x214 ;
  assign n367 = ~x87 & n366 ;
  assign n368 = ( x87 & n365 ) | ( x87 & ~n367 ) | ( n365 & ~n367 ) ;
  assign n369 = n337 | n368 ;
  assign n370 = n347 | n363 ;
  assign n371 = x201 | n339 ;
  assign n372 = n366 | n371 ;
  assign n373 = n370 | n372 ;
  assign n374 = x71 & ~x199 ;
  assign n375 = x194 | x195 ;
  assign n376 = x193 | x196 ;
  assign n377 = n375 | n376 ;
  assign n378 = x65 & ~n377 ;
  assign n379 = x198 | x199 ;
  assign n380 = x70 | x72 ;
  assign n381 = ( x72 & ~n379 ) | ( x72 & n380 ) | ( ~n379 & n380 ) ;
  assign n382 = x197 | n379 ;
  assign n383 = ~n381 & n382 ;
  assign n384 = ( n378 & n381 ) | ( n378 & ~n383 ) | ( n381 & ~n383 ) ;
  assign n385 = n374 | n384 ;
  assign n386 = ~x200 & n385 ;
  assign n387 = x73 | n386 ;
  assign n388 = x183 | x184 ;
  assign n389 = x181 | x182 ;
  assign n390 = x180 | n389 ;
  assign n391 = n388 | n390 ;
  assign n392 = x52 | x57 ;
  assign n393 = ( x57 & ~n391 ) | ( x57 & n392 ) | ( ~n391 & n392 ) ;
  assign n394 = x53 & ~n389 ;
  assign n395 = ( x54 & ~x182 ) | ( x54 & n394 ) | ( ~x182 & n394 ) ;
  assign n396 = x55 | n395 ;
  assign n397 = ~n388 & n396 ;
  assign n398 = ( x56 & ~x184 ) | ( x56 & n397 ) | ( ~x184 & n397 ) ;
  assign n399 = n393 | n398 ;
  assign n400 = x58 & ~x186 ;
  assign n401 = x59 | n400 ;
  assign n402 = ~x187 & n401 ;
  assign n403 = x60 | n402 ;
  assign n404 = x185 | x186 ;
  assign n405 = x187 | n404 ;
  assign n406 = ~n403 & n405 ;
  assign n407 = ( n399 & n403 ) | ( n399 & ~n406 ) | ( n403 & ~n406 ) ;
  assign n408 = x67 & ~x195 ;
  assign n409 = x68 | n408 ;
  assign n410 = n375 & ~n409 ;
  assign n411 = ( x66 & n409 ) | ( x66 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = ~x196 & n411 ;
  assign n413 = x69 | n412 ;
  assign n414 = x191 | x192 ;
  assign n415 = x189 | x190 ;
  assign n416 = x61 & ~n415 ;
  assign n417 = ( x62 & ~x190 ) | ( x62 & n416 ) | ( ~x190 & n416 ) ;
  assign n418 = x63 | n417 ;
  assign n419 = ~n414 & n418 ;
  assign n420 = ( x64 & ~x192 ) | ( x64 & n419 ) | ( ~x192 & n419 ) ;
  assign n421 = n377 & ~n413 ;
  assign n422 = ( n413 & n420 ) | ( n413 & ~n421 ) | ( n420 & ~n421 ) ;
  assign n423 = x188 | n415 ;
  assign n424 = n414 | n423 ;
  assign n425 = n377 | n424 ;
  assign n426 = ~n422 & n425 ;
  assign n427 = ( n407 & n422 ) | ( n407 & ~n426 ) | ( n422 & ~n426 ) ;
  assign n428 = n405 | n425 ;
  assign n429 = x179 | n391 ;
  assign n430 = n428 | n429 ;
  assign n431 = x48 & ~x176 ;
  assign n432 = x49 | n431 ;
  assign n433 = x175 | x176 ;
  assign n434 = ~n432 & n433 ;
  assign n435 = x173 | x174 ;
  assign n436 = x45 & ~n435 ;
  assign n437 = x46 & x174 ;
  assign n438 = ( x46 & x47 ) | ( x46 & ~n437 ) | ( x47 & ~n437 ) ;
  assign n439 = n436 | n438 ;
  assign n440 = ( n432 & ~n434 ) | ( n432 & n439 ) | ( ~n434 & n439 ) ;
  assign n441 = ~x177 & n440 ;
  assign n442 = x50 | n441 ;
  assign n443 = x43 & ~x171 ;
  assign n444 = x44 | n443 ;
  assign n445 = x172 | n435 ;
  assign n446 = n433 | n445 ;
  assign n447 = x177 | n446 ;
  assign n448 = ( x178 & n444 ) | ( x178 & n447 ) | ( n444 & n447 ) ;
  assign n449 = n444 & ~n448 ;
  assign n450 = ( ~x178 & n442 ) | ( ~x178 & n449 ) | ( n442 & n449 ) ;
  assign n451 = x51 | n450 ;
  assign n452 = x168 | x169 ;
  assign n453 = x167 | n452 ;
  assign n454 = x166 | n453 ;
  assign n455 = x164 | x165 ;
  assign n456 = x163 | n455 ;
  assign n457 = n454 | n456 ;
  assign n458 = x34 & ~x162 ;
  assign n459 = x35 | n458 ;
  assign n460 = x161 | x162 ;
  assign n461 = n457 | n460 ;
  assign n462 = x159 | x160 ;
  assign n463 = x31 & ~n462 ;
  assign n464 = ( x32 & ~x160 ) | ( x32 & n463 ) | ( ~x160 & n463 ) ;
  assign n465 = x33 | n464 ;
  assign n466 = ~n461 & n465 ;
  assign n467 = ( ~n457 & n459 ) | ( ~n457 & n466 ) | ( n459 & n466 ) ;
  assign n468 = x41 & ~x169 ;
  assign n469 = x36 & ~n455 ;
  assign n470 = ( x37 & ~x165 ) | ( x37 & n469 ) | ( ~x165 & n469 ) ;
  assign n471 = x38 | n470 ;
  assign n472 = ~n454 & n471 ;
  assign n473 = x39 & ~n453 ;
  assign n474 = ( x40 & ~n452 ) | ( x40 & n473 ) | ( ~n452 & n473 ) ;
  assign n475 = x42 | n474 ;
  assign n476 = n472 | n475 ;
  assign n477 = n468 | n476 ;
  assign n478 = n467 | n477 ;
  assign n479 = x171 | n447 ;
  assign n480 = x170 | x178 ;
  assign n481 = n479 | n480 ;
  assign n482 = n430 | n481 ;
  assign n483 = n478 & ~n482 ;
  assign n484 = ( ~n430 & n451 ) | ( ~n430 & n483 ) | ( n451 & n483 ) ;
  assign n485 = n427 | n484 ;
  assign n486 = x200 | n382 ;
  assign n487 = ~n387 & n486 ;
  assign n488 = ( n387 & n485 ) | ( n387 & ~n487 ) | ( n485 & ~n487 ) ;
  assign n489 = x158 | n462 ;
  assign n490 = n461 | n489 ;
  assign n491 = n482 | n486 ;
  assign n492 = n490 | n491 ;
  assign n493 = x155 | x156 ;
  assign n494 = x153 | x154 ;
  assign n495 = x25 & ~n494 ;
  assign n496 = ( x26 & ~x154 ) | ( x26 & n495 ) | ( ~x154 & n495 ) ;
  assign n497 = x27 | n496 ;
  assign n498 = ~n493 & n497 ;
  assign n499 = ( x28 & ~x156 ) | ( x28 & n498 ) | ( ~x156 & n498 ) ;
  assign n500 = x29 | n499 ;
  assign n501 = ~x157 & n500 ;
  assign n502 = x30 | n501 ;
  assign n503 = x157 | n493 ;
  assign n504 = x152 | n494 ;
  assign n505 = n503 | n504 ;
  assign n506 = x22 & ~x150 ;
  assign n507 = x23 | n506 ;
  assign n508 = ~x151 & n507 ;
  assign n509 = x24 | n508 ;
  assign n510 = x145 | x146 ;
  assign n511 = x144 | n510 ;
  assign n512 = x147 | x148 ;
  assign n513 = n511 | n512 ;
  assign n514 = x141 | x142 ;
  assign n515 = x140 | n514 ;
  assign n516 = x12 | x15 ;
  assign n517 = ( x15 & ~n515 ) | ( x15 & n516 ) | ( ~n515 & n516 ) ;
  assign n518 = x13 & ~n514 ;
  assign n519 = ( x14 & ~x142 ) | ( x14 & n518 ) | ( ~x142 & n518 ) ;
  assign n520 = n517 | n519 ;
  assign n521 = x10 & ~x138 ;
  assign n522 = x11 | n521 ;
  assign n523 = x139 | n515 ;
  assign n524 = ~n520 & n523 ;
  assign n525 = ( n520 & n522 ) | ( n520 & ~n524 ) | ( n522 & ~n524 ) ;
  assign n526 = x143 | n525 ;
  assign n527 = ( x16 & ~x143 ) | ( x16 & n526 ) | ( ~x143 & n526 ) ;
  assign n528 = x143 | n523 ;
  assign n529 = x137 | x138 ;
  assign n530 = n528 | n529 ;
  assign n531 = ~n527 & n530 ;
  assign n532 = x135 | x136 ;
  assign n533 = x6 & ~x134 ;
  assign n534 = x7 | n533 ;
  assign n535 = ~n532 & n534 ;
  assign n536 = ( x8 & ~x136 ) | ( x8 & n535 ) | ( ~x136 & n535 ) ;
  assign n537 = x9 | n536 ;
  assign n538 = ( n527 & ~n531 ) | ( n527 & n537 ) | ( ~n531 & n537 ) ;
  assign n539 = ~n513 & n538 ;
  assign n540 = x17 & ~n510 ;
  assign n541 = ( x18 & ~x146 ) | ( x18 & n540 ) | ( ~x146 & n540 ) ;
  assign n542 = x19 | n541 ;
  assign n543 = ~n512 & n542 ;
  assign n544 = ( x20 & ~x148 ) | ( x20 & n543 ) | ( ~x148 & n543 ) ;
  assign n545 = x21 | n544 ;
  assign n546 = n539 | n545 ;
  assign n547 = x149 | x150 ;
  assign n548 = x151 | n547 ;
  assign n549 = ~n509 & n548 ;
  assign n550 = ( n509 & n546 ) | ( n509 & ~n549 ) | ( n546 & ~n549 ) ;
  assign n551 = ~n505 & n550 ;
  assign n552 = n502 | n551 ;
  assign n553 = ~n492 & n552 ;
  assign n554 = n488 | n553 ;
  assign n555 = n513 | n530 ;
  assign n556 = x133 | x134 ;
  assign n557 = n548 | n556 ;
  assign n558 = n532 | n557 ;
  assign n559 = n505 | n558 ;
  assign n560 = n555 | n559 ;
  assign n561 = n492 | n560 ;
  assign n562 = x130 | x131 ;
  assign n563 = x129 | x132 ;
  assign n564 = n562 | n563 ;
  assign n565 = x128 | n268 ;
  assign n566 = n298 & ~n565 ;
  assign n567 = x126 & ~n257 ;
  assign n568 = ( x127 & ~x255 ) | ( x127 & n567 ) | ( ~x255 & n567 ) ;
  assign n569 = x0 | n568 ;
  assign n570 = x118 & ~x246 ;
  assign n571 = x116 & ~x244 ;
  assign n572 = x117 | n571 ;
  assign n573 = ~x119 & n264 ;
  assign n574 = ( x119 & n572 ) | ( x119 & ~n573 ) | ( n572 & ~n573 ) ;
  assign n575 = n570 | n574 ;
  assign n576 = x120 & ~x248 ;
  assign n577 = x121 | n576 ;
  assign n578 = n263 & ~n577 ;
  assign n579 = ( n575 & n577 ) | ( n575 & ~n578 ) | ( n577 & ~n578 ) ;
  assign n580 = x124 & ~x252 ;
  assign n581 = x122 & ~x250 ;
  assign n582 = x123 | n581 ;
  assign n583 = n259 & ~n580 ;
  assign n584 = ( n580 & n582 ) | ( n580 & ~n583 ) | ( n582 & ~n583 ) ;
  assign n585 = x125 | n584 ;
  assign n586 = n261 & ~n585 ;
  assign n587 = ( n579 & n585 ) | ( n579 & ~n586 ) | ( n585 & ~n586 ) ;
  assign n588 = n569 | n587 ;
  assign n589 = ( ~n258 & n569 ) | ( ~n258 & n588 ) | ( n569 & n588 ) ;
  assign n590 = ( ~x128 & n566 ) | ( ~x128 & n589 ) | ( n566 & n589 ) ;
  assign n591 = x1 | n590 ;
  assign n592 = ~n564 & n591 ;
  assign n593 = n291 | n565 ;
  assign n594 = x230 | n292 ;
  assign n595 = n593 | n594 ;
  assign n596 = n564 | n595 ;
  assign n597 = n336 | n596 ;
  assign n598 = n369 & ~n597 ;
  assign n599 = n334 & ~n596 ;
  assign n600 = x3 & ~x131 ;
  assign n601 = x4 | n600 ;
  assign n602 = n562 & ~n601 ;
  assign n603 = ( x2 & n601 ) | ( x2 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = ~x132 & n603 ;
  assign n605 = x5 | n604 ;
  assign n606 = n599 | n605 ;
  assign n607 = n598 | n606 ;
  assign n608 = n592 | n607 ;
  assign n609 = ~n561 & n608 ;
  assign n610 = n554 | n609 ;
  assign n611 = ~n373 & n610 ;
  assign n612 = n369 | n611 ;
  assign n613 = ~n336 & n612 ;
  assign n614 = n334 | n613 ;
  assign n615 = ~x230 & n614 ;
  assign n616 = ~n292 & n615 ;
  assign n617 = n291 & ~n298 ;
  assign n618 = ( n298 & n616 ) | ( n298 & ~n617 ) | ( n616 & ~n617 ) ;
  assign n619 = ~n268 & n618 ;
  assign n620 = x128 & n589 ;
  assign n621 = ( x128 & n619 ) | ( x128 & n620 ) | ( n619 & n620 ) ;
  assign n622 = ~n593 & n616 ;
  assign n623 = n591 | n622 ;
  assign n624 = x129 & n623 ;
  assign n625 = ~x129 & n623 ;
  assign n626 = x2 | n625 ;
  assign n627 = x130 & n626 ;
  assign n628 = ~x130 & n626 ;
  assign n629 = x3 & x131 ;
  assign n630 = ( x131 & n628 ) | ( x131 & n629 ) | ( n628 & n629 ) ;
  assign n631 = ( n601 & ~n602 ) | ( n601 & n626 ) | ( ~n602 & n626 ) ;
  assign n632 = x132 & n631 ;
  assign n633 = n373 | n597 ;
  assign n634 = n554 & ~n633 ;
  assign n635 = n608 | n634 ;
  assign n636 = x133 & n635 ;
  assign n637 = ~x133 & n635 ;
  assign n638 = x6 & x134 ;
  assign n639 = ( x134 & n637 ) | ( x134 & n638 ) | ( n637 & n638 ) ;
  assign n640 = ~x134 & n637 ;
  assign n641 = n534 | n640 ;
  assign n642 = x135 & n641 ;
  assign n643 = ~x135 & n641 ;
  assign n644 = x8 & x136 ;
  assign n645 = ( x136 & n643 ) | ( x136 & n644 ) | ( n643 & n644 ) ;
  assign n646 = ~n532 & n640 ;
  assign n647 = n537 | n646 ;
  assign n648 = x137 & n647 ;
  assign n649 = ~x137 & n647 ;
  assign n650 = x10 & x138 ;
  assign n651 = ( x138 & n649 ) | ( x138 & n650 ) | ( n649 & n650 ) ;
  assign n652 = ~n522 & n529 ;
  assign n653 = ( n522 & n647 ) | ( n522 & ~n652 ) | ( n647 & ~n652 ) ;
  assign n654 = x139 & n653 ;
  assign n655 = ~x139 & n653 ;
  assign n656 = x12 | n655 ;
  assign n657 = x140 & n656 ;
  assign n658 = ~x140 & n656 ;
  assign n659 = x13 | n658 ;
  assign n660 = x141 & n659 ;
  assign n661 = ~x141 & n659 ;
  assign n662 = x14 & x142 ;
  assign n663 = ( x142 & n661 ) | ( x142 & n662 ) | ( n661 & n662 ) ;
  assign n664 = ( n520 & ~n524 ) | ( n520 & n653 ) | ( ~n524 & n653 ) ;
  assign n665 = x143 & n664 ;
  assign n666 = ( ~n531 & n538 ) | ( ~n531 & n647 ) | ( n538 & n647 ) ;
  assign n667 = x144 & n666 ;
  assign n668 = ~x144 & n666 ;
  assign n669 = x17 | n668 ;
  assign n670 = x145 & n669 ;
  assign n671 = ~x145 & n669 ;
  assign n672 = x18 & x146 ;
  assign n673 = ( x146 & n671 ) | ( x146 & n672 ) | ( n671 & n672 ) ;
  assign n674 = n511 & ~n542 ;
  assign n675 = ( n542 & n666 ) | ( n542 & ~n674 ) | ( n666 & ~n674 ) ;
  assign n676 = x147 & n675 ;
  assign n677 = ~x147 & n675 ;
  assign n678 = x20 & x148 ;
  assign n679 = ( x148 & n677 ) | ( x148 & n678 ) | ( n677 & n678 ) ;
  assign n680 = ~n555 & n646 ;
  assign n681 = n546 | n680 ;
  assign n682 = x149 & n681 ;
  assign n683 = ~x149 & n681 ;
  assign n684 = x22 & x150 ;
  assign n685 = ( x150 & n683 ) | ( x150 & n684 ) | ( n683 & n684 ) ;
  assign n686 = ~n547 & n681 ;
  assign n687 = x151 & n507 ;
  assign n688 = ( x151 & n686 ) | ( x151 & n687 ) | ( n686 & n687 ) ;
  assign n689 = ( ~n549 & n550 ) | ( ~n549 & n680 ) | ( n550 & n680 ) ;
  assign n690 = x152 & n689 ;
  assign n691 = ~x152 & n689 ;
  assign n692 = x25 | n691 ;
  assign n693 = x153 & n692 ;
  assign n694 = ~x153 & n692 ;
  assign n695 = x26 & x154 ;
  assign n696 = ( x154 & n694 ) | ( x154 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ~n494 & n691 ;
  assign n698 = n497 | n697 ;
  assign n699 = x155 & n698 ;
  assign n700 = ~x155 & n698 ;
  assign n701 = x28 & x156 ;
  assign n702 = ( x156 & n700 ) | ( x156 & n701 ) | ( n700 & n701 ) ;
  assign n703 = ~n493 & n697 ;
  assign n704 = x157 & n500 ;
  assign n705 = ( x157 & n703 ) | ( x157 & n704 ) | ( n703 & n704 ) ;
  assign n706 = n488 & ~n633 ;
  assign n707 = n608 | n706 ;
  assign n708 = ~n552 & n560 ;
  assign n709 = ( n552 & n707 ) | ( n552 & ~n708 ) | ( n707 & ~n708 ) ;
  assign n710 = x158 & n709 ;
  assign n711 = ~x158 & n709 ;
  assign n712 = x31 | n711 ;
  assign n713 = x159 & n712 ;
  assign n714 = ~x159 & n712 ;
  assign n715 = x32 & x160 ;
  assign n716 = ( x160 & n714 ) | ( x160 & n715 ) | ( n714 & n715 ) ;
  assign n717 = ~n489 & n709 ;
  assign n718 = n465 | n717 ;
  assign n719 = x161 & n718 ;
  assign n720 = ~x161 & n718 ;
  assign n721 = x34 | n720 ;
  assign n722 = x162 & n721 ;
  assign n723 = ~x162 & n721 ;
  assign n724 = x35 | n723 ;
  assign n725 = x163 & n724 ;
  assign n726 = ~x163 & n724 ;
  assign n727 = x36 | n726 ;
  assign n728 = x164 & n727 ;
  assign n729 = ~x164 & n727 ;
  assign n730 = x37 & x165 ;
  assign n731 = ( x165 & n729 ) | ( x165 & n730 ) | ( n729 & n730 ) ;
  assign n732 = n456 & ~n471 ;
  assign n733 = ( n471 & n724 ) | ( n471 & ~n732 ) | ( n724 & ~n732 ) ;
  assign n734 = x166 & n733 ;
  assign n735 = ~x166 & n733 ;
  assign n736 = x39 | n735 ;
  assign n737 = x167 & n736 ;
  assign n738 = ~x167 & n736 ;
  assign n739 = x40 | n738 ;
  assign n740 = x168 & n739 ;
  assign n741 = ~x168 & n739 ;
  assign n742 = x41 & x169 ;
  assign n743 = ( x169 & n741 ) | ( x169 & n742 ) | ( n741 & n742 ) ;
  assign n744 = ~n490 & n709 ;
  assign n745 = n478 | n744 ;
  assign n746 = x170 & n745 ;
  assign n747 = ~x170 & n745 ;
  assign n748 = x43 | n747 ;
  assign n749 = x171 & n748 ;
  assign n750 = ~x171 & n748 ;
  assign n751 = x44 | n750 ;
  assign n752 = x172 & n751 ;
  assign n753 = ~x172 & n751 ;
  assign n754 = x45 | n753 ;
  assign n755 = x173 & n754 ;
  assign n756 = ~x173 & n754 ;
  assign n757 = ( x174 & n437 ) | ( x174 & n756 ) | ( n437 & n756 ) ;
  assign n758 = ~n439 & n445 ;
  assign n759 = ( n439 & n751 ) | ( n439 & ~n758 ) | ( n751 & ~n758 ) ;
  assign n760 = x175 & n759 ;
  assign n761 = ~x175 & n759 ;
  assign n762 = x48 & x176 ;
  assign n763 = ( x176 & n761 ) | ( x176 & n762 ) | ( n761 & n762 ) ;
  assign n764 = ~n440 & n446 ;
  assign n765 = ( n440 & n751 ) | ( n440 & ~n764 ) | ( n751 & ~n764 ) ;
  assign n766 = x177 & n765 ;
  assign n767 = ~n447 & n751 ;
  assign n768 = x178 & n442 ;
  assign n769 = ( x178 & n767 ) | ( x178 & n768 ) | ( n767 & n768 ) ;
  assign n770 = ~n481 & n745 ;
  assign n771 = n451 | n770 ;
  assign n772 = x179 & n771 ;
  assign n773 = ~x179 & n771 ;
  assign n774 = x52 | n773 ;
  assign n775 = x180 & n774 ;
  assign n776 = ~x180 & n774 ;
  assign n777 = x53 | n776 ;
  assign n778 = x181 & n777 ;
  assign n779 = ~x181 & n777 ;
  assign n780 = x54 & x182 ;
  assign n781 = ( x182 & n779 ) | ( x182 & n780 ) | ( n779 & n780 ) ;
  assign n782 = n390 & ~n396 ;
  assign n783 = ( n396 & n774 ) | ( n396 & ~n782 ) | ( n774 & ~n782 ) ;
  assign n784 = x183 & n783 ;
  assign n785 = ~x183 & n783 ;
  assign n786 = x56 & x184 ;
  assign n787 = ( x184 & n785 ) | ( x184 & n786 ) | ( n785 & n786 ) ;
  assign n788 = ~n391 & n773 ;
  assign n789 = n399 | n788 ;
  assign n790 = x185 & n789 ;
  assign n791 = ~x185 & n789 ;
  assign n792 = x58 & x186 ;
  assign n793 = ( x186 & n791 ) | ( x186 & n792 ) | ( n791 & n792 ) ;
  assign n794 = ~n404 & n789 ;
  assign n795 = x187 & n401 ;
  assign n796 = ( x187 & n794 ) | ( x187 & n795 ) | ( n794 & n795 ) ;
  assign n797 = ( ~n406 & n407 ) | ( ~n406 & n788 ) | ( n407 & n788 ) ;
  assign n798 = x188 & n797 ;
  assign n799 = ~x188 & n797 ;
  assign n800 = x61 | n799 ;
  assign n801 = x189 & n800 ;
  assign n802 = ~x189 & n800 ;
  assign n803 = x62 & x190 ;
  assign n804 = ( x190 & n802 ) | ( x190 & n803 ) | ( n802 & n803 ) ;
  assign n805 = ~n418 & n423 ;
  assign n806 = ( n418 & n797 ) | ( n418 & ~n805 ) | ( n797 & ~n805 ) ;
  assign n807 = x191 & n806 ;
  assign n808 = ~x191 & n806 ;
  assign n809 = x64 & x192 ;
  assign n810 = ( x192 & n808 ) | ( x192 & n809 ) | ( n808 & n809 ) ;
  assign n811 = x65 | n420 ;
  assign n812 = n424 & ~n811 ;
  assign n813 = ( n797 & n811 ) | ( n797 & ~n812 ) | ( n811 & ~n812 ) ;
  assign n814 = x193 & n813 ;
  assign n815 = ~x193 & n813 ;
  assign n816 = x66 | n815 ;
  assign n817 = x194 & n816 ;
  assign n818 = ~x194 & n816 ;
  assign n819 = x67 & x195 ;
  assign n820 = ( x195 & n818 ) | ( x195 & n819 ) | ( n818 & n819 ) ;
  assign n821 = ( ~n410 & n411 ) | ( ~n410 & n815 ) | ( n411 & n815 ) ;
  assign n822 = x196 & n821 ;
  assign n823 = n378 | n427 ;
  assign n824 = n428 & ~n823 ;
  assign n825 = ( n788 & n823 ) | ( n788 & ~n824 ) | ( n823 & ~n824 ) ;
  assign n826 = x197 & n825 ;
  assign n827 = ~x197 & n825 ;
  assign n828 = x70 | n827 ;
  assign n829 = x198 & n828 ;
  assign n830 = ~x198 & n828 ;
  assign n831 = x71 & x199 ;
  assign n832 = ( x199 & n830 ) | ( x199 & n831 ) | ( n830 & n831 ) ;
  assign n833 = n382 & ~n385 ;
  assign n834 = ( n385 & n825 ) | ( n385 & ~n833 ) | ( n825 & ~n833 ) ;
  assign n835 = x200 & n834 ;
  assign n836 = x201 & n610 ;
  assign n837 = ~x201 & n610 ;
  assign n838 = x74 | n837 ;
  assign n839 = x202 & n838 ;
  assign n840 = ~x202 & n838 ;
  assign n841 = x75 | n840 ;
  assign n842 = x203 & n841 ;
  assign n843 = ~x203 & n841 ;
  assign n844 = x76 & x204 ;
  assign n845 = ( x204 & n843 ) | ( x204 & n844 ) | ( n843 & n844 ) ;
  assign n846 = ~n339 & n837 ;
  assign n847 = n344 | n846 ;
  assign n848 = x205 & n847 ;
  assign n849 = ~x205 & n847 ;
  assign n850 = x78 | n849 ;
  assign n851 = x206 & n850 ;
  assign n852 = ~x206 & n850 ;
  assign n853 = x79 | n852 ;
  assign n854 = x207 & n853 ;
  assign n855 = ~x207 & n853 ;
  assign n856 = x80 & x208 ;
  assign n857 = ( x208 & n855 ) | ( x208 & n856 ) | ( n855 & n856 ) ;
  assign n858 = ~n347 & n846 ;
  assign n859 = n354 | n858 ;
  assign n860 = x209 & n859 ;
  assign n861 = ~x209 & n859 ;
  assign n862 = x82 | n861 ;
  assign n863 = x210 & n862 ;
  assign n864 = ~x210 & n862 ;
  assign n865 = x83 & x211 ;
  assign n866 = ( x211 & n864 ) | ( x211 & n865 ) | ( n864 & n865 ) ;
  assign n867 = ( ~n358 & n359 ) | ( ~n358 & n861 ) | ( n359 & n861 ) ;
  assign n868 = x212 & n867 ;
  assign n869 = ( ~n364 & n365 ) | ( ~n364 & n858 ) | ( n365 & n858 ) ;
  assign n870 = x213 & n869 ;
  assign n871 = ~x213 & n869 ;
  assign n872 = x86 & x214 ;
  assign n873 = ( x214 & n871 ) | ( x214 & n872 ) | ( n871 & n872 ) ;
  assign n874 = x215 & n612 ;
  assign n875 = ~x215 & n612 ;
  assign n876 = x88 | n875 ;
  assign n877 = x216 & n876 ;
  assign n878 = ~x216 & n876 ;
  assign n879 = x89 | n878 ;
  assign n880 = x217 & n879 ;
  assign n881 = ~x217 & n879 ;
  assign n882 = x90 | n881 ;
  assign n883 = x218 & n882 ;
  assign n884 = ~x218 & n882 ;
  assign n885 = x91 | n884 ;
  assign n886 = x219 & n885 ;
  assign n887 = ~x219 & n885 ;
  assign n888 = x92 & x220 ;
  assign n889 = ( x220 & n887 ) | ( x220 & n888 ) | ( n887 & n888 ) ;
  assign n890 = ~x220 & n887 ;
  assign n891 = n324 | n890 ;
  assign n892 = x221 & n891 ;
  assign n893 = ( ~n327 & n328 ) | ( ~n327 & n890 ) | ( n328 & n890 ) ;
  assign n894 = x222 & n893 ;
  assign n895 = n307 & ~n330 ;
  assign n896 = ( n330 & n884 ) | ( n330 & ~n895 ) | ( n884 & ~n895 ) ;
  assign n897 = x223 & n896 ;
  assign n898 = ~x223 & n896 ;
  assign n899 = x96 & x224 ;
  assign n900 = ( x224 & n898 ) | ( x224 & n899 ) | ( n898 & n899 ) ;
  assign n901 = n299 & ~n320 ;
  assign n902 = ( n320 & n896 ) | ( n320 & ~n901 ) | ( n896 & ~n901 ) ;
  assign n903 = x225 & n902 ;
  assign n904 = n300 & ~n322 ;
  assign n905 = ( n322 & n896 ) | ( n322 & ~n904 ) | ( n896 & ~n904 ) ;
  assign n906 = x226 & n905 ;
  assign n907 = ~x226 & n905 ;
  assign n908 = x99 | n907 ;
  assign n909 = x227 & n908 ;
  assign n910 = ~x227 & n908 ;
  assign n911 = x100 & x228 ;
  assign n912 = ( x228 & n910 ) | ( x228 & n911 ) | ( n910 & n911 ) ;
  assign n913 = n302 & ~n318 ;
  assign n914 = ( n318 & n905 ) | ( n318 & ~n913 ) | ( n905 & ~n913 ) ;
  assign n915 = x229 & n914 ;
  assign n916 = x230 & n614 ;
  assign n917 = x103 | n615 ;
  assign n918 = x231 & n917 ;
  assign n919 = ~x231 & n917 ;
  assign n920 = x104 & x232 ;
  assign n921 = ( x232 & n919 ) | ( x232 & n920 ) | ( n919 & n920 ) ;
  assign n922 = n295 | n616 ;
  assign n923 = x233 & n922 ;
  assign n924 = ~x233 & n922 ;
  assign n925 = x106 & x234 ;
  assign n926 = ( x234 & n924 ) | ( x234 & n925 ) | ( n924 & n925 ) ;
  assign n927 = ~n289 & n922 ;
  assign n928 = n275 | n927 ;
  assign n929 = x235 & n928 ;
  assign n930 = ~x235 & n928 ;
  assign n931 = x108 & x236 ;
  assign n932 = ( x236 & n930 ) | ( x236 & n931 ) | ( n930 & n931 ) ;
  assign n933 = ~n290 & n922 ;
  assign n934 = n279 | n933 ;
  assign n935 = x237 & n934 ;
  assign n936 = ~x237 & n934 ;
  assign n937 = x110 | n936 ;
  assign n938 = x238 & n937 ;
  assign n939 = ~x238 & n937 ;
  assign n940 = x111 & x239 ;
  assign n941 = ( x239 & n939 ) | ( x239 & n940 ) | ( n939 & n940 ) ;
  assign n942 = n270 & ~n283 ;
  assign n943 = ( n283 & n934 ) | ( n283 & ~n942 ) | ( n934 & ~n942 ) ;
  assign n944 = x240 & n943 ;
  assign n945 = ~x240 & n943 ;
  assign n946 = x113 | n945 ;
  assign n947 = x241 & n946 ;
  assign n948 = ~x241 & n946 ;
  assign n949 = x114 & x242 ;
  assign n950 = ( x242 & n948 ) | ( x242 & n949 ) | ( n948 & n949 ) ;
  assign n951 = x243 & n618 ;
  assign n952 = ~x243 & n618 ;
  assign n953 = x116 | n952 ;
  assign n954 = x244 & n953 ;
  assign n955 = ~x244 & n953 ;
  assign n956 = x117 | n955 ;
  assign n957 = x245 & n956 ;
  assign n958 = ~x245 & n956 ;
  assign n959 = x118 & x246 ;
  assign n960 = ( x246 & n958 ) | ( x246 & n959 ) | ( n958 & n959 ) ;
  assign n961 = n266 & ~n575 ;
  assign n962 = ( n575 & n618 ) | ( n575 & ~n961 ) | ( n618 & ~n961 ) ;
  assign n963 = x247 & n962 ;
  assign n964 = ~x247 & n962 ;
  assign n965 = x120 & x248 ;
  assign n966 = ( x248 & n964 ) | ( x248 & n965 ) | ( n964 & n965 ) ;
  assign n967 = n267 & ~n579 ;
  assign n968 = ( n579 & n618 ) | ( n579 & ~n967 ) | ( n618 & ~n967 ) ;
  assign n969 = x249 & n968 ;
  assign n970 = ~x249 & n968 ;
  assign n971 = x122 | n970 ;
  assign n972 = x250 & n971 ;
  assign n973 = ~x250 & n971 ;
  assign n974 = x123 | n973 ;
  assign n975 = x251 & n974 ;
  assign n976 = ~x251 & n974 ;
  assign n977 = x124 & x252 ;
  assign n978 = ( x252 & n976 ) | ( x252 & n977 ) | ( n976 & n977 ) ;
  assign n979 = ( n585 & ~n586 ) | ( n585 & n968 ) | ( ~n586 & n968 ) ;
  assign n980 = x253 & n979 ;
  assign n981 = ~x253 & n979 ;
  assign n982 = x126 | n981 ;
  assign n983 = x254 & n982 ;
  assign n984 = ~x254 & n982 ;
  assign n985 = x127 & x255 ;
  assign n986 = ( x255 & n984 ) | ( x255 & n985 ) | ( n984 & n985 ) ;
  assign n987 = n561 | n633 ;
  assign y0 = n621 ;
  assign y1 = n624 ;
  assign y2 = n627 ;
  assign y3 = n630 ;
  assign y4 = n632 ;
  assign y5 = n636 ;
  assign y6 = n639 ;
  assign y7 = n642 ;
  assign y8 = n645 ;
  assign y9 = n648 ;
  assign y10 = n651 ;
  assign y11 = n654 ;
  assign y12 = n657 ;
  assign y13 = n660 ;
  assign y14 = n663 ;
  assign y15 = n665 ;
  assign y16 = n667 ;
  assign y17 = n670 ;
  assign y18 = n673 ;
  assign y19 = n676 ;
  assign y20 = n679 ;
  assign y21 = n682 ;
  assign y22 = n685 ;
  assign y23 = n688 ;
  assign y24 = n690 ;
  assign y25 = n693 ;
  assign y26 = n696 ;
  assign y27 = n699 ;
  assign y28 = n702 ;
  assign y29 = n705 ;
  assign y30 = n710 ;
  assign y31 = n713 ;
  assign y32 = n716 ;
  assign y33 = n719 ;
  assign y34 = n722 ;
  assign y35 = n725 ;
  assign y36 = n728 ;
  assign y37 = n731 ;
  assign y38 = n734 ;
  assign y39 = n737 ;
  assign y40 = n740 ;
  assign y41 = n743 ;
  assign y42 = n746 ;
  assign y43 = n749 ;
  assign y44 = n752 ;
  assign y45 = n755 ;
  assign y46 = n757 ;
  assign y47 = n760 ;
  assign y48 = n763 ;
  assign y49 = n766 ;
  assign y50 = n769 ;
  assign y51 = n772 ;
  assign y52 = n775 ;
  assign y53 = n778 ;
  assign y54 = n781 ;
  assign y55 = n784 ;
  assign y56 = n787 ;
  assign y57 = n790 ;
  assign y58 = n793 ;
  assign y59 = n796 ;
  assign y60 = n798 ;
  assign y61 = n801 ;
  assign y62 = n804 ;
  assign y63 = n807 ;
  assign y64 = n810 ;
  assign y65 = n814 ;
  assign y66 = n817 ;
  assign y67 = n820 ;
  assign y68 = n822 ;
  assign y69 = n826 ;
  assign y70 = n829 ;
  assign y71 = n832 ;
  assign y72 = n835 ;
  assign y73 = n836 ;
  assign y74 = n839 ;
  assign y75 = n842 ;
  assign y76 = n845 ;
  assign y77 = n848 ;
  assign y78 = n851 ;
  assign y79 = n854 ;
  assign y80 = n857 ;
  assign y81 = n860 ;
  assign y82 = n863 ;
  assign y83 = n866 ;
  assign y84 = n868 ;
  assign y85 = n870 ;
  assign y86 = n873 ;
  assign y87 = n874 ;
  assign y88 = n877 ;
  assign y89 = n880 ;
  assign y90 = n883 ;
  assign y91 = n886 ;
  assign y92 = n889 ;
  assign y93 = n892 ;
  assign y94 = n894 ;
  assign y95 = n897 ;
  assign y96 = n900 ;
  assign y97 = n903 ;
  assign y98 = n906 ;
  assign y99 = n909 ;
  assign y100 = n912 ;
  assign y101 = n915 ;
  assign y102 = n916 ;
  assign y103 = n918 ;
  assign y104 = n921 ;
  assign y105 = n923 ;
  assign y106 = n926 ;
  assign y107 = n929 ;
  assign y108 = n932 ;
  assign y109 = n935 ;
  assign y110 = n938 ;
  assign y111 = n941 ;
  assign y112 = n944 ;
  assign y113 = n947 ;
  assign y114 = n950 ;
  assign y115 = n951 ;
  assign y116 = n954 ;
  assign y117 = n957 ;
  assign y118 = n960 ;
  assign y119 = n963 ;
  assign y120 = n966 ;
  assign y121 = n969 ;
  assign y122 = n972 ;
  assign y123 = n975 ;
  assign y124 = n978 ;
  assign y125 = n980 ;
  assign y126 = n983 ;
  assign y127 = n986 ;
  assign y128 = n987 ;
endmodule
