module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 ;
  assign n136 = x2 & ~x128 ;
  assign n137 = x1 & ~x128 ;
  assign n138 = ( x1 & n136 ) | ( x1 & ~n137 ) | ( n136 & ~n137 ) ;
  assign n139 = x129 & ~n138 ;
  assign n140 = x4 & ~x128 ;
  assign n141 = x3 & ~x128 ;
  assign n142 = ( x3 & n140 ) | ( x3 & ~n141 ) | ( n140 & ~n141 ) ;
  assign n143 = x129 & ~n142 ;
  assign n144 = ( ~n139 & n142 ) | ( ~n139 & n143 ) | ( n142 & n143 ) ;
  assign n145 = x131 & ~n144 ;
  assign n146 = x10 & ~x128 ;
  assign n147 = x9 & ~x128 ;
  assign n148 = ( x9 & n146 ) | ( x9 & ~n147 ) | ( n146 & ~n147 ) ;
  assign n149 = x129 & ~n148 ;
  assign n150 = x12 & ~x128 ;
  assign n151 = x11 & ~x128 ;
  assign n152 = ( x11 & n150 ) | ( x11 & ~n151 ) | ( n150 & ~n151 ) ;
  assign n153 = x129 & ~n152 ;
  assign n154 = ( ~n149 & n152 ) | ( ~n149 & n153 ) | ( n152 & n153 ) ;
  assign n155 = x131 & ~n154 ;
  assign n156 = ( ~n145 & n154 ) | ( ~n145 & n155 ) | ( n154 & n155 ) ;
  assign n157 = ~x130 & n156 ;
  assign n158 = x6 & ~x128 ;
  assign n159 = x5 & ~x128 ;
  assign n160 = ( x5 & n158 ) | ( x5 & ~n159 ) | ( n158 & ~n159 ) ;
  assign n161 = x129 & ~n160 ;
  assign n162 = x8 & ~x128 ;
  assign n163 = x7 & ~x128 ;
  assign n164 = ( x7 & n162 ) | ( x7 & ~n163 ) | ( n162 & ~n163 ) ;
  assign n165 = x129 & ~n164 ;
  assign n166 = ( ~n161 & n164 ) | ( ~n161 & n165 ) | ( n164 & n165 ) ;
  assign n167 = x131 & ~n166 ;
  assign n168 = x14 & ~x128 ;
  assign n169 = x13 & ~x128 ;
  assign n170 = ( x13 & n168 ) | ( x13 & ~n169 ) | ( n168 & ~n169 ) ;
  assign n171 = x129 & ~n170 ;
  assign n172 = x16 & ~x128 ;
  assign n173 = x15 & ~x128 ;
  assign n174 = ( x15 & n172 ) | ( x15 & ~n173 ) | ( n172 & ~n173 ) ;
  assign n175 = x129 & ~n174 ;
  assign n176 = ( ~n171 & n174 ) | ( ~n171 & n175 ) | ( n174 & n175 ) ;
  assign n177 = x131 & ~n176 ;
  assign n178 = ( ~n167 & n176 ) | ( ~n167 & n177 ) | ( n176 & n177 ) ;
  assign n179 = ~x130 & n178 ;
  assign n180 = ( n156 & ~n157 ) | ( n156 & n179 ) | ( ~n157 & n179 ) ;
  assign n181 = x133 & ~n180 ;
  assign n182 = x34 & ~x128 ;
  assign n183 = x33 & ~x128 ;
  assign n184 = ( x33 & n182 ) | ( x33 & ~n183 ) | ( n182 & ~n183 ) ;
  assign n185 = x129 & ~n184 ;
  assign n186 = x36 & ~x128 ;
  assign n187 = x35 & ~x128 ;
  assign n188 = ( x35 & n186 ) | ( x35 & ~n187 ) | ( n186 & ~n187 ) ;
  assign n189 = x129 & ~n188 ;
  assign n190 = ( ~n185 & n188 ) | ( ~n185 & n189 ) | ( n188 & n189 ) ;
  assign n191 = x131 & ~n190 ;
  assign n192 = x42 & ~x128 ;
  assign n193 = x41 & ~x128 ;
  assign n194 = ( x41 & n192 ) | ( x41 & ~n193 ) | ( n192 & ~n193 ) ;
  assign n195 = x129 & ~n194 ;
  assign n196 = x44 & ~x128 ;
  assign n197 = x43 & ~x128 ;
  assign n198 = ( x43 & n196 ) | ( x43 & ~n197 ) | ( n196 & ~n197 ) ;
  assign n199 = x129 & ~n198 ;
  assign n200 = ( ~n195 & n198 ) | ( ~n195 & n199 ) | ( n198 & n199 ) ;
  assign n201 = x131 & ~n200 ;
  assign n202 = ( ~n191 & n200 ) | ( ~n191 & n201 ) | ( n200 & n201 ) ;
  assign n203 = ~x130 & n202 ;
  assign n204 = x38 & ~x128 ;
  assign n205 = x37 & ~x128 ;
  assign n206 = ( x37 & n204 ) | ( x37 & ~n205 ) | ( n204 & ~n205 ) ;
  assign n207 = x129 & ~n206 ;
  assign n208 = x40 & ~x128 ;
  assign n209 = x39 & ~x128 ;
  assign n210 = ( x39 & n208 ) | ( x39 & ~n209 ) | ( n208 & ~n209 ) ;
  assign n211 = x129 & ~n210 ;
  assign n212 = ( ~n207 & n210 ) | ( ~n207 & n211 ) | ( n210 & n211 ) ;
  assign n213 = x131 & ~n212 ;
  assign n214 = x46 & ~x128 ;
  assign n215 = x45 & ~x128 ;
  assign n216 = ( x45 & n214 ) | ( x45 & ~n215 ) | ( n214 & ~n215 ) ;
  assign n217 = x129 & ~n216 ;
  assign n218 = x48 & ~x128 ;
  assign n219 = x47 & ~x128 ;
  assign n220 = ( x47 & n218 ) | ( x47 & ~n219 ) | ( n218 & ~n219 ) ;
  assign n221 = x129 & ~n220 ;
  assign n222 = ( ~n217 & n220 ) | ( ~n217 & n221 ) | ( n220 & n221 ) ;
  assign n223 = x131 & ~n222 ;
  assign n224 = ( ~n213 & n222 ) | ( ~n213 & n223 ) | ( n222 & n223 ) ;
  assign n225 = ~x130 & n224 ;
  assign n226 = ( n202 & ~n203 ) | ( n202 & n225 ) | ( ~n203 & n225 ) ;
  assign n227 = x133 & ~n226 ;
  assign n228 = ( ~n181 & n226 ) | ( ~n181 & n227 ) | ( n226 & n227 ) ;
  assign n229 = ~x132 & n228 ;
  assign n230 = x18 & ~x128 ;
  assign n231 = x17 & ~x128 ;
  assign n232 = ( x17 & n230 ) | ( x17 & ~n231 ) | ( n230 & ~n231 ) ;
  assign n233 = x129 & ~n232 ;
  assign n234 = x20 & ~x128 ;
  assign n235 = x19 & ~x128 ;
  assign n236 = ( x19 & n234 ) | ( x19 & ~n235 ) | ( n234 & ~n235 ) ;
  assign n237 = x129 & ~n236 ;
  assign n238 = ( ~n233 & n236 ) | ( ~n233 & n237 ) | ( n236 & n237 ) ;
  assign n239 = x131 & ~n238 ;
  assign n240 = x26 & ~x128 ;
  assign n241 = x25 & ~x128 ;
  assign n242 = ( x25 & n240 ) | ( x25 & ~n241 ) | ( n240 & ~n241 ) ;
  assign n243 = x129 & ~n242 ;
  assign n244 = x28 & ~x128 ;
  assign n245 = x27 & ~x128 ;
  assign n246 = ( x27 & n244 ) | ( x27 & ~n245 ) | ( n244 & ~n245 ) ;
  assign n247 = x129 & ~n246 ;
  assign n248 = ( ~n243 & n246 ) | ( ~n243 & n247 ) | ( n246 & n247 ) ;
  assign n249 = x131 & ~n248 ;
  assign n250 = ( ~n239 & n248 ) | ( ~n239 & n249 ) | ( n248 & n249 ) ;
  assign n251 = ~x130 & n250 ;
  assign n252 = x22 & ~x128 ;
  assign n253 = x21 & ~x128 ;
  assign n254 = ( x21 & n252 ) | ( x21 & ~n253 ) | ( n252 & ~n253 ) ;
  assign n255 = x129 & ~n254 ;
  assign n256 = x24 & ~x128 ;
  assign n257 = x23 & ~x128 ;
  assign n258 = ( x23 & n256 ) | ( x23 & ~n257 ) | ( n256 & ~n257 ) ;
  assign n259 = x129 & ~n258 ;
  assign n260 = ( ~n255 & n258 ) | ( ~n255 & n259 ) | ( n258 & n259 ) ;
  assign n261 = x131 & ~n260 ;
  assign n262 = x30 & ~x128 ;
  assign n263 = x29 & ~x128 ;
  assign n264 = ( x29 & n262 ) | ( x29 & ~n263 ) | ( n262 & ~n263 ) ;
  assign n265 = x129 & ~n264 ;
  assign n266 = x32 & ~x128 ;
  assign n267 = x31 & ~x128 ;
  assign n268 = ( x31 & n266 ) | ( x31 & ~n267 ) | ( n266 & ~n267 ) ;
  assign n269 = x129 & ~n268 ;
  assign n270 = ( ~n265 & n268 ) | ( ~n265 & n269 ) | ( n268 & n269 ) ;
  assign n271 = x131 & ~n270 ;
  assign n272 = ( ~n261 & n270 ) | ( ~n261 & n271 ) | ( n270 & n271 ) ;
  assign n273 = ~x130 & n272 ;
  assign n274 = ( n250 & ~n251 ) | ( n250 & n273 ) | ( ~n251 & n273 ) ;
  assign n275 = x133 & ~n274 ;
  assign n276 = x50 & ~x128 ;
  assign n277 = x49 & ~x128 ;
  assign n278 = ( x49 & n276 ) | ( x49 & ~n277 ) | ( n276 & ~n277 ) ;
  assign n279 = x129 & ~n278 ;
  assign n280 = x52 & ~x128 ;
  assign n281 = x51 & ~x128 ;
  assign n282 = ( x51 & n280 ) | ( x51 & ~n281 ) | ( n280 & ~n281 ) ;
  assign n283 = x129 & ~n282 ;
  assign n284 = ( ~n279 & n282 ) | ( ~n279 & n283 ) | ( n282 & n283 ) ;
  assign n285 = x131 & ~n284 ;
  assign n286 = x58 & ~x128 ;
  assign n287 = x57 & ~x128 ;
  assign n288 = ( x57 & n286 ) | ( x57 & ~n287 ) | ( n286 & ~n287 ) ;
  assign n289 = x129 & ~n288 ;
  assign n290 = x60 & ~x128 ;
  assign n291 = x59 & ~x128 ;
  assign n292 = ( x59 & n290 ) | ( x59 & ~n291 ) | ( n290 & ~n291 ) ;
  assign n293 = x129 & ~n292 ;
  assign n294 = ( ~n289 & n292 ) | ( ~n289 & n293 ) | ( n292 & n293 ) ;
  assign n295 = x131 & ~n294 ;
  assign n296 = ( ~n285 & n294 ) | ( ~n285 & n295 ) | ( n294 & n295 ) ;
  assign n297 = ~x130 & n296 ;
  assign n298 = x54 & ~x128 ;
  assign n299 = x53 & ~x128 ;
  assign n300 = ( x53 & n298 ) | ( x53 & ~n299 ) | ( n298 & ~n299 ) ;
  assign n301 = x129 & ~n300 ;
  assign n302 = x56 & ~x128 ;
  assign n303 = x55 & ~x128 ;
  assign n304 = ( x55 & n302 ) | ( x55 & ~n303 ) | ( n302 & ~n303 ) ;
  assign n305 = x129 & ~n304 ;
  assign n306 = ( ~n301 & n304 ) | ( ~n301 & n305 ) | ( n304 & n305 ) ;
  assign n307 = x131 & ~n306 ;
  assign n308 = x62 & ~x128 ;
  assign n309 = x61 & ~x128 ;
  assign n310 = ( x61 & n308 ) | ( x61 & ~n309 ) | ( n308 & ~n309 ) ;
  assign n311 = x129 & ~n310 ;
  assign n312 = x64 & ~x128 ;
  assign n313 = x63 & ~x128 ;
  assign n314 = ( x63 & n312 ) | ( x63 & ~n313 ) | ( n312 & ~n313 ) ;
  assign n315 = x129 & ~n314 ;
  assign n316 = ( ~n311 & n314 ) | ( ~n311 & n315 ) | ( n314 & n315 ) ;
  assign n317 = x131 & ~n316 ;
  assign n318 = ( ~n307 & n316 ) | ( ~n307 & n317 ) | ( n316 & n317 ) ;
  assign n319 = ~x130 & n318 ;
  assign n320 = ( n296 & ~n297 ) | ( n296 & n319 ) | ( ~n297 & n319 ) ;
  assign n321 = x133 & ~n320 ;
  assign n322 = ( ~n275 & n320 ) | ( ~n275 & n321 ) | ( n320 & n321 ) ;
  assign n323 = ~x132 & n322 ;
  assign n324 = ( n228 & ~n229 ) | ( n228 & n323 ) | ( ~n229 & n323 ) ;
  assign n325 = x66 & ~x128 ;
  assign n326 = x65 & ~x128 ;
  assign n327 = ( x65 & n325 ) | ( x65 & ~n326 ) | ( n325 & ~n326 ) ;
  assign n328 = x129 & ~n327 ;
  assign n329 = x68 & ~x128 ;
  assign n330 = x67 & ~x128 ;
  assign n331 = ( x67 & n329 ) | ( x67 & ~n330 ) | ( n329 & ~n330 ) ;
  assign n332 = x129 & ~n331 ;
  assign n333 = ( ~n328 & n331 ) | ( ~n328 & n332 ) | ( n331 & n332 ) ;
  assign n334 = x131 & ~n333 ;
  assign n335 = x74 & ~x128 ;
  assign n336 = x73 & ~x128 ;
  assign n337 = ( x73 & n335 ) | ( x73 & ~n336 ) | ( n335 & ~n336 ) ;
  assign n338 = x129 & ~n337 ;
  assign n339 = x76 & ~x128 ;
  assign n340 = x75 & ~x128 ;
  assign n341 = ( x75 & n339 ) | ( x75 & ~n340 ) | ( n339 & ~n340 ) ;
  assign n342 = x129 & ~n341 ;
  assign n343 = ( ~n338 & n341 ) | ( ~n338 & n342 ) | ( n341 & n342 ) ;
  assign n344 = x131 & ~n343 ;
  assign n345 = ( ~n334 & n343 ) | ( ~n334 & n344 ) | ( n343 & n344 ) ;
  assign n346 = ~x130 & n345 ;
  assign n347 = x70 & ~x128 ;
  assign n348 = x69 & ~x128 ;
  assign n349 = ( x69 & n347 ) | ( x69 & ~n348 ) | ( n347 & ~n348 ) ;
  assign n350 = x129 & ~n349 ;
  assign n351 = x72 & ~x128 ;
  assign n352 = x71 & ~x128 ;
  assign n353 = ( x71 & n351 ) | ( x71 & ~n352 ) | ( n351 & ~n352 ) ;
  assign n354 = x129 & ~n353 ;
  assign n355 = ( ~n350 & n353 ) | ( ~n350 & n354 ) | ( n353 & n354 ) ;
  assign n356 = x131 & ~n355 ;
  assign n357 = x78 & ~x128 ;
  assign n358 = x77 & ~x128 ;
  assign n359 = ( x77 & n357 ) | ( x77 & ~n358 ) | ( n357 & ~n358 ) ;
  assign n360 = x129 & ~n359 ;
  assign n361 = x80 & ~x128 ;
  assign n362 = x79 & ~x128 ;
  assign n363 = ( x79 & n361 ) | ( x79 & ~n362 ) | ( n361 & ~n362 ) ;
  assign n364 = x129 & ~n363 ;
  assign n365 = ( ~n360 & n363 ) | ( ~n360 & n364 ) | ( n363 & n364 ) ;
  assign n366 = x131 & ~n365 ;
  assign n367 = ( ~n356 & n365 ) | ( ~n356 & n366 ) | ( n365 & n366 ) ;
  assign n368 = ~x130 & n367 ;
  assign n369 = ( n345 & ~n346 ) | ( n345 & n368 ) | ( ~n346 & n368 ) ;
  assign n370 = x133 & ~n369 ;
  assign n371 = x98 & ~x128 ;
  assign n372 = x97 & ~x128 ;
  assign n373 = ( x97 & n371 ) | ( x97 & ~n372 ) | ( n371 & ~n372 ) ;
  assign n374 = x129 & ~n373 ;
  assign n375 = x100 & ~x128 ;
  assign n376 = x99 & ~x128 ;
  assign n377 = ( x99 & n375 ) | ( x99 & ~n376 ) | ( n375 & ~n376 ) ;
  assign n378 = x129 & ~n377 ;
  assign n379 = ( ~n374 & n377 ) | ( ~n374 & n378 ) | ( n377 & n378 ) ;
  assign n380 = x131 & ~n379 ;
  assign n381 = x106 & ~x128 ;
  assign n382 = x105 & ~x128 ;
  assign n383 = ( x105 & n381 ) | ( x105 & ~n382 ) | ( n381 & ~n382 ) ;
  assign n384 = x129 & ~n383 ;
  assign n385 = x108 & ~x128 ;
  assign n386 = x107 & ~x128 ;
  assign n387 = ( x107 & n385 ) | ( x107 & ~n386 ) | ( n385 & ~n386 ) ;
  assign n388 = x129 & ~n387 ;
  assign n389 = ( ~n384 & n387 ) | ( ~n384 & n388 ) | ( n387 & n388 ) ;
  assign n390 = x131 & ~n389 ;
  assign n391 = ( ~n380 & n389 ) | ( ~n380 & n390 ) | ( n389 & n390 ) ;
  assign n392 = ~x130 & n391 ;
  assign n393 = x102 & ~x128 ;
  assign n394 = x101 & ~x128 ;
  assign n395 = ( x101 & n393 ) | ( x101 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = x129 & ~n395 ;
  assign n397 = x104 & ~x128 ;
  assign n398 = x103 & ~x128 ;
  assign n399 = ( x103 & n397 ) | ( x103 & ~n398 ) | ( n397 & ~n398 ) ;
  assign n400 = x129 & ~n399 ;
  assign n401 = ( ~n396 & n399 ) | ( ~n396 & n400 ) | ( n399 & n400 ) ;
  assign n402 = x131 & ~n401 ;
  assign n403 = x110 & ~x128 ;
  assign n404 = x109 & ~x128 ;
  assign n405 = ( x109 & n403 ) | ( x109 & ~n404 ) | ( n403 & ~n404 ) ;
  assign n406 = x129 & ~n405 ;
  assign n407 = x112 & ~x128 ;
  assign n408 = x111 & ~x128 ;
  assign n409 = ( x111 & n407 ) | ( x111 & ~n408 ) | ( n407 & ~n408 ) ;
  assign n410 = x129 & ~n409 ;
  assign n411 = ( ~n406 & n409 ) | ( ~n406 & n410 ) | ( n409 & n410 ) ;
  assign n412 = x131 & ~n411 ;
  assign n413 = ( ~n402 & n411 ) | ( ~n402 & n412 ) | ( n411 & n412 ) ;
  assign n414 = ~x130 & n413 ;
  assign n415 = ( n391 & ~n392 ) | ( n391 & n414 ) | ( ~n392 & n414 ) ;
  assign n416 = x133 & ~n415 ;
  assign n417 = ( ~n370 & n415 ) | ( ~n370 & n416 ) | ( n415 & n416 ) ;
  assign n418 = ~x132 & n417 ;
  assign n419 = x82 & ~x128 ;
  assign n420 = x81 & ~x128 ;
  assign n421 = ( x81 & n419 ) | ( x81 & ~n420 ) | ( n419 & ~n420 ) ;
  assign n422 = x129 & ~n421 ;
  assign n423 = x84 & ~x128 ;
  assign n424 = x83 & ~x128 ;
  assign n425 = ( x83 & n423 ) | ( x83 & ~n424 ) | ( n423 & ~n424 ) ;
  assign n426 = x129 & ~n425 ;
  assign n427 = ( ~n422 & n425 ) | ( ~n422 & n426 ) | ( n425 & n426 ) ;
  assign n428 = x131 & ~n427 ;
  assign n429 = x90 & ~x128 ;
  assign n430 = x89 & ~x128 ;
  assign n431 = ( x89 & n429 ) | ( x89 & ~n430 ) | ( n429 & ~n430 ) ;
  assign n432 = x129 & ~n431 ;
  assign n433 = x92 & ~x128 ;
  assign n434 = x91 & ~x128 ;
  assign n435 = ( x91 & n433 ) | ( x91 & ~n434 ) | ( n433 & ~n434 ) ;
  assign n436 = x129 & ~n435 ;
  assign n437 = ( ~n432 & n435 ) | ( ~n432 & n436 ) | ( n435 & n436 ) ;
  assign n438 = x131 & ~n437 ;
  assign n439 = ( ~n428 & n437 ) | ( ~n428 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ~x130 & n439 ;
  assign n441 = x86 & ~x128 ;
  assign n442 = x85 & ~x128 ;
  assign n443 = ( x85 & n441 ) | ( x85 & ~n442 ) | ( n441 & ~n442 ) ;
  assign n444 = x129 & ~n443 ;
  assign n445 = x88 & ~x128 ;
  assign n446 = x87 & ~x128 ;
  assign n447 = ( x87 & n445 ) | ( x87 & ~n446 ) | ( n445 & ~n446 ) ;
  assign n448 = x129 & ~n447 ;
  assign n449 = ( ~n444 & n447 ) | ( ~n444 & n448 ) | ( n447 & n448 ) ;
  assign n450 = x131 & ~n449 ;
  assign n451 = x94 & ~x128 ;
  assign n452 = x93 & ~x128 ;
  assign n453 = ( x93 & n451 ) | ( x93 & ~n452 ) | ( n451 & ~n452 ) ;
  assign n454 = x129 & ~n453 ;
  assign n455 = x96 & ~x128 ;
  assign n456 = x95 & ~x128 ;
  assign n457 = ( x95 & n455 ) | ( x95 & ~n456 ) | ( n455 & ~n456 ) ;
  assign n458 = x129 & ~n457 ;
  assign n459 = ( ~n454 & n457 ) | ( ~n454 & n458 ) | ( n457 & n458 ) ;
  assign n460 = x131 & ~n459 ;
  assign n461 = ( ~n450 & n459 ) | ( ~n450 & n460 ) | ( n459 & n460 ) ;
  assign n462 = ~x130 & n461 ;
  assign n463 = ( n439 & ~n440 ) | ( n439 & n462 ) | ( ~n440 & n462 ) ;
  assign n464 = x133 & ~n463 ;
  assign n465 = x118 & ~x128 ;
  assign n466 = x117 & ~x128 ;
  assign n467 = ( x117 & n465 ) | ( x117 & ~n466 ) | ( n465 & ~n466 ) ;
  assign n468 = x129 & ~n467 ;
  assign n469 = x120 & ~x128 ;
  assign n470 = x119 & ~x128 ;
  assign n471 = ( x119 & n469 ) | ( x119 & ~n470 ) | ( n469 & ~n470 ) ;
  assign n472 = x129 & ~n471 ;
  assign n473 = ( ~n468 & n471 ) | ( ~n468 & n472 ) | ( n471 & n472 ) ;
  assign n474 = x131 & ~n473 ;
  assign n475 = x126 & ~x128 ;
  assign n476 = x125 & ~x128 ;
  assign n477 = ( x125 & n475 ) | ( x125 & ~n476 ) | ( n475 & ~n476 ) ;
  assign n478 = x129 & ~n477 ;
  assign n479 = x0 & ~x128 ;
  assign n480 = x127 & ~x128 ;
  assign n481 = ( x127 & n479 ) | ( x127 & ~n480 ) | ( n479 & ~n480 ) ;
  assign n482 = x129 & ~n481 ;
  assign n483 = ( ~n478 & n481 ) | ( ~n478 & n482 ) | ( n481 & n482 ) ;
  assign n484 = x131 & ~n483 ;
  assign n485 = ( ~n474 & n483 ) | ( ~n474 & n484 ) | ( n483 & n484 ) ;
  assign n486 = ~x130 & n485 ;
  assign n487 = x114 & ~x128 ;
  assign n488 = x113 & ~x128 ;
  assign n489 = ( x113 & n487 ) | ( x113 & ~n488 ) | ( n487 & ~n488 ) ;
  assign n490 = x129 & ~n489 ;
  assign n491 = x116 & ~x128 ;
  assign n492 = x115 & ~x128 ;
  assign n493 = ( x115 & n491 ) | ( x115 & ~n492 ) | ( n491 & ~n492 ) ;
  assign n494 = x129 & ~n493 ;
  assign n495 = ( ~n490 & n493 ) | ( ~n490 & n494 ) | ( n493 & n494 ) ;
  assign n496 = x131 & ~n495 ;
  assign n497 = x122 & ~x128 ;
  assign n498 = x121 & ~x128 ;
  assign n499 = ( x121 & n497 ) | ( x121 & ~n498 ) | ( n497 & ~n498 ) ;
  assign n500 = x129 & ~n499 ;
  assign n501 = x124 & ~x128 ;
  assign n502 = x123 & ~x128 ;
  assign n503 = ( x123 & n501 ) | ( x123 & ~n502 ) | ( n501 & ~n502 ) ;
  assign n504 = x129 & ~n503 ;
  assign n505 = ( ~n500 & n503 ) | ( ~n500 & n504 ) | ( n503 & n504 ) ;
  assign n506 = x131 & ~n505 ;
  assign n507 = ( ~n496 & n505 ) | ( ~n496 & n506 ) | ( n505 & n506 ) ;
  assign n508 = x130 & n507 ;
  assign n509 = n486 | n508 ;
  assign n510 = x133 & ~n509 ;
  assign n511 = ( ~n464 & n509 ) | ( ~n464 & n510 ) | ( n509 & n510 ) ;
  assign n512 = ~x132 & n511 ;
  assign n513 = ( n417 & ~n418 ) | ( n417 & n512 ) | ( ~n418 & n512 ) ;
  assign n514 = ~x134 & n324 ;
  assign n515 = x134 & ~n513 ;
  assign n516 = ( x134 & n514 ) | ( x134 & ~n515 ) | ( n514 & ~n515 ) ;
  assign n517 = ( n324 & n513 ) | ( n324 & ~n516 ) | ( n513 & ~n516 ) ;
  assign n518 = ( x4 & ~n140 ) | ( x4 & n159 ) | ( ~n140 & n159 ) ;
  assign n519 = ( x2 & ~n136 ) | ( x2 & n141 ) | ( ~n136 & n141 ) ;
  assign n520 = x129 & ~n519 ;
  assign n521 = x129 & ~n518 ;
  assign n522 = ( n518 & ~n520 ) | ( n518 & n521 ) | ( ~n520 & n521 ) ;
  assign n523 = x131 & ~n522 ;
  assign n524 = ( x12 & ~n150 ) | ( x12 & n169 ) | ( ~n150 & n169 ) ;
  assign n525 = ( x10 & ~n146 ) | ( x10 & n151 ) | ( ~n146 & n151 ) ;
  assign n526 = x129 & ~n525 ;
  assign n527 = x129 & ~n524 ;
  assign n528 = ( n524 & ~n526 ) | ( n524 & n527 ) | ( ~n526 & n527 ) ;
  assign n529 = x131 & ~n528 ;
  assign n530 = ( ~n523 & n528 ) | ( ~n523 & n529 ) | ( n528 & n529 ) ;
  assign n531 = ~x130 & n530 ;
  assign n532 = ( x8 & n147 ) | ( x8 & ~n162 ) | ( n147 & ~n162 ) ;
  assign n533 = ( x6 & ~n158 ) | ( x6 & n163 ) | ( ~n158 & n163 ) ;
  assign n534 = x129 & ~n533 ;
  assign n535 = x129 & ~n532 ;
  assign n536 = ( n532 & ~n534 ) | ( n532 & n535 ) | ( ~n534 & n535 ) ;
  assign n537 = x131 & ~n536 ;
  assign n538 = ( x16 & ~n172 ) | ( x16 & n231 ) | ( ~n172 & n231 ) ;
  assign n539 = ( x14 & ~n168 ) | ( x14 & n173 ) | ( ~n168 & n173 ) ;
  assign n540 = x129 & ~n539 ;
  assign n541 = x129 & ~n538 ;
  assign n542 = ( n538 & ~n540 ) | ( n538 & n541 ) | ( ~n540 & n541 ) ;
  assign n543 = x131 & ~n542 ;
  assign n544 = ( ~n537 & n542 ) | ( ~n537 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ~x130 & n544 ;
  assign n546 = ( n530 & ~n531 ) | ( n530 & n545 ) | ( ~n531 & n545 ) ;
  assign n547 = x133 & ~n546 ;
  assign n548 = ( x36 & ~n186 ) | ( x36 & n205 ) | ( ~n186 & n205 ) ;
  assign n549 = ( x34 & ~n182 ) | ( x34 & n187 ) | ( ~n182 & n187 ) ;
  assign n550 = x129 & ~n549 ;
  assign n551 = x129 & ~n548 ;
  assign n552 = ( n548 & ~n550 ) | ( n548 & n551 ) | ( ~n550 & n551 ) ;
  assign n553 = x131 & ~n552 ;
  assign n554 = ( x44 & ~n196 ) | ( x44 & n215 ) | ( ~n196 & n215 ) ;
  assign n555 = ( x42 & ~n192 ) | ( x42 & n197 ) | ( ~n192 & n197 ) ;
  assign n556 = x129 & ~n555 ;
  assign n557 = x129 & ~n554 ;
  assign n558 = ( n554 & ~n556 ) | ( n554 & n557 ) | ( ~n556 & n557 ) ;
  assign n559 = x131 & ~n558 ;
  assign n560 = ( ~n553 & n558 ) | ( ~n553 & n559 ) | ( n558 & n559 ) ;
  assign n561 = ~x130 & n560 ;
  assign n562 = ( x40 & n193 ) | ( x40 & ~n208 ) | ( n193 & ~n208 ) ;
  assign n563 = ( x38 & ~n204 ) | ( x38 & n209 ) | ( ~n204 & n209 ) ;
  assign n564 = x129 & ~n563 ;
  assign n565 = x129 & ~n562 ;
  assign n566 = ( n562 & ~n564 ) | ( n562 & n565 ) | ( ~n564 & n565 ) ;
  assign n567 = x131 & ~n566 ;
  assign n568 = ( x48 & ~n218 ) | ( x48 & n277 ) | ( ~n218 & n277 ) ;
  assign n569 = ( x46 & ~n214 ) | ( x46 & n219 ) | ( ~n214 & n219 ) ;
  assign n570 = x129 & ~n569 ;
  assign n571 = x129 & ~n568 ;
  assign n572 = ( n568 & ~n570 ) | ( n568 & n571 ) | ( ~n570 & n571 ) ;
  assign n573 = x131 & ~n572 ;
  assign n574 = ( ~n567 & n572 ) | ( ~n567 & n573 ) | ( n572 & n573 ) ;
  assign n575 = ~x130 & n574 ;
  assign n576 = ( n560 & ~n561 ) | ( n560 & n575 ) | ( ~n561 & n575 ) ;
  assign n577 = x133 & ~n576 ;
  assign n578 = ( ~n547 & n576 ) | ( ~n547 & n577 ) | ( n576 & n577 ) ;
  assign n579 = ~x132 & n578 ;
  assign n580 = ( x20 & ~n234 ) | ( x20 & n253 ) | ( ~n234 & n253 ) ;
  assign n581 = ( x18 & ~n230 ) | ( x18 & n235 ) | ( ~n230 & n235 ) ;
  assign n582 = x129 & ~n581 ;
  assign n583 = x129 & ~n580 ;
  assign n584 = ( n580 & ~n582 ) | ( n580 & n583 ) | ( ~n582 & n583 ) ;
  assign n585 = x131 & ~n584 ;
  assign n586 = ( x28 & ~n244 ) | ( x28 & n263 ) | ( ~n244 & n263 ) ;
  assign n587 = ( x26 & ~n240 ) | ( x26 & n245 ) | ( ~n240 & n245 ) ;
  assign n588 = x129 & ~n587 ;
  assign n589 = x129 & ~n586 ;
  assign n590 = ( n586 & ~n588 ) | ( n586 & n589 ) | ( ~n588 & n589 ) ;
  assign n591 = x131 & ~n590 ;
  assign n592 = ( ~n585 & n590 ) | ( ~n585 & n591 ) | ( n590 & n591 ) ;
  assign n593 = ~x130 & n592 ;
  assign n594 = ( x24 & n241 ) | ( x24 & ~n256 ) | ( n241 & ~n256 ) ;
  assign n595 = ( x22 & ~n252 ) | ( x22 & n257 ) | ( ~n252 & n257 ) ;
  assign n596 = x129 & ~n595 ;
  assign n597 = x129 & ~n594 ;
  assign n598 = ( n594 & ~n596 ) | ( n594 & n597 ) | ( ~n596 & n597 ) ;
  assign n599 = x131 & ~n598 ;
  assign n600 = ( x32 & n183 ) | ( x32 & ~n266 ) | ( n183 & ~n266 ) ;
  assign n601 = ( x30 & ~n262 ) | ( x30 & n267 ) | ( ~n262 & n267 ) ;
  assign n602 = x129 & ~n601 ;
  assign n603 = x129 & ~n600 ;
  assign n604 = ( n600 & ~n602 ) | ( n600 & n603 ) | ( ~n602 & n603 ) ;
  assign n605 = x131 & ~n604 ;
  assign n606 = ( ~n599 & n604 ) | ( ~n599 & n605 ) | ( n604 & n605 ) ;
  assign n607 = ~x130 & n606 ;
  assign n608 = ( n592 & ~n593 ) | ( n592 & n607 ) | ( ~n593 & n607 ) ;
  assign n609 = x133 & ~n608 ;
  assign n610 = ( x52 & ~n280 ) | ( x52 & n299 ) | ( ~n280 & n299 ) ;
  assign n611 = ( x50 & ~n276 ) | ( x50 & n281 ) | ( ~n276 & n281 ) ;
  assign n612 = x129 & ~n611 ;
  assign n613 = x129 & ~n610 ;
  assign n614 = ( n610 & ~n612 ) | ( n610 & n613 ) | ( ~n612 & n613 ) ;
  assign n615 = x131 & ~n614 ;
  assign n616 = ( x60 & ~n290 ) | ( x60 & n309 ) | ( ~n290 & n309 ) ;
  assign n617 = ( x58 & ~n286 ) | ( x58 & n291 ) | ( ~n286 & n291 ) ;
  assign n618 = x129 & ~n617 ;
  assign n619 = x129 & ~n616 ;
  assign n620 = ( n616 & ~n618 ) | ( n616 & n619 ) | ( ~n618 & n619 ) ;
  assign n621 = x131 & ~n620 ;
  assign n622 = ( ~n615 & n620 ) | ( ~n615 & n621 ) | ( n620 & n621 ) ;
  assign n623 = ~x130 & n622 ;
  assign n624 = ( x56 & n287 ) | ( x56 & ~n302 ) | ( n287 & ~n302 ) ;
  assign n625 = ( x54 & ~n298 ) | ( x54 & n303 ) | ( ~n298 & n303 ) ;
  assign n626 = x129 & ~n625 ;
  assign n627 = x129 & ~n624 ;
  assign n628 = ( n624 & ~n626 ) | ( n624 & n627 ) | ( ~n626 & n627 ) ;
  assign n629 = x131 & ~n628 ;
  assign n630 = ( x64 & ~n312 ) | ( x64 & n326 ) | ( ~n312 & n326 ) ;
  assign n631 = ( x62 & ~n308 ) | ( x62 & n313 ) | ( ~n308 & n313 ) ;
  assign n632 = x129 & ~n631 ;
  assign n633 = x129 & ~n630 ;
  assign n634 = ( n630 & ~n632 ) | ( n630 & n633 ) | ( ~n632 & n633 ) ;
  assign n635 = x131 & ~n634 ;
  assign n636 = ( ~n629 & n634 ) | ( ~n629 & n635 ) | ( n634 & n635 ) ;
  assign n637 = ~x130 & n636 ;
  assign n638 = ( n622 & ~n623 ) | ( n622 & n637 ) | ( ~n623 & n637 ) ;
  assign n639 = x133 & ~n638 ;
  assign n640 = ( ~n609 & n638 ) | ( ~n609 & n639 ) | ( n638 & n639 ) ;
  assign n641 = ~x132 & n640 ;
  assign n642 = ( n578 & ~n579 ) | ( n578 & n641 ) | ( ~n579 & n641 ) ;
  assign n643 = ( x68 & ~n329 ) | ( x68 & n348 ) | ( ~n329 & n348 ) ;
  assign n644 = ( x66 & ~n325 ) | ( x66 & n330 ) | ( ~n325 & n330 ) ;
  assign n645 = x129 & ~n644 ;
  assign n646 = x129 & ~n643 ;
  assign n647 = ( n643 & ~n645 ) | ( n643 & n646 ) | ( ~n645 & n646 ) ;
  assign n648 = x131 & ~n647 ;
  assign n649 = ( x76 & ~n339 ) | ( x76 & n358 ) | ( ~n339 & n358 ) ;
  assign n650 = ( x74 & ~n335 ) | ( x74 & n340 ) | ( ~n335 & n340 ) ;
  assign n651 = x129 & ~n650 ;
  assign n652 = x129 & ~n649 ;
  assign n653 = ( n649 & ~n651 ) | ( n649 & n652 ) | ( ~n651 & n652 ) ;
  assign n654 = x131 & ~n653 ;
  assign n655 = ( ~n648 & n653 ) | ( ~n648 & n654 ) | ( n653 & n654 ) ;
  assign n656 = ~x130 & n655 ;
  assign n657 = ( x72 & n336 ) | ( x72 & ~n351 ) | ( n336 & ~n351 ) ;
  assign n658 = ( x70 & ~n347 ) | ( x70 & n352 ) | ( ~n347 & n352 ) ;
  assign n659 = x129 & ~n658 ;
  assign n660 = x129 & ~n657 ;
  assign n661 = ( n657 & ~n659 ) | ( n657 & n660 ) | ( ~n659 & n660 ) ;
  assign n662 = x131 & ~n661 ;
  assign n663 = ( x80 & ~n361 ) | ( x80 & n420 ) | ( ~n361 & n420 ) ;
  assign n664 = ( x78 & ~n357 ) | ( x78 & n362 ) | ( ~n357 & n362 ) ;
  assign n665 = x129 & ~n664 ;
  assign n666 = x129 & ~n663 ;
  assign n667 = ( n663 & ~n665 ) | ( n663 & n666 ) | ( ~n665 & n666 ) ;
  assign n668 = x131 & ~n667 ;
  assign n669 = ( ~n662 & n667 ) | ( ~n662 & n668 ) | ( n667 & n668 ) ;
  assign n670 = ~x130 & n669 ;
  assign n671 = ( n655 & ~n656 ) | ( n655 & n670 ) | ( ~n656 & n670 ) ;
  assign n672 = x133 & ~n671 ;
  assign n673 = ( x100 & ~n375 ) | ( x100 & n394 ) | ( ~n375 & n394 ) ;
  assign n674 = ( x98 & ~n371 ) | ( x98 & n376 ) | ( ~n371 & n376 ) ;
  assign n675 = x129 & ~n674 ;
  assign n676 = x129 & ~n673 ;
  assign n677 = ( n673 & ~n675 ) | ( n673 & n676 ) | ( ~n675 & n676 ) ;
  assign n678 = x131 & ~n677 ;
  assign n679 = ( x108 & ~n385 ) | ( x108 & n404 ) | ( ~n385 & n404 ) ;
  assign n680 = ( x106 & ~n381 ) | ( x106 & n386 ) | ( ~n381 & n386 ) ;
  assign n681 = x129 & ~n680 ;
  assign n682 = x129 & ~n679 ;
  assign n683 = ( n679 & ~n681 ) | ( n679 & n682 ) | ( ~n681 & n682 ) ;
  assign n684 = x131 & ~n683 ;
  assign n685 = ( ~n678 & n683 ) | ( ~n678 & n684 ) | ( n683 & n684 ) ;
  assign n686 = ~x130 & n685 ;
  assign n687 = ( x104 & n382 ) | ( x104 & ~n397 ) | ( n382 & ~n397 ) ;
  assign n688 = ( x102 & ~n393 ) | ( x102 & n398 ) | ( ~n393 & n398 ) ;
  assign n689 = x129 & ~n688 ;
  assign n690 = x129 & ~n687 ;
  assign n691 = ( n687 & ~n689 ) | ( n687 & n690 ) | ( ~n689 & n690 ) ;
  assign n692 = x131 & ~n691 ;
  assign n693 = ( x112 & ~n407 ) | ( x112 & n488 ) | ( ~n407 & n488 ) ;
  assign n694 = ( x110 & ~n403 ) | ( x110 & n408 ) | ( ~n403 & n408 ) ;
  assign n695 = x129 & ~n694 ;
  assign n696 = x129 & ~n693 ;
  assign n697 = ( n693 & ~n695 ) | ( n693 & n696 ) | ( ~n695 & n696 ) ;
  assign n698 = x131 & ~n697 ;
  assign n699 = ( ~n692 & n697 ) | ( ~n692 & n698 ) | ( n697 & n698 ) ;
  assign n700 = ~x130 & n699 ;
  assign n701 = ( n685 & ~n686 ) | ( n685 & n700 ) | ( ~n686 & n700 ) ;
  assign n702 = x133 & ~n701 ;
  assign n703 = ( ~n672 & n701 ) | ( ~n672 & n702 ) | ( n701 & n702 ) ;
  assign n704 = ~x132 & n703 ;
  assign n705 = ( x84 & ~n423 ) | ( x84 & n442 ) | ( ~n423 & n442 ) ;
  assign n706 = ( x82 & ~n419 ) | ( x82 & n424 ) | ( ~n419 & n424 ) ;
  assign n707 = x129 & ~n706 ;
  assign n708 = x129 & ~n705 ;
  assign n709 = ( n705 & ~n707 ) | ( n705 & n708 ) | ( ~n707 & n708 ) ;
  assign n710 = x131 & ~n709 ;
  assign n711 = ( x92 & ~n433 ) | ( x92 & n452 ) | ( ~n433 & n452 ) ;
  assign n712 = ( x90 & ~n429 ) | ( x90 & n434 ) | ( ~n429 & n434 ) ;
  assign n713 = x129 & ~n712 ;
  assign n714 = x129 & ~n711 ;
  assign n715 = ( n711 & ~n713 ) | ( n711 & n714 ) | ( ~n713 & n714 ) ;
  assign n716 = x131 & ~n715 ;
  assign n717 = ( ~n710 & n715 ) | ( ~n710 & n716 ) | ( n715 & n716 ) ;
  assign n718 = ~x130 & n717 ;
  assign n719 = ( x88 & n430 ) | ( x88 & ~n445 ) | ( n430 & ~n445 ) ;
  assign n720 = ( x86 & ~n441 ) | ( x86 & n446 ) | ( ~n441 & n446 ) ;
  assign n721 = x129 & ~n720 ;
  assign n722 = x129 & ~n719 ;
  assign n723 = ( n719 & ~n721 ) | ( n719 & n722 ) | ( ~n721 & n722 ) ;
  assign n724 = x131 & ~n723 ;
  assign n725 = ( x96 & n372 ) | ( x96 & ~n455 ) | ( n372 & ~n455 ) ;
  assign n726 = ( x94 & ~n451 ) | ( x94 & n456 ) | ( ~n451 & n456 ) ;
  assign n727 = x129 & ~n726 ;
  assign n728 = x129 & ~n725 ;
  assign n729 = ( n725 & ~n727 ) | ( n725 & n728 ) | ( ~n727 & n728 ) ;
  assign n730 = x131 & ~n729 ;
  assign n731 = ( ~n724 & n729 ) | ( ~n724 & n730 ) | ( n729 & n730 ) ;
  assign n732 = ~x130 & n731 ;
  assign n733 = ( n717 & ~n718 ) | ( n717 & n732 ) | ( ~n718 & n732 ) ;
  assign n734 = x133 & ~n733 ;
  assign n735 = ( x116 & n466 ) | ( x116 & ~n491 ) | ( n466 & ~n491 ) ;
  assign n736 = ( x114 & ~n487 ) | ( x114 & n492 ) | ( ~n487 & n492 ) ;
  assign n737 = x129 & ~n736 ;
  assign n738 = x129 & ~n735 ;
  assign n739 = ( n735 & ~n737 ) | ( n735 & n738 ) | ( ~n737 & n738 ) ;
  assign n740 = x131 & ~n739 ;
  assign n741 = ( x124 & n476 ) | ( x124 & ~n501 ) | ( n476 & ~n501 ) ;
  assign n742 = ( x122 & ~n497 ) | ( x122 & n502 ) | ( ~n497 & n502 ) ;
  assign n743 = x129 & ~n742 ;
  assign n744 = x129 & ~n741 ;
  assign n745 = ( n741 & ~n743 ) | ( n741 & n744 ) | ( ~n743 & n744 ) ;
  assign n746 = x131 & ~n745 ;
  assign n747 = ( ~n740 & n745 ) | ( ~n740 & n746 ) | ( n745 & n746 ) ;
  assign n748 = ~x130 & n747 ;
  assign n749 = ( x120 & ~n469 ) | ( x120 & n498 ) | ( ~n469 & n498 ) ;
  assign n750 = ( x118 & ~n465 ) | ( x118 & n470 ) | ( ~n465 & n470 ) ;
  assign n751 = x129 & ~n750 ;
  assign n752 = x129 & ~n749 ;
  assign n753 = ( n749 & ~n751 ) | ( n749 & n752 ) | ( ~n751 & n752 ) ;
  assign n754 = x131 & ~n753 ;
  assign n755 = ( x0 & n137 ) | ( x0 & ~n479 ) | ( n137 & ~n479 ) ;
  assign n756 = ( x126 & ~n475 ) | ( x126 & n480 ) | ( ~n475 & n480 ) ;
  assign n757 = x129 & ~n756 ;
  assign n758 = x129 & ~n755 ;
  assign n759 = ( n755 & ~n757 ) | ( n755 & n758 ) | ( ~n757 & n758 ) ;
  assign n760 = x131 & ~n759 ;
  assign n761 = ( ~n754 & n759 ) | ( ~n754 & n760 ) | ( n759 & n760 ) ;
  assign n762 = ~x130 & n761 ;
  assign n763 = ( n747 & ~n748 ) | ( n747 & n762 ) | ( ~n748 & n762 ) ;
  assign n764 = x133 & ~n763 ;
  assign n765 = ( ~n734 & n763 ) | ( ~n734 & n764 ) | ( n763 & n764 ) ;
  assign n766 = ~x132 & n765 ;
  assign n767 = ( n703 & ~n704 ) | ( n703 & n766 ) | ( ~n704 & n766 ) ;
  assign n768 = ~x134 & n642 ;
  assign n769 = x134 & ~n767 ;
  assign n770 = ( x134 & n768 ) | ( x134 & ~n769 ) | ( n768 & ~n769 ) ;
  assign n771 = ( n642 & n767 ) | ( n642 & ~n770 ) | ( n767 & ~n770 ) ;
  assign n772 = ( ~n153 & n170 ) | ( ~n153 & n171 ) | ( n170 & n171 ) ;
  assign n773 = ( ~n143 & n160 ) | ( ~n143 & n161 ) | ( n160 & n161 ) ;
  assign n774 = x131 & ~n773 ;
  assign n775 = x131 & ~n772 ;
  assign n776 = ( n772 & ~n774 ) | ( n772 & n775 ) | ( ~n774 & n775 ) ;
  assign n777 = ~x130 & n776 ;
  assign n778 = ( ~n175 & n232 ) | ( ~n175 & n233 ) | ( n232 & n233 ) ;
  assign n779 = ( n148 & n149 ) | ( n148 & ~n165 ) | ( n149 & ~n165 ) ;
  assign n780 = x131 & ~n779 ;
  assign n781 = x131 & ~n778 ;
  assign n782 = ( n778 & ~n780 ) | ( n778 & n781 ) | ( ~n780 & n781 ) ;
  assign n783 = ~x130 & n782 ;
  assign n784 = ( n776 & ~n777 ) | ( n776 & n783 ) | ( ~n777 & n783 ) ;
  assign n785 = x133 & ~n784 ;
  assign n786 = ( ~n199 & n216 ) | ( ~n199 & n217 ) | ( n216 & n217 ) ;
  assign n787 = ( ~n189 & n206 ) | ( ~n189 & n207 ) | ( n206 & n207 ) ;
  assign n788 = x131 & ~n787 ;
  assign n789 = x131 & ~n786 ;
  assign n790 = ( n786 & ~n788 ) | ( n786 & n789 ) | ( ~n788 & n789 ) ;
  assign n791 = ~x130 & n790 ;
  assign n792 = ( ~n221 & n278 ) | ( ~n221 & n279 ) | ( n278 & n279 ) ;
  assign n793 = ( n194 & n195 ) | ( n194 & ~n211 ) | ( n195 & ~n211 ) ;
  assign n794 = x131 & ~n793 ;
  assign n795 = x131 & ~n792 ;
  assign n796 = ( n792 & ~n794 ) | ( n792 & n795 ) | ( ~n794 & n795 ) ;
  assign n797 = ~x130 & n796 ;
  assign n798 = ( n790 & ~n791 ) | ( n790 & n797 ) | ( ~n791 & n797 ) ;
  assign n799 = x133 & ~n798 ;
  assign n800 = ( ~n785 & n798 ) | ( ~n785 & n799 ) | ( n798 & n799 ) ;
  assign n801 = ~x132 & n800 ;
  assign n802 = ( ~n247 & n264 ) | ( ~n247 & n265 ) | ( n264 & n265 ) ;
  assign n803 = ( ~n237 & n254 ) | ( ~n237 & n255 ) | ( n254 & n255 ) ;
  assign n804 = x131 & ~n803 ;
  assign n805 = x131 & ~n802 ;
  assign n806 = ( n802 & ~n804 ) | ( n802 & n805 ) | ( ~n804 & n805 ) ;
  assign n807 = ~x130 & n806 ;
  assign n808 = ( n184 & n185 ) | ( n184 & ~n269 ) | ( n185 & ~n269 ) ;
  assign n809 = ( n242 & n243 ) | ( n242 & ~n259 ) | ( n243 & ~n259 ) ;
  assign n810 = x131 & ~n809 ;
  assign n811 = x131 & ~n808 ;
  assign n812 = ( n808 & ~n810 ) | ( n808 & n811 ) | ( ~n810 & n811 ) ;
  assign n813 = ~x130 & n812 ;
  assign n814 = ( n806 & ~n807 ) | ( n806 & n813 ) | ( ~n807 & n813 ) ;
  assign n815 = x133 & ~n814 ;
  assign n816 = ( ~n293 & n310 ) | ( ~n293 & n311 ) | ( n310 & n311 ) ;
  assign n817 = ( ~n283 & n300 ) | ( ~n283 & n301 ) | ( n300 & n301 ) ;
  assign n818 = x131 & ~n817 ;
  assign n819 = x131 & ~n816 ;
  assign n820 = ( n816 & ~n818 ) | ( n816 & n819 ) | ( ~n818 & n819 ) ;
  assign n821 = ~x130 & n820 ;
  assign n822 = ( ~n315 & n327 ) | ( ~n315 & n328 ) | ( n327 & n328 ) ;
  assign n823 = ( n288 & n289 ) | ( n288 & ~n305 ) | ( n289 & ~n305 ) ;
  assign n824 = x131 & ~n823 ;
  assign n825 = x131 & ~n822 ;
  assign n826 = ( n822 & ~n824 ) | ( n822 & n825 ) | ( ~n824 & n825 ) ;
  assign n827 = ~x130 & n826 ;
  assign n828 = ( n820 & ~n821 ) | ( n820 & n827 ) | ( ~n821 & n827 ) ;
  assign n829 = x133 & ~n828 ;
  assign n830 = ( ~n815 & n828 ) | ( ~n815 & n829 ) | ( n828 & n829 ) ;
  assign n831 = ~x132 & n830 ;
  assign n832 = ( n800 & ~n801 ) | ( n800 & n831 ) | ( ~n801 & n831 ) ;
  assign n833 = ( ~n342 & n359 ) | ( ~n342 & n360 ) | ( n359 & n360 ) ;
  assign n834 = ( ~n332 & n349 ) | ( ~n332 & n350 ) | ( n349 & n350 ) ;
  assign n835 = x131 & ~n834 ;
  assign n836 = x131 & ~n833 ;
  assign n837 = ( n833 & ~n835 ) | ( n833 & n836 ) | ( ~n835 & n836 ) ;
  assign n838 = ~x130 & n837 ;
  assign n839 = ( ~n364 & n421 ) | ( ~n364 & n422 ) | ( n421 & n422 ) ;
  assign n840 = ( n337 & n338 ) | ( n337 & ~n354 ) | ( n338 & ~n354 ) ;
  assign n841 = x131 & ~n840 ;
  assign n842 = x131 & ~n839 ;
  assign n843 = ( n839 & ~n841 ) | ( n839 & n842 ) | ( ~n841 & n842 ) ;
  assign n844 = ~x130 & n843 ;
  assign n845 = ( n837 & ~n838 ) | ( n837 & n844 ) | ( ~n838 & n844 ) ;
  assign n846 = x133 & ~n845 ;
  assign n847 = ( ~n388 & n405 ) | ( ~n388 & n406 ) | ( n405 & n406 ) ;
  assign n848 = ( ~n378 & n395 ) | ( ~n378 & n396 ) | ( n395 & n396 ) ;
  assign n849 = x131 & ~n848 ;
  assign n850 = x131 & ~n847 ;
  assign n851 = ( n847 & ~n849 ) | ( n847 & n850 ) | ( ~n849 & n850 ) ;
  assign n852 = ~x130 & n851 ;
  assign n853 = ( ~n410 & n489 ) | ( ~n410 & n490 ) | ( n489 & n490 ) ;
  assign n854 = ( n383 & n384 ) | ( n383 & ~n400 ) | ( n384 & ~n400 ) ;
  assign n855 = x131 & ~n854 ;
  assign n856 = x131 & ~n853 ;
  assign n857 = ( n853 & ~n855 ) | ( n853 & n856 ) | ( ~n855 & n856 ) ;
  assign n858 = ~x130 & n857 ;
  assign n859 = ( n851 & ~n852 ) | ( n851 & n858 ) | ( ~n852 & n858 ) ;
  assign n860 = x133 & ~n859 ;
  assign n861 = ( ~n846 & n859 ) | ( ~n846 & n860 ) | ( n859 & n860 ) ;
  assign n862 = ~x132 & n861 ;
  assign n863 = ( ~n436 & n453 ) | ( ~n436 & n454 ) | ( n453 & n454 ) ;
  assign n864 = ( ~n426 & n443 ) | ( ~n426 & n444 ) | ( n443 & n444 ) ;
  assign n865 = x131 & ~n864 ;
  assign n866 = x131 & ~n863 ;
  assign n867 = ( n863 & ~n865 ) | ( n863 & n866 ) | ( ~n865 & n866 ) ;
  assign n868 = ~x130 & n867 ;
  assign n869 = ( n373 & n374 ) | ( n373 & ~n458 ) | ( n374 & ~n458 ) ;
  assign n870 = ( n431 & n432 ) | ( n431 & ~n448 ) | ( n432 & ~n448 ) ;
  assign n871 = x131 & ~n870 ;
  assign n872 = x131 & ~n869 ;
  assign n873 = ( n869 & ~n871 ) | ( n869 & n872 ) | ( ~n871 & n872 ) ;
  assign n874 = ~x130 & n873 ;
  assign n875 = ( n867 & ~n868 ) | ( n867 & n874 ) | ( ~n868 & n874 ) ;
  assign n876 = x133 & ~n875 ;
  assign n877 = ( n477 & n478 ) | ( n477 & ~n504 ) | ( n478 & ~n504 ) ;
  assign n878 = ( n467 & n468 ) | ( n467 & ~n494 ) | ( n468 & ~n494 ) ;
  assign n879 = x131 & ~n878 ;
  assign n880 = x131 & ~n877 ;
  assign n881 = ( n877 & ~n879 ) | ( n877 & n880 ) | ( ~n879 & n880 ) ;
  assign n882 = ~x130 & n881 ;
  assign n883 = ( n138 & n139 ) | ( n138 & ~n482 ) | ( n139 & ~n482 ) ;
  assign n884 = ( ~n472 & n499 ) | ( ~n472 & n500 ) | ( n499 & n500 ) ;
  assign n885 = x131 & ~n884 ;
  assign n886 = x131 & ~n883 ;
  assign n887 = ( n883 & ~n885 ) | ( n883 & n886 ) | ( ~n885 & n886 ) ;
  assign n888 = ~x130 & n887 ;
  assign n889 = ( n881 & ~n882 ) | ( n881 & n888 ) | ( ~n882 & n888 ) ;
  assign n890 = x133 & ~n889 ;
  assign n891 = ( ~n876 & n889 ) | ( ~n876 & n890 ) | ( n889 & n890 ) ;
  assign n892 = ~x132 & n891 ;
  assign n893 = ( n861 & ~n862 ) | ( n861 & n892 ) | ( ~n862 & n892 ) ;
  assign n894 = ~x134 & n832 ;
  assign n895 = x134 & ~n893 ;
  assign n896 = ( x134 & n894 ) | ( x134 & ~n895 ) | ( n894 & ~n895 ) ;
  assign n897 = ( n832 & n893 ) | ( n832 & ~n896 ) | ( n893 & ~n896 ) ;
  assign n898 = ( ~n521 & n533 ) | ( ~n521 & n534 ) | ( n533 & n534 ) ;
  assign n899 = x131 & ~n898 ;
  assign n900 = ( ~n527 & n539 ) | ( ~n527 & n540 ) | ( n539 & n540 ) ;
  assign n901 = x131 & ~n900 ;
  assign n902 = ( ~n899 & n900 ) | ( ~n899 & n901 ) | ( n900 & n901 ) ;
  assign n903 = ~x130 & n902 ;
  assign n904 = ( n525 & n526 ) | ( n525 & ~n535 ) | ( n526 & ~n535 ) ;
  assign n905 = x131 & ~n904 ;
  assign n906 = ( ~n541 & n581 ) | ( ~n541 & n582 ) | ( n581 & n582 ) ;
  assign n907 = x131 & ~n906 ;
  assign n908 = ( ~n905 & n906 ) | ( ~n905 & n907 ) | ( n906 & n907 ) ;
  assign n909 = ~x130 & n908 ;
  assign n910 = ( n902 & ~n903 ) | ( n902 & n909 ) | ( ~n903 & n909 ) ;
  assign n911 = x133 & ~n910 ;
  assign n912 = ( ~n551 & n563 ) | ( ~n551 & n564 ) | ( n563 & n564 ) ;
  assign n913 = x131 & ~n912 ;
  assign n914 = ( ~n557 & n569 ) | ( ~n557 & n570 ) | ( n569 & n570 ) ;
  assign n915 = x131 & ~n914 ;
  assign n916 = ( ~n913 & n914 ) | ( ~n913 & n915 ) | ( n914 & n915 ) ;
  assign n917 = ~x130 & n916 ;
  assign n918 = ( n555 & n556 ) | ( n555 & ~n565 ) | ( n556 & ~n565 ) ;
  assign n919 = x131 & ~n918 ;
  assign n920 = ( ~n571 & n611 ) | ( ~n571 & n612 ) | ( n611 & n612 ) ;
  assign n921 = x131 & ~n920 ;
  assign n922 = ( ~n919 & n920 ) | ( ~n919 & n921 ) | ( n920 & n921 ) ;
  assign n923 = ~x130 & n922 ;
  assign n924 = ( n916 & ~n917 ) | ( n916 & n923 ) | ( ~n917 & n923 ) ;
  assign n925 = x133 & ~n924 ;
  assign n926 = ( ~n911 & n924 ) | ( ~n911 & n925 ) | ( n924 & n925 ) ;
  assign n927 = ~x132 & n926 ;
  assign n928 = ( ~n583 & n595 ) | ( ~n583 & n596 ) | ( n595 & n596 ) ;
  assign n929 = x131 & ~n928 ;
  assign n930 = ( ~n589 & n601 ) | ( ~n589 & n602 ) | ( n601 & n602 ) ;
  assign n931 = x131 & ~n930 ;
  assign n932 = ( ~n929 & n930 ) | ( ~n929 & n931 ) | ( n930 & n931 ) ;
  assign n933 = ~x130 & n932 ;
  assign n934 = ( n587 & n588 ) | ( n587 & ~n597 ) | ( n588 & ~n597 ) ;
  assign n935 = x131 & ~n934 ;
  assign n936 = ( n549 & n550 ) | ( n549 & ~n603 ) | ( n550 & ~n603 ) ;
  assign n937 = x131 & ~n936 ;
  assign n938 = ( ~n935 & n936 ) | ( ~n935 & n937 ) | ( n936 & n937 ) ;
  assign n939 = ~x130 & n938 ;
  assign n940 = ( n932 & ~n933 ) | ( n932 & n939 ) | ( ~n933 & n939 ) ;
  assign n941 = x133 & ~n940 ;
  assign n942 = ( ~n613 & n625 ) | ( ~n613 & n626 ) | ( n625 & n626 ) ;
  assign n943 = x131 & ~n942 ;
  assign n944 = ( ~n619 & n631 ) | ( ~n619 & n632 ) | ( n631 & n632 ) ;
  assign n945 = x131 & ~n944 ;
  assign n946 = ( ~n943 & n944 ) | ( ~n943 & n945 ) | ( n944 & n945 ) ;
  assign n947 = ~x130 & n946 ;
  assign n948 = ( n617 & n618 ) | ( n617 & ~n627 ) | ( n618 & ~n627 ) ;
  assign n949 = x131 & ~n948 ;
  assign n950 = ( ~n633 & n644 ) | ( ~n633 & n645 ) | ( n644 & n645 ) ;
  assign n951 = x131 & ~n950 ;
  assign n952 = ( ~n949 & n950 ) | ( ~n949 & n951 ) | ( n950 & n951 ) ;
  assign n953 = ~x130 & n952 ;
  assign n954 = ( n946 & ~n947 ) | ( n946 & n953 ) | ( ~n947 & n953 ) ;
  assign n955 = x133 & ~n954 ;
  assign n956 = ( ~n941 & n954 ) | ( ~n941 & n955 ) | ( n954 & n955 ) ;
  assign n957 = ~x132 & n956 ;
  assign n958 = ( n926 & ~n927 ) | ( n926 & n957 ) | ( ~n927 & n957 ) ;
  assign n959 = ( ~n646 & n658 ) | ( ~n646 & n659 ) | ( n658 & n659 ) ;
  assign n960 = x131 & ~n959 ;
  assign n961 = ( ~n652 & n664 ) | ( ~n652 & n665 ) | ( n664 & n665 ) ;
  assign n962 = x131 & ~n961 ;
  assign n963 = ( ~n960 & n961 ) | ( ~n960 & n962 ) | ( n961 & n962 ) ;
  assign n964 = ~x130 & n963 ;
  assign n965 = ( n650 & n651 ) | ( n650 & ~n660 ) | ( n651 & ~n660 ) ;
  assign n966 = x131 & ~n965 ;
  assign n967 = ( ~n666 & n706 ) | ( ~n666 & n707 ) | ( n706 & n707 ) ;
  assign n968 = x131 & ~n967 ;
  assign n969 = ( ~n966 & n967 ) | ( ~n966 & n968 ) | ( n967 & n968 ) ;
  assign n970 = ~x130 & n969 ;
  assign n971 = ( n963 & ~n964 ) | ( n963 & n970 ) | ( ~n964 & n970 ) ;
  assign n972 = x133 & ~n971 ;
  assign n973 = ( ~n676 & n688 ) | ( ~n676 & n689 ) | ( n688 & n689 ) ;
  assign n974 = x131 & ~n973 ;
  assign n975 = ( ~n682 & n694 ) | ( ~n682 & n695 ) | ( n694 & n695 ) ;
  assign n976 = x131 & ~n975 ;
  assign n977 = ( ~n974 & n975 ) | ( ~n974 & n976 ) | ( n975 & n976 ) ;
  assign n978 = ~x130 & n977 ;
  assign n979 = ( n680 & n681 ) | ( n680 & ~n690 ) | ( n681 & ~n690 ) ;
  assign n980 = x131 & ~n979 ;
  assign n981 = ( ~n696 & n736 ) | ( ~n696 & n737 ) | ( n736 & n737 ) ;
  assign n982 = x131 & ~n981 ;
  assign n983 = ( ~n980 & n981 ) | ( ~n980 & n982 ) | ( n981 & n982 ) ;
  assign n984 = ~x130 & n983 ;
  assign n985 = ( n977 & ~n978 ) | ( n977 & n984 ) | ( ~n978 & n984 ) ;
  assign n986 = x133 & ~n985 ;
  assign n987 = ( ~n972 & n985 ) | ( ~n972 & n986 ) | ( n985 & n986 ) ;
  assign n988 = ~x132 & n987 ;
  assign n989 = ( ~n708 & n720 ) | ( ~n708 & n721 ) | ( n720 & n721 ) ;
  assign n990 = x131 & ~n989 ;
  assign n991 = ( ~n714 & n726 ) | ( ~n714 & n727 ) | ( n726 & n727 ) ;
  assign n992 = x131 & ~n991 ;
  assign n993 = ( ~n990 & n991 ) | ( ~n990 & n992 ) | ( n991 & n992 ) ;
  assign n994 = ~x130 & n993 ;
  assign n995 = ( n712 & n713 ) | ( n712 & ~n722 ) | ( n713 & ~n722 ) ;
  assign n996 = x131 & ~n995 ;
  assign n997 = ( n674 & n675 ) | ( n674 & ~n728 ) | ( n675 & ~n728 ) ;
  assign n998 = x131 & ~n997 ;
  assign n999 = ( ~n996 & n997 ) | ( ~n996 & n998 ) | ( n997 & n998 ) ;
  assign n1000 = ~x130 & n999 ;
  assign n1001 = ( n993 & ~n994 ) | ( n993 & n1000 ) | ( ~n994 & n1000 ) ;
  assign n1002 = x133 & ~n1001 ;
  assign n1003 = ( ~n738 & n750 ) | ( ~n738 & n751 ) | ( n750 & n751 ) ;
  assign n1004 = x131 & ~n1003 ;
  assign n1005 = ( ~n744 & n756 ) | ( ~n744 & n757 ) | ( n756 & n757 ) ;
  assign n1006 = x131 & ~n1005 ;
  assign n1007 = ( ~n1004 & n1005 ) | ( ~n1004 & n1006 ) | ( n1005 & n1006 ) ;
  assign n1008 = ~x130 & n1007 ;
  assign n1009 = ( n742 & n743 ) | ( n742 & ~n752 ) | ( n743 & ~n752 ) ;
  assign n1010 = x131 & ~n1009 ;
  assign n1011 = ( n519 & n520 ) | ( n519 & ~n758 ) | ( n520 & ~n758 ) ;
  assign n1012 = x131 & ~n1011 ;
  assign n1013 = ( ~n1010 & n1011 ) | ( ~n1010 & n1012 ) | ( n1011 & n1012 ) ;
  assign n1014 = ~x130 & n1013 ;
  assign n1015 = ( n1007 & ~n1008 ) | ( n1007 & n1014 ) | ( ~n1008 & n1014 ) ;
  assign n1016 = x133 & ~n1015 ;
  assign n1017 = ( ~n1002 & n1015 ) | ( ~n1002 & n1016 ) | ( n1015 & n1016 ) ;
  assign n1018 = ~x132 & n1017 ;
  assign n1019 = ( n987 & ~n988 ) | ( n987 & n1018 ) | ( ~n988 & n1018 ) ;
  assign n1020 = ~x134 & n958 ;
  assign n1021 = x134 & ~n1019 ;
  assign n1022 = ( x134 & n1020 ) | ( x134 & ~n1021 ) | ( n1020 & ~n1021 ) ;
  assign n1023 = ( n958 & n1019 ) | ( n958 & ~n1022 ) | ( n1019 & ~n1022 ) ;
  assign n1024 = ( ~n155 & n238 ) | ( ~n155 & n239 ) | ( n238 & n239 ) ;
  assign n1025 = ~x130 & n1024 ;
  assign n1026 = ( n178 & ~n179 ) | ( n178 & n1025 ) | ( ~n179 & n1025 ) ;
  assign n1027 = ~x133 & n1026 ;
  assign n1028 = ( ~n201 & n284 ) | ( ~n201 & n285 ) | ( n284 & n285 ) ;
  assign n1029 = ~x130 & n1028 ;
  assign n1030 = ( n224 & ~n225 ) | ( n224 & n1029 ) | ( ~n225 & n1029 ) ;
  assign n1031 = ~x133 & n1030 ;
  assign n1032 = ( n1026 & ~n1027 ) | ( n1026 & n1031 ) | ( ~n1027 & n1031 ) ;
  assign n1033 = x132 & ~n1032 ;
  assign n1034 = ( n190 & n191 ) | ( n190 & ~n249 ) | ( n191 & ~n249 ) ;
  assign n1035 = ~x130 & n1034 ;
  assign n1036 = ( n272 & ~n273 ) | ( n272 & n1035 ) | ( ~n273 & n1035 ) ;
  assign n1037 = ~x133 & n1036 ;
  assign n1038 = ( ~n295 & n333 ) | ( ~n295 & n334 ) | ( n333 & n334 ) ;
  assign n1039 = ~x130 & n1038 ;
  assign n1040 = ( n318 & ~n319 ) | ( n318 & n1039 ) | ( ~n319 & n1039 ) ;
  assign n1041 = ~x133 & n1040 ;
  assign n1042 = ( n1036 & ~n1037 ) | ( n1036 & n1041 ) | ( ~n1037 & n1041 ) ;
  assign n1043 = ~x132 & n1042 ;
  assign n1044 = ( x132 & ~n1033 ) | ( x132 & n1043 ) | ( ~n1033 & n1043 ) ;
  assign n1045 = ( ~n344 & n427 ) | ( ~n344 & n428 ) | ( n427 & n428 ) ;
  assign n1046 = ~x130 & n1045 ;
  assign n1047 = ( n367 & ~n368 ) | ( n367 & n1046 ) | ( ~n368 & n1046 ) ;
  assign n1048 = ~x133 & n1047 ;
  assign n1049 = ( ~n390 & n495 ) | ( ~n390 & n496 ) | ( n495 & n496 ) ;
  assign n1050 = ~x130 & n1049 ;
  assign n1051 = ( n413 & ~n414 ) | ( n413 & n1050 ) | ( ~n414 & n1050 ) ;
  assign n1052 = ~x133 & n1051 ;
  assign n1053 = ( n1047 & ~n1048 ) | ( n1047 & n1052 ) | ( ~n1048 & n1052 ) ;
  assign n1054 = x132 & ~n1053 ;
  assign n1055 = ( n379 & n380 ) | ( n379 & ~n438 ) | ( n380 & ~n438 ) ;
  assign n1056 = ~x130 & n1055 ;
  assign n1057 = ( n461 & ~n462 ) | ( n461 & n1056 ) | ( ~n462 & n1056 ) ;
  assign n1058 = ~x133 & n1057 ;
  assign n1059 = ( n144 & n145 ) | ( n144 & ~n506 ) | ( n145 & ~n506 ) ;
  assign n1060 = ~x130 & n1059 ;
  assign n1061 = ( n485 & ~n486 ) | ( n485 & n1060 ) | ( ~n486 & n1060 ) ;
  assign n1062 = ~x133 & n1061 ;
  assign n1063 = ( n1057 & ~n1058 ) | ( n1057 & n1062 ) | ( ~n1058 & n1062 ) ;
  assign n1064 = ~x132 & n1063 ;
  assign n1065 = ( x132 & ~n1054 ) | ( x132 & n1064 ) | ( ~n1054 & n1064 ) ;
  assign n1066 = ~x134 & n1044 ;
  assign n1067 = x134 & ~n1065 ;
  assign n1068 = ( x134 & n1066 ) | ( x134 & ~n1067 ) | ( n1066 & ~n1067 ) ;
  assign n1069 = ( n1044 & n1065 ) | ( n1044 & ~n1068 ) | ( n1065 & ~n1068 ) ;
  assign n1070 = ( ~n529 & n584 ) | ( ~n529 & n585 ) | ( n584 & n585 ) ;
  assign n1071 = ~x130 & n1070 ;
  assign n1072 = ( n544 & ~n545 ) | ( n544 & n1071 ) | ( ~n545 & n1071 ) ;
  assign n1073 = ~x133 & n1072 ;
  assign n1074 = ( ~n559 & n614 ) | ( ~n559 & n615 ) | ( n614 & n615 ) ;
  assign n1075 = ~x130 & n1074 ;
  assign n1076 = ( n574 & ~n575 ) | ( n574 & n1075 ) | ( ~n575 & n1075 ) ;
  assign n1077 = ~x133 & n1076 ;
  assign n1078 = ( n1072 & ~n1073 ) | ( n1072 & n1077 ) | ( ~n1073 & n1077 ) ;
  assign n1079 = x132 & ~n1078 ;
  assign n1080 = ( n552 & n553 ) | ( n552 & ~n591 ) | ( n553 & ~n591 ) ;
  assign n1081 = ~x130 & n1080 ;
  assign n1082 = ( n606 & ~n607 ) | ( n606 & n1081 ) | ( ~n607 & n1081 ) ;
  assign n1083 = ~x133 & n1082 ;
  assign n1084 = ( ~n621 & n647 ) | ( ~n621 & n648 ) | ( n647 & n648 ) ;
  assign n1085 = ~x130 & n1084 ;
  assign n1086 = ( n636 & ~n637 ) | ( n636 & n1085 ) | ( ~n637 & n1085 ) ;
  assign n1087 = ~x133 & n1086 ;
  assign n1088 = ( n1082 & ~n1083 ) | ( n1082 & n1087 ) | ( ~n1083 & n1087 ) ;
  assign n1089 = ~x132 & n1088 ;
  assign n1090 = ( x132 & ~n1079 ) | ( x132 & n1089 ) | ( ~n1079 & n1089 ) ;
  assign n1091 = ( ~n654 & n709 ) | ( ~n654 & n710 ) | ( n709 & n710 ) ;
  assign n1092 = ~x130 & n1091 ;
  assign n1093 = ( n669 & ~n670 ) | ( n669 & n1092 ) | ( ~n670 & n1092 ) ;
  assign n1094 = ~x133 & n1093 ;
  assign n1095 = ( ~n684 & n739 ) | ( ~n684 & n740 ) | ( n739 & n740 ) ;
  assign n1096 = ~x130 & n1095 ;
  assign n1097 = ( n699 & ~n700 ) | ( n699 & n1096 ) | ( ~n700 & n1096 ) ;
  assign n1098 = ~x133 & n1097 ;
  assign n1099 = ( n1093 & ~n1094 ) | ( n1093 & n1098 ) | ( ~n1094 & n1098 ) ;
  assign n1100 = x132 & ~n1099 ;
  assign n1101 = ( n677 & n678 ) | ( n677 & ~n716 ) | ( n678 & ~n716 ) ;
  assign n1102 = ~x130 & n1101 ;
  assign n1103 = ( n731 & ~n732 ) | ( n731 & n1102 ) | ( ~n732 & n1102 ) ;
  assign n1104 = ~x133 & n1103 ;
  assign n1105 = ( n522 & n523 ) | ( n522 & ~n746 ) | ( n523 & ~n746 ) ;
  assign n1106 = ~x130 & n1105 ;
  assign n1107 = ( n761 & ~n762 ) | ( n761 & n1106 ) | ( ~n762 & n1106 ) ;
  assign n1108 = ~x133 & n1107 ;
  assign n1109 = ( n1103 & ~n1104 ) | ( n1103 & n1108 ) | ( ~n1104 & n1108 ) ;
  assign n1110 = ~x132 & n1109 ;
  assign n1111 = ( x132 & ~n1100 ) | ( x132 & n1110 ) | ( ~n1100 & n1110 ) ;
  assign n1112 = ~x134 & n1090 ;
  assign n1113 = x134 & ~n1111 ;
  assign n1114 = ( x134 & n1112 ) | ( x134 & ~n1113 ) | ( n1112 & ~n1113 ) ;
  assign n1115 = ( n1090 & n1111 ) | ( n1090 & ~n1114 ) | ( n1111 & ~n1114 ) ;
  assign n1116 = ( ~n789 & n817 ) | ( ~n789 & n818 ) | ( n817 & n818 ) ;
  assign n1117 = ~x130 & n1116 ;
  assign n1118 = ( n796 & ~n797 ) | ( n796 & n1117 ) | ( ~n797 & n1117 ) ;
  assign n1119 = x133 & n1118 ;
  assign n1120 = ( ~n775 & n803 ) | ( ~n775 & n804 ) | ( n803 & n804 ) ;
  assign n1121 = ~x130 & n1120 ;
  assign n1122 = ( n782 & ~n783 ) | ( n782 & n1121 ) | ( ~n783 & n1121 ) ;
  assign n1123 = x133 & n1122 ;
  assign n1124 = ( n1118 & ~n1119 ) | ( n1118 & n1123 ) | ( ~n1119 & n1123 ) ;
  assign n1125 = x132 & ~n1124 ;
  assign n1126 = ( ~n819 & n834 ) | ( ~n819 & n835 ) | ( n834 & n835 ) ;
  assign n1127 = ~x130 & n1126 ;
  assign n1128 = ( n826 & ~n827 ) | ( n826 & n1127 ) | ( ~n827 & n1127 ) ;
  assign n1129 = x133 & n1128 ;
  assign n1130 = ( n787 & n788 ) | ( n787 & ~n805 ) | ( n788 & ~n805 ) ;
  assign n1131 = ~x130 & n1130 ;
  assign n1132 = ( n812 & ~n813 ) | ( n812 & n1131 ) | ( ~n813 & n1131 ) ;
  assign n1133 = x133 & n1132 ;
  assign n1134 = ( n1128 & ~n1129 ) | ( n1128 & n1133 ) | ( ~n1129 & n1133 ) ;
  assign n1135 = ~x132 & n1134 ;
  assign n1136 = ( x132 & ~n1125 ) | ( x132 & n1135 ) | ( ~n1125 & n1135 ) ;
  assign n1137 = ( ~n850 & n878 ) | ( ~n850 & n879 ) | ( n878 & n879 ) ;
  assign n1138 = ~x130 & n1137 ;
  assign n1139 = ( n857 & ~n858 ) | ( n857 & n1138 ) | ( ~n858 & n1138 ) ;
  assign n1140 = x133 & n1139 ;
  assign n1141 = ( ~n836 & n864 ) | ( ~n836 & n865 ) | ( n864 & n865 ) ;
  assign n1142 = ~x130 & n1141 ;
  assign n1143 = ( n843 & ~n844 ) | ( n843 & n1142 ) | ( ~n844 & n1142 ) ;
  assign n1144 = x133 & n1143 ;
  assign n1145 = ( n1139 & ~n1140 ) | ( n1139 & n1144 ) | ( ~n1140 & n1144 ) ;
  assign n1146 = x132 & ~n1145 ;
  assign n1147 = ( n773 & n774 ) | ( n773 & ~n880 ) | ( n774 & ~n880 ) ;
  assign n1148 = ~x130 & n1147 ;
  assign n1149 = ( n887 & ~n888 ) | ( n887 & n1148 ) | ( ~n888 & n1148 ) ;
  assign n1150 = x133 & n1149 ;
  assign n1151 = ( n848 & n849 ) | ( n848 & ~n866 ) | ( n849 & ~n866 ) ;
  assign n1152 = ~x130 & n1151 ;
  assign n1153 = ( n873 & ~n874 ) | ( n873 & n1152 ) | ( ~n874 & n1152 ) ;
  assign n1154 = x133 & n1153 ;
  assign n1155 = ( n1149 & ~n1150 ) | ( n1149 & n1154 ) | ( ~n1150 & n1154 ) ;
  assign n1156 = ~x132 & n1155 ;
  assign n1157 = ( x132 & ~n1146 ) | ( x132 & n1156 ) | ( ~n1146 & n1156 ) ;
  assign n1158 = ~x134 & n1136 ;
  assign n1159 = x134 & ~n1157 ;
  assign n1160 = ( x134 & n1158 ) | ( x134 & ~n1159 ) | ( n1158 & ~n1159 ) ;
  assign n1161 = ( n1136 & n1157 ) | ( n1136 & ~n1160 ) | ( n1157 & ~n1160 ) ;
  assign n1162 = ( ~n915 & n942 ) | ( ~n915 & n943 ) | ( n942 & n943 ) ;
  assign n1163 = ~x130 & n1162 ;
  assign n1164 = ( n922 & ~n923 ) | ( n922 & n1163 ) | ( ~n923 & n1163 ) ;
  assign n1165 = x133 & n1164 ;
  assign n1166 = ( ~n901 & n928 ) | ( ~n901 & n929 ) | ( n928 & n929 ) ;
  assign n1167 = ~x130 & n1166 ;
  assign n1168 = ( n908 & ~n909 ) | ( n908 & n1167 ) | ( ~n909 & n1167 ) ;
  assign n1169 = x133 & n1168 ;
  assign n1170 = ( n1164 & ~n1165 ) | ( n1164 & n1169 ) | ( ~n1165 & n1169 ) ;
  assign n1171 = x132 & ~n1170 ;
  assign n1172 = ( ~n945 & n959 ) | ( ~n945 & n960 ) | ( n959 & n960 ) ;
  assign n1173 = ~x130 & n1172 ;
  assign n1174 = ( n952 & ~n953 ) | ( n952 & n1173 ) | ( ~n953 & n1173 ) ;
  assign n1175 = x133 & n1174 ;
  assign n1176 = ( n912 & n913 ) | ( n912 & ~n931 ) | ( n913 & ~n931 ) ;
  assign n1177 = ~x130 & n1176 ;
  assign n1178 = ( n938 & ~n939 ) | ( n938 & n1177 ) | ( ~n939 & n1177 ) ;
  assign n1179 = x133 & n1178 ;
  assign n1180 = ( n1174 & ~n1175 ) | ( n1174 & n1179 ) | ( ~n1175 & n1179 ) ;
  assign n1181 = ~x132 & n1180 ;
  assign n1182 = ( x132 & ~n1171 ) | ( x132 & n1181 ) | ( ~n1171 & n1181 ) ;
  assign n1183 = ( ~n976 & n1003 ) | ( ~n976 & n1004 ) | ( n1003 & n1004 ) ;
  assign n1184 = ~x130 & n1183 ;
  assign n1185 = ( n983 & ~n984 ) | ( n983 & n1184 ) | ( ~n984 & n1184 ) ;
  assign n1186 = x133 & n1185 ;
  assign n1187 = ( ~n962 & n989 ) | ( ~n962 & n990 ) | ( n989 & n990 ) ;
  assign n1188 = ~x130 & n1187 ;
  assign n1189 = ( n969 & ~n970 ) | ( n969 & n1188 ) | ( ~n970 & n1188 ) ;
  assign n1190 = x133 & n1189 ;
  assign n1191 = ( n1185 & ~n1186 ) | ( n1185 & n1190 ) | ( ~n1186 & n1190 ) ;
  assign n1192 = x132 & ~n1191 ;
  assign n1193 = ( n898 & n899 ) | ( n898 & ~n1006 ) | ( n899 & ~n1006 ) ;
  assign n1194 = ~x130 & n1193 ;
  assign n1195 = ( n1013 & ~n1014 ) | ( n1013 & n1194 ) | ( ~n1014 & n1194 ) ;
  assign n1196 = x133 & n1195 ;
  assign n1197 = ( n973 & n974 ) | ( n973 & ~n992 ) | ( n974 & ~n992 ) ;
  assign n1198 = ~x130 & n1197 ;
  assign n1199 = ( n999 & ~n1000 ) | ( n999 & n1198 ) | ( ~n1000 & n1198 ) ;
  assign n1200 = x133 & n1199 ;
  assign n1201 = ( n1195 & ~n1196 ) | ( n1195 & n1200 ) | ( ~n1196 & n1200 ) ;
  assign n1202 = ~x132 & n1201 ;
  assign n1203 = ( x132 & ~n1192 ) | ( x132 & n1202 ) | ( ~n1192 & n1202 ) ;
  assign n1204 = ~x134 & n1182 ;
  assign n1205 = x134 & ~n1203 ;
  assign n1206 = ( x134 & n1204 ) | ( x134 & ~n1205 ) | ( n1204 & ~n1205 ) ;
  assign n1207 = ( n1182 & n1203 ) | ( n1182 & ~n1206 ) | ( n1203 & ~n1206 ) ;
  assign n1208 = ( ~n177 & n260 ) | ( ~n177 & n261 ) | ( n260 & n261 ) ;
  assign n1209 = ~x130 & n1208 ;
  assign n1210 = ( n1024 & ~n1025 ) | ( n1024 & n1209 ) | ( ~n1025 & n1209 ) ;
  assign n1211 = x133 & ~n1210 ;
  assign n1212 = ( ~n223 & n306 ) | ( ~n223 & n307 ) | ( n306 & n307 ) ;
  assign n1213 = ~x130 & n1212 ;
  assign n1214 = ( n1028 & ~n1029 ) | ( n1028 & n1213 ) | ( ~n1029 & n1213 ) ;
  assign n1215 = x133 & ~n1214 ;
  assign n1216 = ( ~n1211 & n1214 ) | ( ~n1211 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1217 = ~x132 & n1216 ;
  assign n1218 = ( n212 & n213 ) | ( n212 & ~n271 ) | ( n213 & ~n271 ) ;
  assign n1219 = ~x130 & n1218 ;
  assign n1220 = ( n1034 & ~n1035 ) | ( n1034 & n1219 ) | ( ~n1035 & n1219 ) ;
  assign n1221 = x133 & ~n1220 ;
  assign n1222 = ( ~n317 & n355 ) | ( ~n317 & n356 ) | ( n355 & n356 ) ;
  assign n1223 = ~x130 & n1222 ;
  assign n1224 = ( n1038 & ~n1039 ) | ( n1038 & n1223 ) | ( ~n1039 & n1223 ) ;
  assign n1225 = x133 & ~n1224 ;
  assign n1226 = ( ~n1221 & n1224 ) | ( ~n1221 & n1225 ) | ( n1224 & n1225 ) ;
  assign n1227 = ~x132 & n1226 ;
  assign n1228 = ( n1216 & ~n1217 ) | ( n1216 & n1227 ) | ( ~n1217 & n1227 ) ;
  assign n1229 = ( ~n366 & n449 ) | ( ~n366 & n450 ) | ( n449 & n450 ) ;
  assign n1230 = ~x130 & n1229 ;
  assign n1231 = ( n1045 & ~n1046 ) | ( n1045 & n1230 ) | ( ~n1046 & n1230 ) ;
  assign n1232 = x133 & ~n1231 ;
  assign n1233 = ( ~n412 & n473 ) | ( ~n412 & n474 ) | ( n473 & n474 ) ;
  assign n1234 = ~x130 & n1233 ;
  assign n1235 = ( n1049 & ~n1050 ) | ( n1049 & n1234 ) | ( ~n1050 & n1234 ) ;
  assign n1236 = x133 & ~n1235 ;
  assign n1237 = ( ~n1232 & n1235 ) | ( ~n1232 & n1236 ) | ( n1235 & n1236 ) ;
  assign n1238 = ~x132 & n1237 ;
  assign n1239 = ( n401 & n402 ) | ( n401 & ~n460 ) | ( n402 & ~n460 ) ;
  assign n1240 = ~x130 & n1239 ;
  assign n1241 = ( n1055 & ~n1056 ) | ( n1055 & n1240 ) | ( ~n1056 & n1240 ) ;
  assign n1242 = x133 & ~n1241 ;
  assign n1243 = ( n166 & n167 ) | ( n166 & ~n484 ) | ( n167 & ~n484 ) ;
  assign n1244 = ~x130 & n1243 ;
  assign n1245 = ( n1059 & ~n1060 ) | ( n1059 & n1244 ) | ( ~n1060 & n1244 ) ;
  assign n1246 = x133 & ~n1245 ;
  assign n1247 = ( ~n1242 & n1245 ) | ( ~n1242 & n1246 ) | ( n1245 & n1246 ) ;
  assign n1248 = ~x132 & n1247 ;
  assign n1249 = ( n1237 & ~n1238 ) | ( n1237 & n1248 ) | ( ~n1238 & n1248 ) ;
  assign n1250 = ~x134 & n1228 ;
  assign n1251 = x134 & ~n1249 ;
  assign n1252 = ( x134 & n1250 ) | ( x134 & ~n1251 ) | ( n1250 & ~n1251 ) ;
  assign n1253 = ( n1228 & n1249 ) | ( n1228 & ~n1252 ) | ( n1249 & ~n1252 ) ;
  assign n1254 = ( ~n543 & n598 ) | ( ~n543 & n599 ) | ( n598 & n599 ) ;
  assign n1255 = ~x130 & n1254 ;
  assign n1256 = ( n1070 & ~n1071 ) | ( n1070 & n1255 ) | ( ~n1071 & n1255 ) ;
  assign n1257 = x133 & ~n1256 ;
  assign n1258 = ( ~n573 & n628 ) | ( ~n573 & n629 ) | ( n628 & n629 ) ;
  assign n1259 = ~x130 & n1258 ;
  assign n1260 = ( n1074 & ~n1075 ) | ( n1074 & n1259 ) | ( ~n1075 & n1259 ) ;
  assign n1261 = x133 & ~n1260 ;
  assign n1262 = ( ~n1257 & n1260 ) | ( ~n1257 & n1261 ) | ( n1260 & n1261 ) ;
  assign n1263 = ~x132 & n1262 ;
  assign n1264 = ( n566 & n567 ) | ( n566 & ~n605 ) | ( n567 & ~n605 ) ;
  assign n1265 = ~x130 & n1264 ;
  assign n1266 = ( n1080 & ~n1081 ) | ( n1080 & n1265 ) | ( ~n1081 & n1265 ) ;
  assign n1267 = x133 & ~n1266 ;
  assign n1268 = ( ~n635 & n661 ) | ( ~n635 & n662 ) | ( n661 & n662 ) ;
  assign n1269 = ~x130 & n1268 ;
  assign n1270 = ( n1084 & ~n1085 ) | ( n1084 & n1269 ) | ( ~n1085 & n1269 ) ;
  assign n1271 = x133 & ~n1270 ;
  assign n1272 = ( ~n1267 & n1270 ) | ( ~n1267 & n1271 ) | ( n1270 & n1271 ) ;
  assign n1273 = ~x132 & n1272 ;
  assign n1274 = ( n1262 & ~n1263 ) | ( n1262 & n1273 ) | ( ~n1263 & n1273 ) ;
  assign n1275 = ( ~n668 & n723 ) | ( ~n668 & n724 ) | ( n723 & n724 ) ;
  assign n1276 = ~x130 & n1275 ;
  assign n1277 = ( n1091 & ~n1092 ) | ( n1091 & n1276 ) | ( ~n1092 & n1276 ) ;
  assign n1278 = x133 & ~n1277 ;
  assign n1279 = ( ~n698 & n753 ) | ( ~n698 & n754 ) | ( n753 & n754 ) ;
  assign n1280 = ~x130 & n1279 ;
  assign n1281 = ( n1095 & ~n1096 ) | ( n1095 & n1280 ) | ( ~n1096 & n1280 ) ;
  assign n1282 = x133 & ~n1281 ;
  assign n1283 = ( ~n1278 & n1281 ) | ( ~n1278 & n1282 ) | ( n1281 & n1282 ) ;
  assign n1284 = ~x132 & n1283 ;
  assign n1285 = ( n691 & n692 ) | ( n691 & ~n730 ) | ( n692 & ~n730 ) ;
  assign n1286 = ~x130 & n1285 ;
  assign n1287 = ( n1101 & ~n1102 ) | ( n1101 & n1286 ) | ( ~n1102 & n1286 ) ;
  assign n1288 = x133 & ~n1287 ;
  assign n1289 = ( n536 & n537 ) | ( n536 & ~n760 ) | ( n537 & ~n760 ) ;
  assign n1290 = ~x130 & n1289 ;
  assign n1291 = ( n1105 & ~n1106 ) | ( n1105 & n1290 ) | ( ~n1106 & n1290 ) ;
  assign n1292 = x133 & ~n1291 ;
  assign n1293 = ( ~n1288 & n1291 ) | ( ~n1288 & n1292 ) | ( n1291 & n1292 ) ;
  assign n1294 = ~x132 & n1293 ;
  assign n1295 = ( n1283 & ~n1284 ) | ( n1283 & n1294 ) | ( ~n1284 & n1294 ) ;
  assign n1296 = ~x134 & n1274 ;
  assign n1297 = x134 & ~n1295 ;
  assign n1298 = ( x134 & n1296 ) | ( x134 & ~n1297 ) | ( n1296 & ~n1297 ) ;
  assign n1299 = ( n1274 & n1295 ) | ( n1274 & ~n1298 ) | ( n1295 & ~n1298 ) ;
  assign n1300 = ( ~n795 & n823 ) | ( ~n795 & n824 ) | ( n823 & n824 ) ;
  assign n1301 = ~x130 & n1300 ;
  assign n1302 = ( n1116 & ~n1117 ) | ( n1116 & n1301 ) | ( ~n1117 & n1301 ) ;
  assign n1303 = ( ~n781 & n809 ) | ( ~n781 & n810 ) | ( n809 & n810 ) ;
  assign n1304 = ~x130 & n1303 ;
  assign n1305 = ( n1120 & ~n1121 ) | ( n1120 & n1304 ) | ( ~n1121 & n1304 ) ;
  assign n1306 = x133 & ~n1305 ;
  assign n1307 = x133 & ~n1302 ;
  assign n1308 = ( n1302 & ~n1306 ) | ( n1302 & n1307 ) | ( ~n1306 & n1307 ) ;
  assign n1309 = ~x132 & n1308 ;
  assign n1310 = ( ~n825 & n840 ) | ( ~n825 & n841 ) | ( n840 & n841 ) ;
  assign n1311 = ~x130 & n1310 ;
  assign n1312 = ( n1126 & ~n1127 ) | ( n1126 & n1311 ) | ( ~n1127 & n1311 ) ;
  assign n1313 = ( n793 & n794 ) | ( n793 & ~n811 ) | ( n794 & ~n811 ) ;
  assign n1314 = ~x130 & n1313 ;
  assign n1315 = ( n1130 & ~n1131 ) | ( n1130 & n1314 ) | ( ~n1131 & n1314 ) ;
  assign n1316 = x133 & ~n1315 ;
  assign n1317 = x133 & ~n1312 ;
  assign n1318 = ( n1312 & ~n1316 ) | ( n1312 & n1317 ) | ( ~n1316 & n1317 ) ;
  assign n1319 = ~x132 & n1318 ;
  assign n1320 = ( n1308 & ~n1309 ) | ( n1308 & n1319 ) | ( ~n1309 & n1319 ) ;
  assign n1321 = ( ~n856 & n884 ) | ( ~n856 & n885 ) | ( n884 & n885 ) ;
  assign n1322 = ~x130 & n1321 ;
  assign n1323 = ( n1137 & ~n1138 ) | ( n1137 & n1322 ) | ( ~n1138 & n1322 ) ;
  assign n1324 = ( ~n842 & n870 ) | ( ~n842 & n871 ) | ( n870 & n871 ) ;
  assign n1325 = ~x130 & n1324 ;
  assign n1326 = ( n1141 & ~n1142 ) | ( n1141 & n1325 ) | ( ~n1142 & n1325 ) ;
  assign n1327 = x133 & ~n1326 ;
  assign n1328 = x133 & ~n1323 ;
  assign n1329 = ( n1323 & ~n1327 ) | ( n1323 & n1328 ) | ( ~n1327 & n1328 ) ;
  assign n1330 = ~x132 & n1329 ;
  assign n1331 = ( n779 & n780 ) | ( n779 & ~n886 ) | ( n780 & ~n886 ) ;
  assign n1332 = ~x130 & n1331 ;
  assign n1333 = ( n1147 & ~n1148 ) | ( n1147 & n1332 ) | ( ~n1148 & n1332 ) ;
  assign n1334 = ( n854 & n855 ) | ( n854 & ~n872 ) | ( n855 & ~n872 ) ;
  assign n1335 = ~x130 & n1334 ;
  assign n1336 = ( n1151 & ~n1152 ) | ( n1151 & n1335 ) | ( ~n1152 & n1335 ) ;
  assign n1337 = x133 & ~n1336 ;
  assign n1338 = x133 & ~n1333 ;
  assign n1339 = ( n1333 & ~n1337 ) | ( n1333 & n1338 ) | ( ~n1337 & n1338 ) ;
  assign n1340 = ~x132 & n1339 ;
  assign n1341 = ( n1329 & ~n1330 ) | ( n1329 & n1340 ) | ( ~n1330 & n1340 ) ;
  assign n1342 = ~x134 & n1320 ;
  assign n1343 = x134 & ~n1341 ;
  assign n1344 = ( x134 & n1342 ) | ( x134 & ~n1343 ) | ( n1342 & ~n1343 ) ;
  assign n1345 = ( n1320 & n1341 ) | ( n1320 & ~n1344 ) | ( n1341 & ~n1344 ) ;
  assign n1346 = ( ~n921 & n948 ) | ( ~n921 & n949 ) | ( n948 & n949 ) ;
  assign n1347 = ~x130 & n1346 ;
  assign n1348 = ( n1162 & ~n1163 ) | ( n1162 & n1347 ) | ( ~n1163 & n1347 ) ;
  assign n1349 = ( ~n907 & n934 ) | ( ~n907 & n935 ) | ( n934 & n935 ) ;
  assign n1350 = ~x130 & n1349 ;
  assign n1351 = ( n1166 & ~n1167 ) | ( n1166 & n1350 ) | ( ~n1167 & n1350 ) ;
  assign n1352 = x133 & ~n1351 ;
  assign n1353 = x133 & ~n1348 ;
  assign n1354 = ( n1348 & ~n1352 ) | ( n1348 & n1353 ) | ( ~n1352 & n1353 ) ;
  assign n1355 = ~x132 & n1354 ;
  assign n1356 = ( ~n951 & n965 ) | ( ~n951 & n966 ) | ( n965 & n966 ) ;
  assign n1357 = ~x130 & n1356 ;
  assign n1358 = ( n1172 & ~n1173 ) | ( n1172 & n1357 ) | ( ~n1173 & n1357 ) ;
  assign n1359 = ( n918 & n919 ) | ( n918 & ~n937 ) | ( n919 & ~n937 ) ;
  assign n1360 = ~x130 & n1359 ;
  assign n1361 = ( n1176 & ~n1177 ) | ( n1176 & n1360 ) | ( ~n1177 & n1360 ) ;
  assign n1362 = x133 & ~n1361 ;
  assign n1363 = x133 & ~n1358 ;
  assign n1364 = ( n1358 & ~n1362 ) | ( n1358 & n1363 ) | ( ~n1362 & n1363 ) ;
  assign n1365 = ~x132 & n1364 ;
  assign n1366 = ( n1354 & ~n1355 ) | ( n1354 & n1365 ) | ( ~n1355 & n1365 ) ;
  assign n1367 = ( ~n982 & n1009 ) | ( ~n982 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1368 = ~x130 & n1367 ;
  assign n1369 = ( n1183 & ~n1184 ) | ( n1183 & n1368 ) | ( ~n1184 & n1368 ) ;
  assign n1370 = ( ~n968 & n995 ) | ( ~n968 & n996 ) | ( n995 & n996 ) ;
  assign n1371 = ~x130 & n1370 ;
  assign n1372 = ( n1187 & ~n1188 ) | ( n1187 & n1371 ) | ( ~n1188 & n1371 ) ;
  assign n1373 = x133 & ~n1372 ;
  assign n1374 = x133 & ~n1369 ;
  assign n1375 = ( n1369 & ~n1373 ) | ( n1369 & n1374 ) | ( ~n1373 & n1374 ) ;
  assign n1376 = ~x132 & n1375 ;
  assign n1377 = ( n904 & n905 ) | ( n904 & ~n1012 ) | ( n905 & ~n1012 ) ;
  assign n1378 = ~x130 & n1377 ;
  assign n1379 = ( n1193 & ~n1194 ) | ( n1193 & n1378 ) | ( ~n1194 & n1378 ) ;
  assign n1380 = ( n979 & n980 ) | ( n979 & ~n998 ) | ( n980 & ~n998 ) ;
  assign n1381 = ~x130 & n1380 ;
  assign n1382 = ( n1197 & ~n1198 ) | ( n1197 & n1381 ) | ( ~n1198 & n1381 ) ;
  assign n1383 = x133 & ~n1382 ;
  assign n1384 = x133 & ~n1379 ;
  assign n1385 = ( n1379 & ~n1383 ) | ( n1379 & n1384 ) | ( ~n1383 & n1384 ) ;
  assign n1386 = ~x132 & n1385 ;
  assign n1387 = ( n1375 & ~n1376 ) | ( n1375 & n1386 ) | ( ~n1376 & n1386 ) ;
  assign n1388 = ~x134 & n1366 ;
  assign n1389 = x134 & ~n1387 ;
  assign n1390 = ( x134 & n1388 ) | ( x134 & ~n1389 ) | ( n1388 & ~n1389 ) ;
  assign n1391 = ( n1366 & n1387 ) | ( n1366 & ~n1390 ) | ( n1387 & ~n1390 ) ;
  assign n1392 = ( n297 & n1212 ) | ( n297 & ~n1213 ) | ( n1212 & ~n1213 ) ;
  assign n1393 = ( n251 & n1208 ) | ( n251 & ~n1209 ) | ( n1208 & ~n1209 ) ;
  assign n1394 = x133 & ~n1393 ;
  assign n1395 = x133 & ~n1392 ;
  assign n1396 = ( n1392 & ~n1394 ) | ( n1392 & n1395 ) | ( ~n1394 & n1395 ) ;
  assign n1397 = ~x132 & n1396 ;
  assign n1398 = ( n346 & n1222 ) | ( n346 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1399 = ( n203 & n1218 ) | ( n203 & ~n1219 ) | ( n1218 & ~n1219 ) ;
  assign n1400 = x133 & ~n1399 ;
  assign n1401 = x133 & ~n1398 ;
  assign n1402 = ( n1398 & ~n1400 ) | ( n1398 & n1401 ) | ( ~n1400 & n1401 ) ;
  assign n1403 = ~x132 & n1402 ;
  assign n1404 = ( n1396 & ~n1397 ) | ( n1396 & n1403 ) | ( ~n1397 & n1403 ) ;
  assign n1405 = ( n440 & n1229 ) | ( n440 & ~n1230 ) | ( n1229 & ~n1230 ) ;
  assign n1406 = x133 & ~n1405 ;
  assign n1407 = ~x130 & n507 ;
  assign n1408 = ( n1233 & ~n1234 ) | ( n1233 & n1407 ) | ( ~n1234 & n1407 ) ;
  assign n1409 = x133 & ~n1408 ;
  assign n1410 = ( ~n1406 & n1408 ) | ( ~n1406 & n1409 ) | ( n1408 & n1409 ) ;
  assign n1411 = ~x132 & n1410 ;
  assign n1412 = ( n157 & n1243 ) | ( n157 & ~n1244 ) | ( n1243 & ~n1244 ) ;
  assign n1413 = ( n392 & n1239 ) | ( n392 & ~n1240 ) | ( n1239 & ~n1240 ) ;
  assign n1414 = x133 & ~n1413 ;
  assign n1415 = x133 & ~n1412 ;
  assign n1416 = ( n1412 & ~n1414 ) | ( n1412 & n1415 ) | ( ~n1414 & n1415 ) ;
  assign n1417 = ~x132 & n1416 ;
  assign n1418 = ( n1410 & ~n1411 ) | ( n1410 & n1417 ) | ( ~n1411 & n1417 ) ;
  assign n1419 = ~x134 & n1404 ;
  assign n1420 = x134 & ~n1418 ;
  assign n1421 = ( x134 & n1419 ) | ( x134 & ~n1420 ) | ( n1419 & ~n1420 ) ;
  assign n1422 = ( n1404 & n1418 ) | ( n1404 & ~n1421 ) | ( n1418 & ~n1421 ) ;
  assign n1423 = ( n623 & n1258 ) | ( n623 & ~n1259 ) | ( n1258 & ~n1259 ) ;
  assign n1424 = ( n593 & n1254 ) | ( n593 & ~n1255 ) | ( n1254 & ~n1255 ) ;
  assign n1425 = x133 & ~n1424 ;
  assign n1426 = x133 & ~n1423 ;
  assign n1427 = ( n1423 & ~n1425 ) | ( n1423 & n1426 ) | ( ~n1425 & n1426 ) ;
  assign n1428 = ~x132 & n1427 ;
  assign n1429 = ( n656 & n1268 ) | ( n656 & ~n1269 ) | ( n1268 & ~n1269 ) ;
  assign n1430 = ( n561 & n1264 ) | ( n561 & ~n1265 ) | ( n1264 & ~n1265 ) ;
  assign n1431 = x133 & ~n1430 ;
  assign n1432 = x133 & ~n1429 ;
  assign n1433 = ( n1429 & ~n1431 ) | ( n1429 & n1432 ) | ( ~n1431 & n1432 ) ;
  assign n1434 = ~x132 & n1433 ;
  assign n1435 = ( n1427 & ~n1428 ) | ( n1427 & n1434 ) | ( ~n1428 & n1434 ) ;
  assign n1436 = ( n748 & n1279 ) | ( n748 & ~n1280 ) | ( n1279 & ~n1280 ) ;
  assign n1437 = ( n718 & n1275 ) | ( n718 & ~n1276 ) | ( n1275 & ~n1276 ) ;
  assign n1438 = x133 & ~n1437 ;
  assign n1439 = x133 & ~n1436 ;
  assign n1440 = ( n1436 & ~n1438 ) | ( n1436 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1441 = ~x132 & n1440 ;
  assign n1442 = ( n531 & n1289 ) | ( n531 & ~n1290 ) | ( n1289 & ~n1290 ) ;
  assign n1443 = ( n686 & n1285 ) | ( n686 & ~n1286 ) | ( n1285 & ~n1286 ) ;
  assign n1444 = x133 & ~n1443 ;
  assign n1445 = x133 & ~n1442 ;
  assign n1446 = ( n1442 & ~n1444 ) | ( n1442 & n1445 ) | ( ~n1444 & n1445 ) ;
  assign n1447 = ~x132 & n1446 ;
  assign n1448 = ( n1440 & ~n1441 ) | ( n1440 & n1447 ) | ( ~n1441 & n1447 ) ;
  assign n1449 = ~x134 & n1435 ;
  assign n1450 = x134 & ~n1448 ;
  assign n1451 = ( x134 & n1449 ) | ( x134 & ~n1450 ) | ( n1449 & ~n1450 ) ;
  assign n1452 = ( n1435 & n1448 ) | ( n1435 & ~n1451 ) | ( n1448 & ~n1451 ) ;
  assign n1453 = ( n821 & n1300 ) | ( n821 & ~n1301 ) | ( n1300 & ~n1301 ) ;
  assign n1454 = ( n807 & n1303 ) | ( n807 & ~n1304 ) | ( n1303 & ~n1304 ) ;
  assign n1455 = x133 & ~n1454 ;
  assign n1456 = x133 & ~n1453 ;
  assign n1457 = ( n1453 & ~n1455 ) | ( n1453 & n1456 ) | ( ~n1455 & n1456 ) ;
  assign n1458 = ~x132 & n1457 ;
  assign n1459 = ( n838 & n1310 ) | ( n838 & ~n1311 ) | ( n1310 & ~n1311 ) ;
  assign n1460 = ( n791 & n1313 ) | ( n791 & ~n1314 ) | ( n1313 & ~n1314 ) ;
  assign n1461 = x133 & ~n1460 ;
  assign n1462 = x133 & ~n1459 ;
  assign n1463 = ( n1459 & ~n1461 ) | ( n1459 & n1462 ) | ( ~n1461 & n1462 ) ;
  assign n1464 = ~x132 & n1463 ;
  assign n1465 = ( n1457 & ~n1458 ) | ( n1457 & n1464 ) | ( ~n1458 & n1464 ) ;
  assign n1466 = ( n882 & n1321 ) | ( n882 & ~n1322 ) | ( n1321 & ~n1322 ) ;
  assign n1467 = ( n868 & n1324 ) | ( n868 & ~n1325 ) | ( n1324 & ~n1325 ) ;
  assign n1468 = x133 & ~n1467 ;
  assign n1469 = x133 & ~n1466 ;
  assign n1470 = ( n1466 & ~n1468 ) | ( n1466 & n1469 ) | ( ~n1468 & n1469 ) ;
  assign n1471 = ~x132 & n1470 ;
  assign n1472 = ( n777 & n1331 ) | ( n777 & ~n1332 ) | ( n1331 & ~n1332 ) ;
  assign n1473 = ( n852 & n1334 ) | ( n852 & ~n1335 ) | ( n1334 & ~n1335 ) ;
  assign n1474 = x133 & ~n1473 ;
  assign n1475 = x133 & ~n1472 ;
  assign n1476 = ( n1472 & ~n1474 ) | ( n1472 & n1475 ) | ( ~n1474 & n1475 ) ;
  assign n1477 = ~x132 & n1476 ;
  assign n1478 = ( n1470 & ~n1471 ) | ( n1470 & n1477 ) | ( ~n1471 & n1477 ) ;
  assign n1479 = ~x134 & n1465 ;
  assign n1480 = x134 & ~n1478 ;
  assign n1481 = ( x134 & n1479 ) | ( x134 & ~n1480 ) | ( n1479 & ~n1480 ) ;
  assign n1482 = ( n1465 & n1478 ) | ( n1465 & ~n1481 ) | ( n1478 & ~n1481 ) ;
  assign n1483 = ( n947 & n1346 ) | ( n947 & ~n1347 ) | ( n1346 & ~n1347 ) ;
  assign n1484 = ( n933 & n1349 ) | ( n933 & ~n1350 ) | ( n1349 & ~n1350 ) ;
  assign n1485 = x133 & ~n1484 ;
  assign n1486 = x133 & ~n1483 ;
  assign n1487 = ( n1483 & ~n1485 ) | ( n1483 & n1486 ) | ( ~n1485 & n1486 ) ;
  assign n1488 = ~x132 & n1487 ;
  assign n1489 = ( n964 & n1356 ) | ( n964 & ~n1357 ) | ( n1356 & ~n1357 ) ;
  assign n1490 = ( n917 & n1359 ) | ( n917 & ~n1360 ) | ( n1359 & ~n1360 ) ;
  assign n1491 = x133 & ~n1490 ;
  assign n1492 = x133 & ~n1489 ;
  assign n1493 = ( n1489 & ~n1491 ) | ( n1489 & n1492 ) | ( ~n1491 & n1492 ) ;
  assign n1494 = ~x132 & n1493 ;
  assign n1495 = ( n1487 & ~n1488 ) | ( n1487 & n1494 ) | ( ~n1488 & n1494 ) ;
  assign n1496 = ( n1008 & n1367 ) | ( n1008 & ~n1368 ) | ( n1367 & ~n1368 ) ;
  assign n1497 = ( n994 & n1370 ) | ( n994 & ~n1371 ) | ( n1370 & ~n1371 ) ;
  assign n1498 = x133 & ~n1497 ;
  assign n1499 = x133 & ~n1496 ;
  assign n1500 = ( n1496 & ~n1498 ) | ( n1496 & n1499 ) | ( ~n1498 & n1499 ) ;
  assign n1501 = ~x132 & n1500 ;
  assign n1502 = ( n903 & n1377 ) | ( n903 & ~n1378 ) | ( n1377 & ~n1378 ) ;
  assign n1503 = ( n978 & n1380 ) | ( n978 & ~n1381 ) | ( n1380 & ~n1381 ) ;
  assign n1504 = x133 & ~n1503 ;
  assign n1505 = x133 & ~n1502 ;
  assign n1506 = ( n1502 & ~n1504 ) | ( n1502 & n1505 ) | ( ~n1504 & n1505 ) ;
  assign n1507 = ~x132 & n1506 ;
  assign n1508 = ( n1500 & ~n1501 ) | ( n1500 & n1507 ) | ( ~n1501 & n1507 ) ;
  assign n1509 = ~x134 & n1495 ;
  assign n1510 = x134 & ~n1508 ;
  assign n1511 = ( x134 & n1509 ) | ( x134 & ~n1510 ) | ( n1509 & ~n1510 ) ;
  assign n1512 = ( n1495 & n1508 ) | ( n1495 & ~n1511 ) | ( n1508 & ~n1511 ) ;
  assign n1513 = ( ~n227 & n369 ) | ( ~n227 & n370 ) | ( n369 & n370 ) ;
  assign n1514 = ~x132 & n1513 ;
  assign n1515 = ( n322 & ~n323 ) | ( n322 & n1514 ) | ( ~n323 & n1514 ) ;
  assign n1516 = ( n180 & n181 ) | ( n180 & ~n416 ) | ( n181 & ~n416 ) ;
  assign n1517 = ~x132 & n1516 ;
  assign n1518 = ( n511 & ~n512 ) | ( n511 & n1517 ) | ( ~n512 & n1517 ) ;
  assign n1519 = ~x134 & n1515 ;
  assign n1520 = x134 & ~n1518 ;
  assign n1521 = ( x134 & n1519 ) | ( x134 & ~n1520 ) | ( n1519 & ~n1520 ) ;
  assign n1522 = ( n1515 & n1518 ) | ( n1515 & ~n1521 ) | ( n1518 & ~n1521 ) ;
  assign n1523 = ( ~n577 & n671 ) | ( ~n577 & n672 ) | ( n671 & n672 ) ;
  assign n1524 = ~x132 & n1523 ;
  assign n1525 = ( n640 & ~n641 ) | ( n640 & n1524 ) | ( ~n641 & n1524 ) ;
  assign n1526 = ( n546 & n547 ) | ( n546 & ~n702 ) | ( n547 & ~n702 ) ;
  assign n1527 = ~x132 & n1526 ;
  assign n1528 = ( n765 & ~n766 ) | ( n765 & n1527 ) | ( ~n766 & n1527 ) ;
  assign n1529 = ~x134 & n1525 ;
  assign n1530 = x134 & ~n1528 ;
  assign n1531 = ( x134 & n1529 ) | ( x134 & ~n1530 ) | ( n1529 & ~n1530 ) ;
  assign n1532 = ( n1525 & n1528 ) | ( n1525 & ~n1531 ) | ( n1528 & ~n1531 ) ;
  assign n1533 = ( ~n799 & n845 ) | ( ~n799 & n846 ) | ( n845 & n846 ) ;
  assign n1534 = ~x132 & n1533 ;
  assign n1535 = ( n830 & ~n831 ) | ( n830 & n1534 ) | ( ~n831 & n1534 ) ;
  assign n1536 = ( n784 & n785 ) | ( n784 & ~n860 ) | ( n785 & ~n860 ) ;
  assign n1537 = ~x132 & n1536 ;
  assign n1538 = ( n891 & ~n892 ) | ( n891 & n1537 ) | ( ~n892 & n1537 ) ;
  assign n1539 = ~x134 & n1535 ;
  assign n1540 = x134 & ~n1538 ;
  assign n1541 = ( x134 & n1539 ) | ( x134 & ~n1540 ) | ( n1539 & ~n1540 ) ;
  assign n1542 = ( n1535 & n1538 ) | ( n1535 & ~n1541 ) | ( n1538 & ~n1541 ) ;
  assign n1543 = ( ~n925 & n971 ) | ( ~n925 & n972 ) | ( n971 & n972 ) ;
  assign n1544 = ~x132 & n1543 ;
  assign n1545 = ( n956 & ~n957 ) | ( n956 & n1544 ) | ( ~n957 & n1544 ) ;
  assign n1546 = ( n910 & n911 ) | ( n910 & ~n986 ) | ( n911 & ~n986 ) ;
  assign n1547 = ~x132 & n1546 ;
  assign n1548 = ( n1017 & ~n1018 ) | ( n1017 & n1547 ) | ( ~n1018 & n1547 ) ;
  assign n1549 = ~x134 & n1545 ;
  assign n1550 = x134 & ~n1548 ;
  assign n1551 = ( x134 & n1549 ) | ( x134 & ~n1550 ) | ( n1549 & ~n1550 ) ;
  assign n1552 = ( n1545 & n1548 ) | ( n1545 & ~n1551 ) | ( n1548 & ~n1551 ) ;
  assign n1553 = ( n1027 & n1051 ) | ( n1027 & ~n1052 ) | ( n1051 & ~n1052 ) ;
  assign n1554 = ~x132 & n1553 ;
  assign n1555 = ( n1063 & ~n1064 ) | ( n1063 & n1554 ) | ( ~n1064 & n1554 ) ;
  assign n1556 = ( n1030 & ~n1031 ) | ( n1030 & n1048 ) | ( ~n1031 & n1048 ) ;
  assign n1557 = ~x132 & n1556 ;
  assign n1558 = ( n1042 & ~n1043 ) | ( n1042 & n1557 ) | ( ~n1043 & n1557 ) ;
  assign n1559 = ~x134 & n1558 ;
  assign n1560 = x134 & ~n1555 ;
  assign n1561 = ( x134 & n1559 ) | ( x134 & ~n1560 ) | ( n1559 & ~n1560 ) ;
  assign n1562 = ( n1555 & n1558 ) | ( n1555 & ~n1561 ) | ( n1558 & ~n1561 ) ;
  assign n1563 = ( n1073 & n1097 ) | ( n1073 & ~n1098 ) | ( n1097 & ~n1098 ) ;
  assign n1564 = ~x132 & n1563 ;
  assign n1565 = ( n1109 & ~n1110 ) | ( n1109 & n1564 ) | ( ~n1110 & n1564 ) ;
  assign n1566 = ( n1076 & ~n1077 ) | ( n1076 & n1094 ) | ( ~n1077 & n1094 ) ;
  assign n1567 = ~x132 & n1566 ;
  assign n1568 = ( n1088 & ~n1089 ) | ( n1088 & n1567 ) | ( ~n1089 & n1567 ) ;
  assign n1569 = ~x134 & n1568 ;
  assign n1570 = x134 & ~n1565 ;
  assign n1571 = ( x134 & n1569 ) | ( x134 & ~n1570 ) | ( n1569 & ~n1570 ) ;
  assign n1572 = ( n1565 & n1568 ) | ( n1565 & ~n1571 ) | ( n1568 & ~n1571 ) ;
  assign n1573 = ( n1119 & n1143 ) | ( n1119 & ~n1144 ) | ( n1143 & ~n1144 ) ;
  assign n1574 = ~x132 & n1573 ;
  assign n1575 = ( n1134 & ~n1135 ) | ( n1134 & n1574 ) | ( ~n1135 & n1574 ) ;
  assign n1576 = ( n1122 & ~n1123 ) | ( n1122 & n1140 ) | ( ~n1123 & n1140 ) ;
  assign n1577 = ~x132 & n1576 ;
  assign n1578 = ( n1155 & ~n1156 ) | ( n1155 & n1577 ) | ( ~n1156 & n1577 ) ;
  assign n1579 = ~x134 & n1575 ;
  assign n1580 = x134 & ~n1578 ;
  assign n1581 = ( x134 & n1579 ) | ( x134 & ~n1580 ) | ( n1579 & ~n1580 ) ;
  assign n1582 = ( n1575 & n1578 ) | ( n1575 & ~n1581 ) | ( n1578 & ~n1581 ) ;
  assign n1583 = ( n1165 & n1189 ) | ( n1165 & ~n1190 ) | ( n1189 & ~n1190 ) ;
  assign n1584 = ~x132 & n1583 ;
  assign n1585 = ( n1180 & ~n1181 ) | ( n1180 & n1584 ) | ( ~n1181 & n1584 ) ;
  assign n1586 = ( n1168 & ~n1169 ) | ( n1168 & n1186 ) | ( ~n1169 & n1186 ) ;
  assign n1587 = ~x132 & n1586 ;
  assign n1588 = ( n1201 & ~n1202 ) | ( n1201 & n1587 ) | ( ~n1202 & n1587 ) ;
  assign n1589 = ~x134 & n1585 ;
  assign n1590 = x134 & ~n1588 ;
  assign n1591 = ( x134 & n1589 ) | ( x134 & ~n1590 ) | ( n1589 & ~n1590 ) ;
  assign n1592 = ( n1585 & n1588 ) | ( n1585 & ~n1591 ) | ( n1588 & ~n1591 ) ;
  assign n1593 = ( ~n1215 & n1231 ) | ( ~n1215 & n1232 ) | ( n1231 & n1232 ) ;
  assign n1594 = ~x132 & n1593 ;
  assign n1595 = ( n1226 & ~n1227 ) | ( n1226 & n1594 ) | ( ~n1227 & n1594 ) ;
  assign n1596 = ( n1210 & n1211 ) | ( n1210 & ~n1236 ) | ( n1211 & ~n1236 ) ;
  assign n1597 = ~x132 & n1596 ;
  assign n1598 = ( n1247 & ~n1248 ) | ( n1247 & n1597 ) | ( ~n1248 & n1597 ) ;
  assign n1599 = ~x134 & n1595 ;
  assign n1600 = x134 & ~n1598 ;
  assign n1601 = ( x134 & n1599 ) | ( x134 & ~n1600 ) | ( n1599 & ~n1600 ) ;
  assign n1602 = ( n1595 & n1598 ) | ( n1595 & ~n1601 ) | ( n1598 & ~n1601 ) ;
  assign n1603 = ( ~n1261 & n1277 ) | ( ~n1261 & n1278 ) | ( n1277 & n1278 ) ;
  assign n1604 = ~x132 & n1603 ;
  assign n1605 = ( n1272 & ~n1273 ) | ( n1272 & n1604 ) | ( ~n1273 & n1604 ) ;
  assign n1606 = ( n1256 & n1257 ) | ( n1256 & ~n1282 ) | ( n1257 & ~n1282 ) ;
  assign n1607 = ~x132 & n1606 ;
  assign n1608 = ( n1293 & ~n1294 ) | ( n1293 & n1607 ) | ( ~n1294 & n1607 ) ;
  assign n1609 = ~x134 & n1605 ;
  assign n1610 = x134 & ~n1608 ;
  assign n1611 = ( x134 & n1609 ) | ( x134 & ~n1610 ) | ( n1609 & ~n1610 ) ;
  assign n1612 = ( n1605 & n1608 ) | ( n1605 & ~n1611 ) | ( n1608 & ~n1611 ) ;
  assign n1613 = ( ~n1307 & n1326 ) | ( ~n1307 & n1327 ) | ( n1326 & n1327 ) ;
  assign n1614 = ~x132 & n1613 ;
  assign n1615 = ( n1318 & ~n1319 ) | ( n1318 & n1614 ) | ( ~n1319 & n1614 ) ;
  assign n1616 = ( n1305 & n1306 ) | ( n1305 & ~n1328 ) | ( n1306 & ~n1328 ) ;
  assign n1617 = ~x132 & n1616 ;
  assign n1618 = ( n1339 & ~n1340 ) | ( n1339 & n1617 ) | ( ~n1340 & n1617 ) ;
  assign n1619 = ~x134 & n1615 ;
  assign n1620 = x134 & ~n1618 ;
  assign n1621 = ( x134 & n1619 ) | ( x134 & ~n1620 ) | ( n1619 & ~n1620 ) ;
  assign n1622 = ( n1615 & n1618 ) | ( n1615 & ~n1621 ) | ( n1618 & ~n1621 ) ;
  assign n1623 = ( ~n1353 & n1372 ) | ( ~n1353 & n1373 ) | ( n1372 & n1373 ) ;
  assign n1624 = ~x132 & n1623 ;
  assign n1625 = ( n1364 & ~n1365 ) | ( n1364 & n1624 ) | ( ~n1365 & n1624 ) ;
  assign n1626 = ( n1351 & n1352 ) | ( n1351 & ~n1374 ) | ( n1352 & ~n1374 ) ;
  assign n1627 = ~x132 & n1626 ;
  assign n1628 = ( n1385 & ~n1386 ) | ( n1385 & n1627 ) | ( ~n1386 & n1627 ) ;
  assign n1629 = ~x134 & n1625 ;
  assign n1630 = x134 & ~n1628 ;
  assign n1631 = ( x134 & n1629 ) | ( x134 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1632 = ( n1625 & n1628 ) | ( n1625 & ~n1631 ) | ( n1628 & ~n1631 ) ;
  assign n1633 = ( ~n1395 & n1405 ) | ( ~n1395 & n1406 ) | ( n1405 & n1406 ) ;
  assign n1634 = ~x132 & n1633 ;
  assign n1635 = ( n1402 & ~n1403 ) | ( n1402 & n1634 ) | ( ~n1403 & n1634 ) ;
  assign n1636 = ( n1393 & n1394 ) | ( n1393 & ~n1409 ) | ( n1394 & ~n1409 ) ;
  assign n1637 = ~x132 & n1636 ;
  assign n1638 = ( n1416 & ~n1417 ) | ( n1416 & n1637 ) | ( ~n1417 & n1637 ) ;
  assign n1639 = ~x134 & n1635 ;
  assign n1640 = x134 & ~n1638 ;
  assign n1641 = ( x134 & n1639 ) | ( x134 & ~n1640 ) | ( n1639 & ~n1640 ) ;
  assign n1642 = ( n1635 & n1638 ) | ( n1635 & ~n1641 ) | ( n1638 & ~n1641 ) ;
  assign n1643 = ( ~n1426 & n1437 ) | ( ~n1426 & n1438 ) | ( n1437 & n1438 ) ;
  assign n1644 = ~x132 & n1643 ;
  assign n1645 = ( n1433 & ~n1434 ) | ( n1433 & n1644 ) | ( ~n1434 & n1644 ) ;
  assign n1646 = ( n1424 & n1425 ) | ( n1424 & ~n1439 ) | ( n1425 & ~n1439 ) ;
  assign n1647 = ~x132 & n1646 ;
  assign n1648 = ( n1446 & ~n1447 ) | ( n1446 & n1647 ) | ( ~n1447 & n1647 ) ;
  assign n1649 = ~x134 & n1645 ;
  assign n1650 = x134 & ~n1648 ;
  assign n1651 = ( x134 & n1649 ) | ( x134 & ~n1650 ) | ( n1649 & ~n1650 ) ;
  assign n1652 = ( n1645 & n1648 ) | ( n1645 & ~n1651 ) | ( n1648 & ~n1651 ) ;
  assign n1653 = ( ~n1456 & n1467 ) | ( ~n1456 & n1468 ) | ( n1467 & n1468 ) ;
  assign n1654 = ~x132 & n1653 ;
  assign n1655 = ( n1463 & ~n1464 ) | ( n1463 & n1654 ) | ( ~n1464 & n1654 ) ;
  assign n1656 = ( n1454 & n1455 ) | ( n1454 & ~n1469 ) | ( n1455 & ~n1469 ) ;
  assign n1657 = ~x132 & n1656 ;
  assign n1658 = ( n1476 & ~n1477 ) | ( n1476 & n1657 ) | ( ~n1477 & n1657 ) ;
  assign n1659 = ~x134 & n1655 ;
  assign n1660 = x134 & ~n1658 ;
  assign n1661 = ( x134 & n1659 ) | ( x134 & ~n1660 ) | ( n1659 & ~n1660 ) ;
  assign n1662 = ( n1655 & n1658 ) | ( n1655 & ~n1661 ) | ( n1658 & ~n1661 ) ;
  assign n1663 = ( ~n1486 & n1497 ) | ( ~n1486 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1664 = ~x132 & n1663 ;
  assign n1665 = ( n1493 & ~n1494 ) | ( n1493 & n1664 ) | ( ~n1494 & n1664 ) ;
  assign n1666 = ( n1484 & n1485 ) | ( n1484 & ~n1499 ) | ( n1485 & ~n1499 ) ;
  assign n1667 = ~x132 & n1666 ;
  assign n1668 = ( n1506 & ~n1507 ) | ( n1506 & n1667 ) | ( ~n1507 & n1667 ) ;
  assign n1669 = ~x134 & n1665 ;
  assign n1670 = x134 & ~n1668 ;
  assign n1671 = ( x134 & n1669 ) | ( x134 & ~n1670 ) | ( n1669 & ~n1670 ) ;
  assign n1672 = ( n1665 & n1668 ) | ( n1665 & ~n1671 ) | ( n1668 & ~n1671 ) ;
  assign n1673 = ( ~n321 & n463 ) | ( ~n321 & n464 ) | ( n463 & n464 ) ;
  assign n1674 = ~x132 & n1673 ;
  assign n1675 = ( n1513 & ~n1514 ) | ( n1513 & n1674 ) | ( ~n1514 & n1674 ) ;
  assign n1676 = ( n274 & n275 ) | ( n274 & ~n510 ) | ( n275 & ~n510 ) ;
  assign n1677 = ~x132 & n1676 ;
  assign n1678 = ( n1516 & ~n1517 ) | ( n1516 & n1677 ) | ( ~n1517 & n1677 ) ;
  assign n1679 = ~x134 & n1675 ;
  assign n1680 = x134 & ~n1678 ;
  assign n1681 = ( x134 & n1679 ) | ( x134 & ~n1680 ) | ( n1679 & ~n1680 ) ;
  assign n1682 = ( n1675 & n1678 ) | ( n1675 & ~n1681 ) | ( n1678 & ~n1681 ) ;
  assign n1683 = ( ~n639 & n733 ) | ( ~n639 & n734 ) | ( n733 & n734 ) ;
  assign n1684 = ~x132 & n1683 ;
  assign n1685 = ( n1523 & ~n1524 ) | ( n1523 & n1684 ) | ( ~n1524 & n1684 ) ;
  assign n1686 = ( n608 & n609 ) | ( n608 & ~n764 ) | ( n609 & ~n764 ) ;
  assign n1687 = ~x132 & n1686 ;
  assign n1688 = ( n1526 & ~n1527 ) | ( n1526 & n1687 ) | ( ~n1527 & n1687 ) ;
  assign n1689 = ~x134 & n1685 ;
  assign n1690 = x134 & ~n1688 ;
  assign n1691 = ( x134 & n1689 ) | ( x134 & ~n1690 ) | ( n1689 & ~n1690 ) ;
  assign n1692 = ( n1685 & n1688 ) | ( n1685 & ~n1691 ) | ( n1688 & ~n1691 ) ;
  assign n1693 = ( ~n829 & n875 ) | ( ~n829 & n876 ) | ( n875 & n876 ) ;
  assign n1694 = ~x132 & n1693 ;
  assign n1695 = ( n1533 & ~n1534 ) | ( n1533 & n1694 ) | ( ~n1534 & n1694 ) ;
  assign n1696 = ( n814 & n815 ) | ( n814 & ~n890 ) | ( n815 & ~n890 ) ;
  assign n1697 = ~x132 & n1696 ;
  assign n1698 = ( n1536 & ~n1537 ) | ( n1536 & n1697 ) | ( ~n1537 & n1697 ) ;
  assign n1699 = ~x134 & n1695 ;
  assign n1700 = x134 & ~n1698 ;
  assign n1701 = ( x134 & n1699 ) | ( x134 & ~n1700 ) | ( n1699 & ~n1700 ) ;
  assign n1702 = ( n1695 & n1698 ) | ( n1695 & ~n1701 ) | ( n1698 & ~n1701 ) ;
  assign n1703 = ( ~n955 & n1001 ) | ( ~n955 & n1002 ) | ( n1001 & n1002 ) ;
  assign n1704 = ~x132 & n1703 ;
  assign n1705 = ( n1543 & ~n1544 ) | ( n1543 & n1704 ) | ( ~n1544 & n1704 ) ;
  assign n1706 = ( n940 & n941 ) | ( n940 & ~n1016 ) | ( n941 & ~n1016 ) ;
  assign n1707 = ~x132 & n1706 ;
  assign n1708 = ( n1546 & ~n1547 ) | ( n1546 & n1707 ) | ( ~n1547 & n1707 ) ;
  assign n1709 = ~x134 & n1705 ;
  assign n1710 = x134 & ~n1708 ;
  assign n1711 = ( x134 & n1709 ) | ( x134 & ~n1710 ) | ( n1709 & ~n1710 ) ;
  assign n1712 = ( n1705 & n1708 ) | ( n1705 & ~n1711 ) | ( n1708 & ~n1711 ) ;
  assign n1713 = ( n1040 & ~n1041 ) | ( n1040 & n1058 ) | ( ~n1041 & n1058 ) ;
  assign n1714 = ~x132 & n1713 ;
  assign n1715 = ( n1556 & ~n1557 ) | ( n1556 & n1714 ) | ( ~n1557 & n1714 ) ;
  assign n1716 = ( n1037 & n1061 ) | ( n1037 & ~n1062 ) | ( n1061 & ~n1062 ) ;
  assign n1717 = ~x132 & n1716 ;
  assign n1718 = ( n1553 & ~n1554 ) | ( n1553 & n1717 ) | ( ~n1554 & n1717 ) ;
  assign n1719 = ~x134 & n1715 ;
  assign n1720 = x134 & ~n1718 ;
  assign n1721 = ( x134 & n1719 ) | ( x134 & ~n1720 ) | ( n1719 & ~n1720 ) ;
  assign n1722 = ( n1715 & n1718 ) | ( n1715 & ~n1721 ) | ( n1718 & ~n1721 ) ;
  assign n1723 = ( n1086 & ~n1087 ) | ( n1086 & n1104 ) | ( ~n1087 & n1104 ) ;
  assign n1724 = ~x132 & n1723 ;
  assign n1725 = ( n1566 & ~n1567 ) | ( n1566 & n1724 ) | ( ~n1567 & n1724 ) ;
  assign n1726 = ( n1083 & n1107 ) | ( n1083 & ~n1108 ) | ( n1107 & ~n1108 ) ;
  assign n1727 = ~x132 & n1726 ;
  assign n1728 = ( n1563 & ~n1564 ) | ( n1563 & n1727 ) | ( ~n1564 & n1727 ) ;
  assign n1729 = ~x134 & n1725 ;
  assign n1730 = x134 & ~n1728 ;
  assign n1731 = ( x134 & n1729 ) | ( x134 & ~n1730 ) | ( n1729 & ~n1730 ) ;
  assign n1732 = ( n1725 & n1728 ) | ( n1725 & ~n1731 ) | ( n1728 & ~n1731 ) ;
  assign n1733 = ( n1129 & n1153 ) | ( n1129 & ~n1154 ) | ( n1153 & ~n1154 ) ;
  assign n1734 = ~x132 & n1733 ;
  assign n1735 = ( n1573 & ~n1574 ) | ( n1573 & n1734 ) | ( ~n1574 & n1734 ) ;
  assign n1736 = ( n1132 & ~n1133 ) | ( n1132 & n1150 ) | ( ~n1133 & n1150 ) ;
  assign n1737 = ~x132 & n1736 ;
  assign n1738 = ( n1576 & ~n1577 ) | ( n1576 & n1737 ) | ( ~n1577 & n1737 ) ;
  assign n1739 = ~x134 & n1735 ;
  assign n1740 = x134 & ~n1738 ;
  assign n1741 = ( x134 & n1739 ) | ( x134 & ~n1740 ) | ( n1739 & ~n1740 ) ;
  assign n1742 = ( n1735 & n1738 ) | ( n1735 & ~n1741 ) | ( n1738 & ~n1741 ) ;
  assign n1743 = ( n1175 & n1199 ) | ( n1175 & ~n1200 ) | ( n1199 & ~n1200 ) ;
  assign n1744 = ~x132 & n1743 ;
  assign n1745 = ( n1583 & ~n1584 ) | ( n1583 & n1744 ) | ( ~n1584 & n1744 ) ;
  assign n1746 = ( n1178 & ~n1179 ) | ( n1178 & n1196 ) | ( ~n1179 & n1196 ) ;
  assign n1747 = ~x132 & n1746 ;
  assign n1748 = ( n1586 & ~n1587 ) | ( n1586 & n1747 ) | ( ~n1587 & n1747 ) ;
  assign n1749 = ~x134 & n1745 ;
  assign n1750 = x134 & ~n1748 ;
  assign n1751 = ( x134 & n1749 ) | ( x134 & ~n1750 ) | ( n1749 & ~n1750 ) ;
  assign n1752 = ( n1745 & n1748 ) | ( n1745 & ~n1751 ) | ( n1748 & ~n1751 ) ;
  assign n1753 = ( ~n1225 & n1241 ) | ( ~n1225 & n1242 ) | ( n1241 & n1242 ) ;
  assign n1754 = ~x132 & n1753 ;
  assign n1755 = ( n1593 & ~n1594 ) | ( n1593 & n1754 ) | ( ~n1594 & n1754 ) ;
  assign n1756 = ( n1220 & n1221 ) | ( n1220 & ~n1246 ) | ( n1221 & ~n1246 ) ;
  assign n1757 = ~x132 & n1756 ;
  assign n1758 = ( n1596 & ~n1597 ) | ( n1596 & n1757 ) | ( ~n1597 & n1757 ) ;
  assign n1759 = ~x134 & n1755 ;
  assign n1760 = x134 & ~n1758 ;
  assign n1761 = ( x134 & n1759 ) | ( x134 & ~n1760 ) | ( n1759 & ~n1760 ) ;
  assign n1762 = ( n1755 & n1758 ) | ( n1755 & ~n1761 ) | ( n1758 & ~n1761 ) ;
  assign n1763 = ( ~n1271 & n1287 ) | ( ~n1271 & n1288 ) | ( n1287 & n1288 ) ;
  assign n1764 = ~x132 & n1763 ;
  assign n1765 = ( n1603 & ~n1604 ) | ( n1603 & n1764 ) | ( ~n1604 & n1764 ) ;
  assign n1766 = ( n1266 & n1267 ) | ( n1266 & ~n1292 ) | ( n1267 & ~n1292 ) ;
  assign n1767 = ~x132 & n1766 ;
  assign n1768 = ( n1606 & ~n1607 ) | ( n1606 & n1767 ) | ( ~n1607 & n1767 ) ;
  assign n1769 = ~x134 & n1765 ;
  assign n1770 = x134 & ~n1768 ;
  assign n1771 = ( x134 & n1769 ) | ( x134 & ~n1770 ) | ( n1769 & ~n1770 ) ;
  assign n1772 = ( n1765 & n1768 ) | ( n1765 & ~n1771 ) | ( n1768 & ~n1771 ) ;
  assign n1773 = ( ~n1317 & n1336 ) | ( ~n1317 & n1337 ) | ( n1336 & n1337 ) ;
  assign n1774 = ~x132 & n1773 ;
  assign n1775 = ( n1613 & ~n1614 ) | ( n1613 & n1774 ) | ( ~n1614 & n1774 ) ;
  assign n1776 = ( n1315 & n1316 ) | ( n1315 & ~n1338 ) | ( n1316 & ~n1338 ) ;
  assign n1777 = ~x132 & n1776 ;
  assign n1778 = ( n1616 & ~n1617 ) | ( n1616 & n1777 ) | ( ~n1617 & n1777 ) ;
  assign n1779 = ~x134 & n1775 ;
  assign n1780 = x134 & ~n1778 ;
  assign n1781 = ( x134 & n1779 ) | ( x134 & ~n1780 ) | ( n1779 & ~n1780 ) ;
  assign n1782 = ( n1775 & n1778 ) | ( n1775 & ~n1781 ) | ( n1778 & ~n1781 ) ;
  assign n1783 = ( ~n1363 & n1382 ) | ( ~n1363 & n1383 ) | ( n1382 & n1383 ) ;
  assign n1784 = ~x132 & n1783 ;
  assign n1785 = ( n1623 & ~n1624 ) | ( n1623 & n1784 ) | ( ~n1624 & n1784 ) ;
  assign n1786 = ( n1361 & n1362 ) | ( n1361 & ~n1384 ) | ( n1362 & ~n1384 ) ;
  assign n1787 = ~x132 & n1786 ;
  assign n1788 = ( n1626 & ~n1627 ) | ( n1626 & n1787 ) | ( ~n1627 & n1787 ) ;
  assign n1789 = ~x134 & n1785 ;
  assign n1790 = x134 & ~n1788 ;
  assign n1791 = ( x134 & n1789 ) | ( x134 & ~n1790 ) | ( n1789 & ~n1790 ) ;
  assign n1792 = ( n1785 & n1788 ) | ( n1785 & ~n1791 ) | ( n1788 & ~n1791 ) ;
  assign n1793 = ( ~n1401 & n1413 ) | ( ~n1401 & n1414 ) | ( n1413 & n1414 ) ;
  assign n1794 = ~x132 & n1793 ;
  assign n1795 = ( n1633 & ~n1634 ) | ( n1633 & n1794 ) | ( ~n1634 & n1794 ) ;
  assign n1796 = ( n1399 & n1400 ) | ( n1399 & ~n1415 ) | ( n1400 & ~n1415 ) ;
  assign n1797 = ~x132 & n1796 ;
  assign n1798 = ( n1636 & ~n1637 ) | ( n1636 & n1797 ) | ( ~n1637 & n1797 ) ;
  assign n1799 = ~x134 & n1795 ;
  assign n1800 = x134 & ~n1798 ;
  assign n1801 = ( x134 & n1799 ) | ( x134 & ~n1800 ) | ( n1799 & ~n1800 ) ;
  assign n1802 = ( n1795 & n1798 ) | ( n1795 & ~n1801 ) | ( n1798 & ~n1801 ) ;
  assign n1803 = ( ~n1432 & n1443 ) | ( ~n1432 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1804 = ~x132 & n1803 ;
  assign n1805 = ( n1643 & ~n1644 ) | ( n1643 & n1804 ) | ( ~n1644 & n1804 ) ;
  assign n1806 = ( n1430 & n1431 ) | ( n1430 & ~n1445 ) | ( n1431 & ~n1445 ) ;
  assign n1807 = ~x132 & n1806 ;
  assign n1808 = ( n1646 & ~n1647 ) | ( n1646 & n1807 ) | ( ~n1647 & n1807 ) ;
  assign n1809 = ~x134 & n1805 ;
  assign n1810 = x134 & ~n1808 ;
  assign n1811 = ( x134 & n1809 ) | ( x134 & ~n1810 ) | ( n1809 & ~n1810 ) ;
  assign n1812 = ( n1805 & n1808 ) | ( n1805 & ~n1811 ) | ( n1808 & ~n1811 ) ;
  assign n1813 = ( ~n1462 & n1473 ) | ( ~n1462 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1814 = ~x132 & n1813 ;
  assign n1815 = ( n1653 & ~n1654 ) | ( n1653 & n1814 ) | ( ~n1654 & n1814 ) ;
  assign n1816 = ( n1460 & n1461 ) | ( n1460 & ~n1475 ) | ( n1461 & ~n1475 ) ;
  assign n1817 = ~x132 & n1816 ;
  assign n1818 = ( n1656 & ~n1657 ) | ( n1656 & n1817 ) | ( ~n1657 & n1817 ) ;
  assign n1819 = ~x134 & n1815 ;
  assign n1820 = x134 & ~n1818 ;
  assign n1821 = ( x134 & n1819 ) | ( x134 & ~n1820 ) | ( n1819 & ~n1820 ) ;
  assign n1822 = ( n1815 & n1818 ) | ( n1815 & ~n1821 ) | ( n1818 & ~n1821 ) ;
  assign n1823 = ( ~n1492 & n1503 ) | ( ~n1492 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1824 = ~x132 & n1823 ;
  assign n1825 = ( n1663 & ~n1664 ) | ( n1663 & n1824 ) | ( ~n1664 & n1824 ) ;
  assign n1826 = ( n1490 & n1491 ) | ( n1490 & ~n1505 ) | ( n1491 & ~n1505 ) ;
  assign n1827 = ~x132 & n1826 ;
  assign n1828 = ( n1666 & ~n1667 ) | ( n1666 & n1827 ) | ( ~n1667 & n1827 ) ;
  assign n1829 = ~x134 & n1825 ;
  assign n1830 = x134 & ~n1828 ;
  assign n1831 = ( x134 & n1829 ) | ( x134 & ~n1830 ) | ( n1829 & ~n1830 ) ;
  assign n1832 = ( n1825 & n1828 ) | ( n1825 & ~n1831 ) | ( n1828 & ~n1831 ) ;
  assign n1833 = ( n418 & n1673 ) | ( n418 & ~n1674 ) | ( n1673 & ~n1674 ) ;
  assign n1834 = ( n229 & n1676 ) | ( n229 & ~n1677 ) | ( n1676 & ~n1677 ) ;
  assign n1835 = ~x134 & n1833 ;
  assign n1836 = x134 & ~n1834 ;
  assign n1837 = ( x134 & n1835 ) | ( x134 & ~n1836 ) | ( n1835 & ~n1836 ) ;
  assign n1838 = ( n1833 & n1834 ) | ( n1833 & ~n1837 ) | ( n1834 & ~n1837 ) ;
  assign n1839 = ( n704 & n1683 ) | ( n704 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1840 = ( n579 & n1686 ) | ( n579 & ~n1687 ) | ( n1686 & ~n1687 ) ;
  assign n1841 = ~x134 & n1839 ;
  assign n1842 = x134 & ~n1840 ;
  assign n1843 = ( x134 & n1841 ) | ( x134 & ~n1842 ) | ( n1841 & ~n1842 ) ;
  assign n1844 = ( n1839 & n1840 ) | ( n1839 & ~n1843 ) | ( n1840 & ~n1843 ) ;
  assign n1845 = ( n862 & n1693 ) | ( n862 & ~n1694 ) | ( n1693 & ~n1694 ) ;
  assign n1846 = ( n801 & n1696 ) | ( n801 & ~n1697 ) | ( n1696 & ~n1697 ) ;
  assign n1847 = ~x134 & n1845 ;
  assign n1848 = x134 & ~n1846 ;
  assign n1849 = ( x134 & n1847 ) | ( x134 & ~n1848 ) | ( n1847 & ~n1848 ) ;
  assign n1850 = ( n1845 & n1846 ) | ( n1845 & ~n1849 ) | ( n1846 & ~n1849 ) ;
  assign n1851 = ( n988 & n1703 ) | ( n988 & ~n1704 ) | ( n1703 & ~n1704 ) ;
  assign n1852 = ( n927 & n1706 ) | ( n927 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1853 = ~x134 & n1851 ;
  assign n1854 = x134 & ~n1852 ;
  assign n1855 = ( x134 & n1853 ) | ( x134 & ~n1854 ) | ( n1853 & ~n1854 ) ;
  assign n1856 = ( n1851 & n1852 ) | ( n1851 & ~n1855 ) | ( n1852 & ~n1855 ) ;
  assign n1857 = x132 & ~n1713 ;
  assign n1858 = ( n1053 & n1054 ) | ( n1053 & ~n1857 ) | ( n1054 & ~n1857 ) ;
  assign n1859 = x132 & ~n1716 ;
  assign n1860 = ( n1032 & n1033 ) | ( n1032 & ~n1859 ) | ( n1033 & ~n1859 ) ;
  assign n1861 = ~x134 & n1858 ;
  assign n1862 = x134 & ~n1860 ;
  assign n1863 = ( x134 & n1861 ) | ( x134 & ~n1862 ) | ( n1861 & ~n1862 ) ;
  assign n1864 = ( n1858 & n1860 ) | ( n1858 & ~n1863 ) | ( n1860 & ~n1863 ) ;
  assign n1865 = x132 & ~n1723 ;
  assign n1866 = ( n1099 & n1100 ) | ( n1099 & ~n1865 ) | ( n1100 & ~n1865 ) ;
  assign n1867 = x132 & ~n1726 ;
  assign n1868 = ( n1078 & n1079 ) | ( n1078 & ~n1867 ) | ( n1079 & ~n1867 ) ;
  assign n1869 = ~x134 & n1866 ;
  assign n1870 = x134 & ~n1868 ;
  assign n1871 = ( x134 & n1869 ) | ( x134 & ~n1870 ) | ( n1869 & ~n1870 ) ;
  assign n1872 = ( n1866 & n1868 ) | ( n1866 & ~n1871 ) | ( n1868 & ~n1871 ) ;
  assign n1873 = x132 & ~n1733 ;
  assign n1874 = ( n1145 & n1146 ) | ( n1145 & ~n1873 ) | ( n1146 & ~n1873 ) ;
  assign n1875 = x132 & ~n1736 ;
  assign n1876 = ( n1124 & n1125 ) | ( n1124 & ~n1875 ) | ( n1125 & ~n1875 ) ;
  assign n1877 = ~x134 & n1874 ;
  assign n1878 = x134 & ~n1876 ;
  assign n1879 = ( x134 & n1877 ) | ( x134 & ~n1878 ) | ( n1877 & ~n1878 ) ;
  assign n1880 = ( n1874 & n1876 ) | ( n1874 & ~n1879 ) | ( n1876 & ~n1879 ) ;
  assign n1881 = x132 & ~n1743 ;
  assign n1882 = ( n1191 & n1192 ) | ( n1191 & ~n1881 ) | ( n1192 & ~n1881 ) ;
  assign n1883 = x132 & ~n1746 ;
  assign n1884 = ( n1170 & n1171 ) | ( n1170 & ~n1883 ) | ( n1171 & ~n1883 ) ;
  assign n1885 = ~x134 & n1882 ;
  assign n1886 = x134 & ~n1884 ;
  assign n1887 = ( x134 & n1885 ) | ( x134 & ~n1886 ) | ( n1885 & ~n1886 ) ;
  assign n1888 = ( n1882 & n1884 ) | ( n1882 & ~n1887 ) | ( n1884 & ~n1887 ) ;
  assign n1889 = ( n1238 & n1753 ) | ( n1238 & ~n1754 ) | ( n1753 & ~n1754 ) ;
  assign n1890 = ( n1217 & n1756 ) | ( n1217 & ~n1757 ) | ( n1756 & ~n1757 ) ;
  assign n1891 = ~x134 & n1889 ;
  assign n1892 = x134 & ~n1890 ;
  assign n1893 = ( x134 & n1891 ) | ( x134 & ~n1892 ) | ( n1891 & ~n1892 ) ;
  assign n1894 = ( n1889 & n1890 ) | ( n1889 & ~n1893 ) | ( n1890 & ~n1893 ) ;
  assign n1895 = ( n1263 & n1766 ) | ( n1263 & ~n1767 ) | ( n1766 & ~n1767 ) ;
  assign n1896 = ( n1284 & n1763 ) | ( n1284 & ~n1764 ) | ( n1763 & ~n1764 ) ;
  assign n1897 = ~x134 & n1896 ;
  assign n1898 = x134 & ~n1895 ;
  assign n1899 = ( x134 & n1897 ) | ( x134 & ~n1898 ) | ( n1897 & ~n1898 ) ;
  assign n1900 = ( n1895 & n1896 ) | ( n1895 & ~n1899 ) | ( n1896 & ~n1899 ) ;
  assign n1901 = ( n1330 & n1773 ) | ( n1330 & ~n1774 ) | ( n1773 & ~n1774 ) ;
  assign n1902 = ( n1309 & n1776 ) | ( n1309 & ~n1777 ) | ( n1776 & ~n1777 ) ;
  assign n1903 = ~x134 & n1901 ;
  assign n1904 = x134 & ~n1902 ;
  assign n1905 = ( x134 & n1903 ) | ( x134 & ~n1904 ) | ( n1903 & ~n1904 ) ;
  assign n1906 = ( n1901 & n1902 ) | ( n1901 & ~n1905 ) | ( n1902 & ~n1905 ) ;
  assign n1907 = ( n1355 & n1786 ) | ( n1355 & ~n1787 ) | ( n1786 & ~n1787 ) ;
  assign n1908 = ( n1376 & n1783 ) | ( n1376 & ~n1784 ) | ( n1783 & ~n1784 ) ;
  assign n1909 = ~x134 & n1908 ;
  assign n1910 = x134 & ~n1907 ;
  assign n1911 = ( x134 & n1909 ) | ( x134 & ~n1910 ) | ( n1909 & ~n1910 ) ;
  assign n1912 = ( n1907 & n1908 ) | ( n1907 & ~n1911 ) | ( n1908 & ~n1911 ) ;
  assign n1913 = ( n1397 & n1796 ) | ( n1397 & ~n1797 ) | ( n1796 & ~n1797 ) ;
  assign n1914 = ( n1411 & n1793 ) | ( n1411 & ~n1794 ) | ( n1793 & ~n1794 ) ;
  assign n1915 = ~x134 & n1914 ;
  assign n1916 = x134 & ~n1913 ;
  assign n1917 = ( x134 & n1915 ) | ( x134 & ~n1916 ) | ( n1915 & ~n1916 ) ;
  assign n1918 = ( n1913 & n1914 ) | ( n1913 & ~n1917 ) | ( n1914 & ~n1917 ) ;
  assign n1919 = ( n1428 & n1806 ) | ( n1428 & ~n1807 ) | ( n1806 & ~n1807 ) ;
  assign n1920 = ( n1441 & n1803 ) | ( n1441 & ~n1804 ) | ( n1803 & ~n1804 ) ;
  assign n1921 = ~x134 & n1920 ;
  assign n1922 = x134 & ~n1919 ;
  assign n1923 = ( x134 & n1921 ) | ( x134 & ~n1922 ) | ( n1921 & ~n1922 ) ;
  assign n1924 = ( n1919 & n1920 ) | ( n1919 & ~n1923 ) | ( n1920 & ~n1923 ) ;
  assign n1925 = ( n1471 & n1813 ) | ( n1471 & ~n1814 ) | ( n1813 & ~n1814 ) ;
  assign n1926 = ( n1458 & n1816 ) | ( n1458 & ~n1817 ) | ( n1816 & ~n1817 ) ;
  assign n1927 = ~x134 & n1925 ;
  assign n1928 = x134 & ~n1926 ;
  assign n1929 = ( x134 & n1927 ) | ( x134 & ~n1928 ) | ( n1927 & ~n1928 ) ;
  assign n1930 = ( n1925 & n1926 ) | ( n1925 & ~n1929 ) | ( n1926 & ~n1929 ) ;
  assign n1931 = ( n1488 & n1826 ) | ( n1488 & ~n1827 ) | ( n1826 & ~n1827 ) ;
  assign n1932 = ( n1501 & n1823 ) | ( n1501 & ~n1824 ) | ( n1823 & ~n1824 ) ;
  assign n1933 = ~x134 & n1932 ;
  assign n1934 = x134 & ~n1931 ;
  assign n1935 = ( x134 & n1933 ) | ( x134 & ~n1934 ) | ( n1933 & ~n1934 ) ;
  assign n1936 = ( n1931 & n1932 ) | ( n1931 & ~n1935 ) | ( n1932 & ~n1935 ) ;
  assign y0 = n517 ;
  assign y1 = n771 ;
  assign y2 = n897 ;
  assign y3 = n1023 ;
  assign y4 = n1069 ;
  assign y5 = n1115 ;
  assign y6 = n1161 ;
  assign y7 = n1207 ;
  assign y8 = n1253 ;
  assign y9 = n1299 ;
  assign y10 = n1345 ;
  assign y11 = n1391 ;
  assign y12 = n1422 ;
  assign y13 = n1452 ;
  assign y14 = n1482 ;
  assign y15 = n1512 ;
  assign y16 = n1522 ;
  assign y17 = n1532 ;
  assign y18 = n1542 ;
  assign y19 = n1552 ;
  assign y20 = n1562 ;
  assign y21 = n1572 ;
  assign y22 = n1582 ;
  assign y23 = n1592 ;
  assign y24 = n1602 ;
  assign y25 = n1612 ;
  assign y26 = n1622 ;
  assign y27 = n1632 ;
  assign y28 = n1642 ;
  assign y29 = n1652 ;
  assign y30 = n1662 ;
  assign y31 = n1672 ;
  assign y32 = n1682 ;
  assign y33 = n1692 ;
  assign y34 = n1702 ;
  assign y35 = n1712 ;
  assign y36 = n1722 ;
  assign y37 = n1732 ;
  assign y38 = n1742 ;
  assign y39 = n1752 ;
  assign y40 = n1762 ;
  assign y41 = n1772 ;
  assign y42 = n1782 ;
  assign y43 = n1792 ;
  assign y44 = n1802 ;
  assign y45 = n1812 ;
  assign y46 = n1822 ;
  assign y47 = n1832 ;
  assign y48 = n1838 ;
  assign y49 = n1844 ;
  assign y50 = n1850 ;
  assign y51 = n1856 ;
  assign y52 = n1864 ;
  assign y53 = n1872 ;
  assign y54 = n1880 ;
  assign y55 = n1888 ;
  assign y56 = n1894 ;
  assign y57 = n1900 ;
  assign y58 = n1906 ;
  assign y59 = n1912 ;
  assign y60 = n1918 ;
  assign y61 = n1924 ;
  assign y62 = n1930 ;
  assign y63 = n1936 ;
  assign y64 = n516 ;
  assign y65 = n770 ;
  assign y66 = n896 ;
  assign y67 = n1022 ;
  assign y68 = n1068 ;
  assign y69 = n1114 ;
  assign y70 = n1160 ;
  assign y71 = n1206 ;
  assign y72 = n1252 ;
  assign y73 = n1298 ;
  assign y74 = n1344 ;
  assign y75 = n1390 ;
  assign y76 = n1421 ;
  assign y77 = n1451 ;
  assign y78 = n1481 ;
  assign y79 = n1511 ;
  assign y80 = n1521 ;
  assign y81 = n1531 ;
  assign y82 = n1541 ;
  assign y83 = n1551 ;
  assign y84 = n1561 ;
  assign y85 = n1571 ;
  assign y86 = n1581 ;
  assign y87 = n1591 ;
  assign y88 = n1601 ;
  assign y89 = n1611 ;
  assign y90 = n1621 ;
  assign y91 = n1631 ;
  assign y92 = n1641 ;
  assign y93 = n1651 ;
  assign y94 = n1661 ;
  assign y95 = n1671 ;
  assign y96 = n1681 ;
  assign y97 = n1691 ;
  assign y98 = n1701 ;
  assign y99 = n1711 ;
  assign y100 = n1721 ;
  assign y101 = n1731 ;
  assign y102 = n1741 ;
  assign y103 = n1751 ;
  assign y104 = n1761 ;
  assign y105 = n1771 ;
  assign y106 = n1781 ;
  assign y107 = n1791 ;
  assign y108 = n1801 ;
  assign y109 = n1811 ;
  assign y110 = n1821 ;
  assign y111 = n1831 ;
  assign y112 = n1837 ;
  assign y113 = n1843 ;
  assign y114 = n1849 ;
  assign y115 = n1855 ;
  assign y116 = n1863 ;
  assign y117 = n1871 ;
  assign y118 = n1879 ;
  assign y119 = n1887 ;
  assign y120 = n1893 ;
  assign y121 = n1899 ;
  assign y122 = n1905 ;
  assign y123 = n1911 ;
  assign y124 = n1917 ;
  assign y125 = n1923 ;
  assign y126 = n1929 ;
  assign y127 = n1935 ;
endmodule
