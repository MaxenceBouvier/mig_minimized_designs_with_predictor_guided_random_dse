module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 ;
  assign n1002 = ( x835 & x836 ) | ( x835 & x837 ) | ( x836 & x837 ) ;
  assign n1003 = ( ~x835 & x836 ) | ( ~x835 & x837 ) | ( x836 & x837 ) ;
  assign n1004 = ( x835 & ~n1002 ) | ( x835 & n1003 ) | ( ~n1002 & n1003 ) ;
  assign n1005 = ( x838 & x839 ) | ( x838 & x840 ) | ( x839 & x840 ) ;
  assign n1006 = ( ~x838 & x839 ) | ( ~x838 & x840 ) | ( x839 & x840 ) ;
  assign n1007 = ( x838 & ~n1005 ) | ( x838 & n1006 ) | ( ~n1005 & n1006 ) ;
  assign n1008 = n1004 & n1007 ;
  assign n1009 = n1004 | n1007 ;
  assign n1010 = ~n1008 & n1009 ;
  assign n1011 = ( x841 & x842 ) | ( x841 & x843 ) | ( x842 & x843 ) ;
  assign n1012 = ( ~x841 & x842 ) | ( ~x841 & x843 ) | ( x842 & x843 ) ;
  assign n1013 = ( x841 & ~n1011 ) | ( x841 & n1012 ) | ( ~n1011 & n1012 ) ;
  assign n1014 = ( x844 & x845 ) | ( x844 & x846 ) | ( x845 & x846 ) ;
  assign n1015 = ( ~x844 & x845 ) | ( ~x844 & x846 ) | ( x845 & x846 ) ;
  assign n1016 = ( x844 & ~n1014 ) | ( x844 & n1015 ) | ( ~n1014 & n1015 ) ;
  assign n1017 = ( n1010 & n1013 ) | ( n1010 & n1016 ) | ( n1013 & n1016 ) ;
  assign n1018 = ( ~n1010 & n1013 ) | ( ~n1010 & n1016 ) | ( n1013 & n1016 ) ;
  assign n1019 = ( n1010 & ~n1017 ) | ( n1010 & n1018 ) | ( ~n1017 & n1018 ) ;
  assign n1020 = ( x829 & x830 ) | ( x829 & x831 ) | ( x830 & x831 ) ;
  assign n1021 = ( ~x829 & x830 ) | ( ~x829 & x831 ) | ( x830 & x831 ) ;
  assign n1022 = ( x829 & ~n1020 ) | ( x829 & n1021 ) | ( ~n1020 & n1021 ) ;
  assign n1023 = ( x832 & x833 ) | ( x832 & x834 ) | ( x833 & x834 ) ;
  assign n1024 = ( ~x832 & x833 ) | ( ~x832 & x834 ) | ( x833 & x834 ) ;
  assign n1025 = ( x832 & ~n1023 ) | ( x832 & n1024 ) | ( ~n1023 & n1024 ) ;
  assign n1026 = ( x823 & x824 ) | ( x823 & x825 ) | ( x824 & x825 ) ;
  assign n1027 = ( ~x823 & x824 ) | ( ~x823 & x825 ) | ( x824 & x825 ) ;
  assign n1028 = ( x823 & ~n1026 ) | ( x823 & n1027 ) | ( ~n1026 & n1027 ) ;
  assign n1029 = ( x826 & x827 ) | ( x826 & x828 ) | ( x827 & x828 ) ;
  assign n1030 = ( ~x826 & x827 ) | ( ~x826 & x828 ) | ( x827 & x828 ) ;
  assign n1031 = ( x826 & ~n1029 ) | ( x826 & n1030 ) | ( ~n1029 & n1030 ) ;
  assign n1032 = n1028 & n1031 ;
  assign n1033 = n1028 | n1031 ;
  assign n1034 = ~n1032 & n1033 ;
  assign n1035 = ( n1022 & n1025 ) | ( n1022 & n1034 ) | ( n1025 & n1034 ) ;
  assign n1036 = ( ~n1022 & n1025 ) | ( ~n1022 & n1034 ) | ( n1025 & n1034 ) ;
  assign n1037 = ( n1022 & ~n1035 ) | ( n1022 & n1036 ) | ( ~n1035 & n1036 ) ;
  assign n1038 = n1019 & n1037 ;
  assign n1039 = n1019 | n1037 ;
  assign n1040 = ~n1038 & n1039 ;
  assign n1041 = ( x814 & x815 ) | ( x814 & x816 ) | ( x815 & x816 ) ;
  assign n1042 = ( ~x814 & x815 ) | ( ~x814 & x816 ) | ( x815 & x816 ) ;
  assign n1043 = ( x814 & ~n1041 ) | ( x814 & n1042 ) | ( ~n1041 & n1042 ) ;
  assign n1044 = ( x811 & x812 ) | ( x811 & x813 ) | ( x812 & x813 ) ;
  assign n1045 = ( ~x811 & x812 ) | ( ~x811 & x813 ) | ( x812 & x813 ) ;
  assign n1046 = ( x811 & ~n1044 ) | ( x811 & n1045 ) | ( ~n1044 & n1045 ) ;
  assign n1047 = n1043 & n1046 ;
  assign n1048 = n1043 | n1046 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = ( x817 & x818 ) | ( x817 & x819 ) | ( x818 & x819 ) ;
  assign n1051 = ( ~x817 & x818 ) | ( ~x817 & x819 ) | ( x818 & x819 ) ;
  assign n1052 = ( x817 & ~n1050 ) | ( x817 & n1051 ) | ( ~n1050 & n1051 ) ;
  assign n1053 = ( x820 & x821 ) | ( x820 & x822 ) | ( x821 & x822 ) ;
  assign n1054 = ( ~x820 & x821 ) | ( ~x820 & x822 ) | ( x821 & x822 ) ;
  assign n1055 = ( x820 & ~n1053 ) | ( x820 & n1054 ) | ( ~n1053 & n1054 ) ;
  assign n1056 = ( n1049 & n1052 ) | ( n1049 & n1055 ) | ( n1052 & n1055 ) ;
  assign n1057 = ( ~n1049 & n1052 ) | ( ~n1049 & n1055 ) | ( n1052 & n1055 ) ;
  assign n1058 = ( n1049 & ~n1056 ) | ( n1049 & n1057 ) | ( ~n1056 & n1057 ) ;
  assign n1059 = ( x802 & x803 ) | ( x802 & x804 ) | ( x803 & x804 ) ;
  assign n1060 = ( ~x802 & x803 ) | ( ~x802 & x804 ) | ( x803 & x804 ) ;
  assign n1061 = ( x802 & ~n1059 ) | ( x802 & n1060 ) | ( ~n1059 & n1060 ) ;
  assign n1062 = ( x799 & x800 ) | ( x799 & x801 ) | ( x800 & x801 ) ;
  assign n1063 = ( ~x799 & x800 ) | ( ~x799 & x801 ) | ( x800 & x801 ) ;
  assign n1064 = ( x799 & ~n1062 ) | ( x799 & n1063 ) | ( ~n1062 & n1063 ) ;
  assign n1065 = n1061 & n1064 ;
  assign n1066 = n1061 | n1064 ;
  assign n1067 = ~n1065 & n1066 ;
  assign n1068 = ( x805 & x806 ) | ( x805 & x807 ) | ( x806 & x807 ) ;
  assign n1069 = ( ~x805 & x806 ) | ( ~x805 & x807 ) | ( x806 & x807 ) ;
  assign n1070 = ( x805 & ~n1068 ) | ( x805 & n1069 ) | ( ~n1068 & n1069 ) ;
  assign n1071 = ( x808 & x809 ) | ( x808 & x810 ) | ( x809 & x810 ) ;
  assign n1072 = ( ~x808 & x809 ) | ( ~x808 & x810 ) | ( x809 & x810 ) ;
  assign n1073 = ( x808 & ~n1071 ) | ( x808 & n1072 ) | ( ~n1071 & n1072 ) ;
  assign n1074 = ( n1067 & n1070 ) | ( n1067 & n1073 ) | ( n1070 & n1073 ) ;
  assign n1075 = ( ~n1067 & n1070 ) | ( ~n1067 & n1073 ) | ( n1070 & n1073 ) ;
  assign n1076 = ( n1067 & ~n1074 ) | ( n1067 & n1075 ) | ( ~n1074 & n1075 ) ;
  assign n1077 = n1058 & n1076 ;
  assign n1078 = n1058 | n1076 ;
  assign n1079 = ~n1077 & n1078 ;
  assign n1080 = ( x778 & x779 ) | ( x778 & x780 ) | ( x779 & x780 ) ;
  assign n1081 = ( ~x778 & x779 ) | ( ~x778 & x780 ) | ( x779 & x780 ) ;
  assign n1082 = ( x778 & ~n1080 ) | ( x778 & n1081 ) | ( ~n1080 & n1081 ) ;
  assign n1083 = ( x775 & x776 ) | ( x775 & x777 ) | ( x776 & x777 ) ;
  assign n1084 = ( ~x775 & x776 ) | ( ~x775 & x777 ) | ( x776 & x777 ) ;
  assign n1085 = ( x775 & ~n1083 ) | ( x775 & n1084 ) | ( ~n1083 & n1084 ) ;
  assign n1086 = n1082 & n1085 ;
  assign n1087 = n1082 | n1085 ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = ( ~x781 & x782 ) | ( ~x781 & x783 ) | ( x782 & x783 ) ;
  assign n1090 = ( x781 & x782 ) | ( x781 & x783 ) | ( x782 & x783 ) ;
  assign n1091 = ( x781 & n1089 ) | ( x781 & ~n1090 ) | ( n1089 & ~n1090 ) ;
  assign n1092 = ( ~x784 & x785 ) | ( ~x784 & x786 ) | ( x785 & x786 ) ;
  assign n1093 = ( x784 & x785 ) | ( x784 & x786 ) | ( x785 & x786 ) ;
  assign n1094 = ( x784 & n1092 ) | ( x784 & ~n1093 ) | ( n1092 & ~n1093 ) ;
  assign n1095 = ( n1088 & n1091 ) | ( n1088 & n1094 ) | ( n1091 & n1094 ) ;
  assign n1096 = ( ~n1088 & n1091 ) | ( ~n1088 & n1094 ) | ( n1091 & n1094 ) ;
  assign n1097 = ( n1088 & ~n1095 ) | ( n1088 & n1096 ) | ( ~n1095 & n1096 ) ;
  assign n1098 = ( x793 & x794 ) | ( x793 & x795 ) | ( x794 & x795 ) ;
  assign n1099 = ( ~x793 & x794 ) | ( ~x793 & x795 ) | ( x794 & x795 ) ;
  assign n1100 = ( x793 & ~n1098 ) | ( x793 & n1099 ) | ( ~n1098 & n1099 ) ;
  assign n1101 = ( x796 & x797 ) | ( x796 & x798 ) | ( x797 & x798 ) ;
  assign n1102 = ( ~x796 & x797 ) | ( ~x796 & x798 ) | ( x797 & x798 ) ;
  assign n1103 = ( x796 & ~n1101 ) | ( x796 & n1102 ) | ( ~n1101 & n1102 ) ;
  assign n1104 = ( x790 & x791 ) | ( x790 & x792 ) | ( x791 & x792 ) ;
  assign n1105 = ( ~x790 & x791 ) | ( ~x790 & x792 ) | ( x791 & x792 ) ;
  assign n1106 = ( x790 & ~n1104 ) | ( x790 & n1105 ) | ( ~n1104 & n1105 ) ;
  assign n1107 = ( x787 & x788 ) | ( x787 & x789 ) | ( x788 & x789 ) ;
  assign n1108 = ( ~x787 & x788 ) | ( ~x787 & x789 ) | ( x788 & x789 ) ;
  assign n1109 = ( x787 & ~n1107 ) | ( x787 & n1108 ) | ( ~n1107 & n1108 ) ;
  assign n1110 = n1106 & n1109 ;
  assign n1111 = n1106 | n1109 ;
  assign n1112 = ~n1110 & n1111 ;
  assign n1113 = ( n1100 & n1103 ) | ( n1100 & n1112 ) | ( n1103 & n1112 ) ;
  assign n1114 = ( ~n1100 & n1103 ) | ( ~n1100 & n1112 ) | ( n1103 & n1112 ) ;
  assign n1115 = ( n1100 & ~n1113 ) | ( n1100 & n1114 ) | ( ~n1113 & n1114 ) ;
  assign n1116 = n1097 & n1115 ;
  assign n1117 = n1097 | n1115 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = ( ~x772 & x773 ) | ( ~x772 & x774 ) | ( x773 & x774 ) ;
  assign n1120 = ( x772 & x773 ) | ( x772 & x774 ) | ( x773 & x774 ) ;
  assign n1121 = ( x772 & n1119 ) | ( x772 & ~n1120 ) | ( n1119 & ~n1120 ) ;
  assign n1122 = ( ~x769 & x770 ) | ( ~x769 & x771 ) | ( x770 & x771 ) ;
  assign n1123 = ( x769 & x770 ) | ( x769 & x771 ) | ( x770 & x771 ) ;
  assign n1124 = ( x769 & n1122 ) | ( x769 & ~n1123 ) | ( n1122 & ~n1123 ) ;
  assign n1125 = ( x766 & x767 ) | ( x766 & x768 ) | ( x767 & x768 ) ;
  assign n1126 = ( ~x766 & x767 ) | ( ~x766 & x768 ) | ( x767 & x768 ) ;
  assign n1127 = ( x766 & ~n1125 ) | ( x766 & n1126 ) | ( ~n1125 & n1126 ) ;
  assign n1128 = ( x763 & x764 ) | ( x763 & x765 ) | ( x764 & x765 ) ;
  assign n1129 = ( ~x763 & x764 ) | ( ~x763 & x765 ) | ( x764 & x765 ) ;
  assign n1130 = ( x763 & ~n1128 ) | ( x763 & n1129 ) | ( ~n1128 & n1129 ) ;
  assign n1131 = n1127 & n1130 ;
  assign n1132 = n1127 | n1130 ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ( n1121 & n1124 ) | ( n1121 & n1133 ) | ( n1124 & n1133 ) ;
  assign n1135 = ( ~n1121 & n1124 ) | ( ~n1121 & n1133 ) | ( n1124 & n1133 ) ;
  assign n1136 = ( n1121 & ~n1134 ) | ( n1121 & n1135 ) | ( ~n1134 & n1135 ) ;
  assign n1137 = ( x751 & x752 ) | ( x751 & x753 ) | ( x752 & x753 ) ;
  assign n1138 = ( ~x751 & x752 ) | ( ~x751 & x753 ) | ( x752 & x753 ) ;
  assign n1139 = ( x751 & ~n1137 ) | ( x751 & n1138 ) | ( ~n1137 & n1138 ) ;
  assign n1140 = ( x754 & x755 ) | ( x754 & x756 ) | ( x755 & x756 ) ;
  assign n1141 = ( ~x754 & x755 ) | ( ~x754 & x756 ) | ( x755 & x756 ) ;
  assign n1142 = ( x754 & ~n1140 ) | ( x754 & n1141 ) | ( ~n1140 & n1141 ) ;
  assign n1143 = n1139 & n1142 ;
  assign n1144 = n1139 | n1142 ;
  assign n1145 = ~n1143 & n1144 ;
  assign n1146 = ( x760 & x761 ) | ( x760 & x762 ) | ( x761 & x762 ) ;
  assign n1147 = ( ~x760 & x761 ) | ( ~x760 & x762 ) | ( x761 & x762 ) ;
  assign n1148 = ( x760 & ~n1146 ) | ( x760 & n1147 ) | ( ~n1146 & n1147 ) ;
  assign n1149 = ( x757 & x758 ) | ( x757 & x759 ) | ( x758 & x759 ) ;
  assign n1150 = ( ~x757 & x758 ) | ( ~x757 & x759 ) | ( x758 & x759 ) ;
  assign n1151 = ( x757 & ~n1149 ) | ( x757 & n1150 ) | ( ~n1149 & n1150 ) ;
  assign n1152 = ( n1145 & n1148 ) | ( n1145 & n1151 ) | ( n1148 & n1151 ) ;
  assign n1153 = ( ~n1145 & n1148 ) | ( ~n1145 & n1151 ) | ( n1148 & n1151 ) ;
  assign n1154 = ( n1145 & ~n1152 ) | ( n1145 & n1153 ) | ( ~n1152 & n1153 ) ;
  assign n1155 = n1136 & n1154 ;
  assign n1156 = n1136 | n1154 ;
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = n1118 & n1157 ;
  assign n1159 = n1118 | n1157 ;
  assign n1160 = ~n1158 & n1159 ;
  assign n1161 = ( n1040 & n1079 ) | ( n1040 & n1160 ) | ( n1079 & n1160 ) ;
  assign n1162 = ( ~n1040 & n1079 ) | ( ~n1040 & n1160 ) | ( n1079 & n1160 ) ;
  assign n1163 = ( n1040 & ~n1161 ) | ( n1040 & n1162 ) | ( ~n1161 & n1162 ) ;
  assign n1164 = ( ~x664 & x665 ) | ( ~x664 & x666 ) | ( x665 & x666 ) ;
  assign n1165 = ( x664 & x665 ) | ( x664 & x666 ) | ( x665 & x666 ) ;
  assign n1166 = ( x664 & n1164 ) | ( x664 & ~n1165 ) | ( n1164 & ~n1165 ) ;
  assign n1167 = ( ~x661 & x662 ) | ( ~x661 & x663 ) | ( x662 & x663 ) ;
  assign n1168 = ( x661 & x662 ) | ( x661 & x663 ) | ( x662 & x663 ) ;
  assign n1169 = ( x661 & n1167 ) | ( x661 & ~n1168 ) | ( n1167 & ~n1168 ) ;
  assign n1170 = ( x655 & x656 ) | ( x655 & x657 ) | ( x656 & x657 ) ;
  assign n1171 = ( ~x655 & x656 ) | ( ~x655 & x657 ) | ( x656 & x657 ) ;
  assign n1172 = ( x655 & ~n1170 ) | ( x655 & n1171 ) | ( ~n1170 & n1171 ) ;
  assign n1173 = ( x658 & x659 ) | ( x658 & x660 ) | ( x659 & x660 ) ;
  assign n1174 = ( ~x658 & x659 ) | ( ~x658 & x660 ) | ( x659 & x660 ) ;
  assign n1175 = ( x658 & ~n1173 ) | ( x658 & n1174 ) | ( ~n1173 & n1174 ) ;
  assign n1176 = n1172 & n1175 ;
  assign n1177 = n1172 | n1175 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1179 = ( n1166 & n1169 ) | ( n1166 & n1178 ) | ( n1169 & n1178 ) ;
  assign n1180 = ( ~n1166 & n1169 ) | ( ~n1166 & n1178 ) | ( n1169 & n1178 ) ;
  assign n1181 = ( n1166 & ~n1179 ) | ( n1166 & n1180 ) | ( ~n1179 & n1180 ) ;
  assign n1182 = ( x667 & x668 ) | ( x667 & x669 ) | ( x668 & x669 ) ;
  assign n1183 = ( ~x667 & x668 ) | ( ~x667 & x669 ) | ( x668 & x669 ) ;
  assign n1184 = ( x667 & ~n1182 ) | ( x667 & n1183 ) | ( ~n1182 & n1183 ) ;
  assign n1185 = ( x670 & x671 ) | ( x670 & x672 ) | ( x671 & x672 ) ;
  assign n1186 = ( ~x670 & x671 ) | ( ~x670 & x672 ) | ( x671 & x672 ) ;
  assign n1187 = ( x670 & ~n1185 ) | ( x670 & n1186 ) | ( ~n1185 & n1186 ) ;
  assign n1188 = n1184 & n1187 ;
  assign n1189 = n1184 | n1187 ;
  assign n1190 = ~n1188 & n1189 ;
  assign n1191 = ( x676 & x677 ) | ( x676 & x678 ) | ( x677 & x678 ) ;
  assign n1192 = ( ~x676 & x677 ) | ( ~x676 & x678 ) | ( x677 & x678 ) ;
  assign n1193 = ( x676 & ~n1191 ) | ( x676 & n1192 ) | ( ~n1191 & n1192 ) ;
  assign n1194 = ( x673 & x674 ) | ( x673 & x675 ) | ( x674 & x675 ) ;
  assign n1195 = ( ~x673 & x674 ) | ( ~x673 & x675 ) | ( x674 & x675 ) ;
  assign n1196 = ( x673 & ~n1194 ) | ( x673 & n1195 ) | ( ~n1194 & n1195 ) ;
  assign n1197 = ( n1190 & n1193 ) | ( n1190 & n1196 ) | ( n1193 & n1196 ) ;
  assign n1198 = ( ~n1190 & n1193 ) | ( ~n1190 & n1196 ) | ( n1193 & n1196 ) ;
  assign n1199 = ( n1190 & ~n1197 ) | ( n1190 & n1198 ) | ( ~n1197 & n1198 ) ;
  assign n1200 = n1181 & n1199 ;
  assign n1201 = n1181 | n1199 ;
  assign n1202 = ~n1200 & n1201 ;
  assign n1203 = ( ~x688 & x689 ) | ( ~x688 & x690 ) | ( x689 & x690 ) ;
  assign n1204 = ( x688 & x689 ) | ( x688 & x690 ) | ( x689 & x690 ) ;
  assign n1205 = ( x688 & n1203 ) | ( x688 & ~n1204 ) | ( n1203 & ~n1204 ) ;
  assign n1206 = ( ~x685 & x686 ) | ( ~x685 & x687 ) | ( x686 & x687 ) ;
  assign n1207 = ( x685 & x686 ) | ( x685 & x687 ) | ( x686 & x687 ) ;
  assign n1208 = ( x685 & n1206 ) | ( x685 & ~n1207 ) | ( n1206 & ~n1207 ) ;
  assign n1209 = ( x679 & x680 ) | ( x679 & x681 ) | ( x680 & x681 ) ;
  assign n1210 = ( ~x679 & x680 ) | ( ~x679 & x681 ) | ( x680 & x681 ) ;
  assign n1211 = ( x679 & ~n1209 ) | ( x679 & n1210 ) | ( ~n1209 & n1210 ) ;
  assign n1212 = ( x682 & x683 ) | ( x682 & x684 ) | ( x683 & x684 ) ;
  assign n1213 = ( ~x682 & x683 ) | ( ~x682 & x684 ) | ( x683 & x684 ) ;
  assign n1214 = ( x682 & ~n1212 ) | ( x682 & n1213 ) | ( ~n1212 & n1213 ) ;
  assign n1215 = n1211 & n1214 ;
  assign n1216 = n1211 | n1214 ;
  assign n1217 = ~n1215 & n1216 ;
  assign n1218 = ( n1205 & n1208 ) | ( n1205 & n1217 ) | ( n1208 & n1217 ) ;
  assign n1219 = ( ~n1205 & n1208 ) | ( ~n1205 & n1217 ) | ( n1208 & n1217 ) ;
  assign n1220 = ( n1205 & ~n1218 ) | ( n1205 & n1219 ) | ( ~n1218 & n1219 ) ;
  assign n1221 = ( x694 & x695 ) | ( x694 & x696 ) | ( x695 & x696 ) ;
  assign n1222 = ( ~x694 & x695 ) | ( ~x694 & x696 ) | ( x695 & x696 ) ;
  assign n1223 = ( x694 & ~n1221 ) | ( x694 & n1222 ) | ( ~n1221 & n1222 ) ;
  assign n1224 = ( x691 & x692 ) | ( x691 & x693 ) | ( x692 & x693 ) ;
  assign n1225 = ( ~x691 & x692 ) | ( ~x691 & x693 ) | ( x692 & x693 ) ;
  assign n1226 = ( x691 & ~n1224 ) | ( x691 & n1225 ) | ( ~n1224 & n1225 ) ;
  assign n1227 = n1223 & n1226 ;
  assign n1228 = n1223 | n1226 ;
  assign n1229 = ~n1227 & n1228 ;
  assign n1230 = ( ~x697 & x698 ) | ( ~x697 & x699 ) | ( x698 & x699 ) ;
  assign n1231 = ( x697 & x698 ) | ( x697 & x699 ) | ( x698 & x699 ) ;
  assign n1232 = ( x697 & n1230 ) | ( x697 & ~n1231 ) | ( n1230 & ~n1231 ) ;
  assign n1233 = ( ~x700 & x701 ) | ( ~x700 & x702 ) | ( x701 & x702 ) ;
  assign n1234 = ( x700 & x701 ) | ( x700 & x702 ) | ( x701 & x702 ) ;
  assign n1235 = ( x700 & n1233 ) | ( x700 & ~n1234 ) | ( n1233 & ~n1234 ) ;
  assign n1236 = ( n1229 & n1232 ) | ( n1229 & n1235 ) | ( n1232 & n1235 ) ;
  assign n1237 = ( ~n1229 & n1232 ) | ( ~n1229 & n1235 ) | ( n1232 & n1235 ) ;
  assign n1238 = ( n1229 & ~n1236 ) | ( n1229 & n1237 ) | ( ~n1236 & n1237 ) ;
  assign n1239 = n1220 & n1238 ;
  assign n1240 = n1220 | n1238 ;
  assign n1241 = ~n1239 & n1240 ;
  assign n1242 = n1202 & n1241 ;
  assign n1243 = n1202 | n1241 ;
  assign n1244 = ~n1242 & n1243 ;
  assign n1245 = ( x742 & x743 ) | ( x742 & x744 ) | ( x743 & x744 ) ;
  assign n1246 = ( ~x742 & x743 ) | ( ~x742 & x744 ) | ( x743 & x744 ) ;
  assign n1247 = ( x742 & ~n1245 ) | ( x742 & n1246 ) | ( ~n1245 & n1246 ) ;
  assign n1248 = ( x739 & x740 ) | ( x739 & x741 ) | ( x740 & x741 ) ;
  assign n1249 = ( ~x739 & x740 ) | ( ~x739 & x741 ) | ( x740 & x741 ) ;
  assign n1250 = ( x739 & ~n1248 ) | ( x739 & n1249 ) | ( ~n1248 & n1249 ) ;
  assign n1251 = n1247 & n1250 ;
  assign n1252 = n1247 | n1250 ;
  assign n1253 = ~n1251 & n1252 ;
  assign n1254 = ( x745 & x746 ) | ( x745 & x747 ) | ( x746 & x747 ) ;
  assign n1255 = ( ~x745 & x746 ) | ( ~x745 & x747 ) | ( x746 & x747 ) ;
  assign n1256 = ( x745 & ~n1254 ) | ( x745 & n1255 ) | ( ~n1254 & n1255 ) ;
  assign n1257 = ( x748 & x749 ) | ( x748 & x750 ) | ( x749 & x750 ) ;
  assign n1258 = ( ~x748 & x749 ) | ( ~x748 & x750 ) | ( x749 & x750 ) ;
  assign n1259 = ( x748 & ~n1257 ) | ( x748 & n1258 ) | ( ~n1257 & n1258 ) ;
  assign n1260 = ( n1253 & n1256 ) | ( n1253 & n1259 ) | ( n1256 & n1259 ) ;
  assign n1261 = ( ~n1253 & n1256 ) | ( ~n1253 & n1259 ) | ( n1256 & n1259 ) ;
  assign n1262 = ( n1253 & ~n1260 ) | ( n1253 & n1261 ) | ( ~n1260 & n1261 ) ;
  assign n1263 = ( x727 & x728 ) | ( x727 & x729 ) | ( x728 & x729 ) ;
  assign n1264 = ( ~x727 & x728 ) | ( ~x727 & x729 ) | ( x728 & x729 ) ;
  assign n1265 = ( x727 & ~n1263 ) | ( x727 & n1264 ) | ( ~n1263 & n1264 ) ;
  assign n1266 = ( x730 & x731 ) | ( x730 & x732 ) | ( x731 & x732 ) ;
  assign n1267 = ( ~x730 & x731 ) | ( ~x730 & x732 ) | ( x731 & x732 ) ;
  assign n1268 = ( x730 & ~n1266 ) | ( x730 & n1267 ) | ( ~n1266 & n1267 ) ;
  assign n1269 = n1265 & n1268 ;
  assign n1270 = n1265 | n1268 ;
  assign n1271 = ~n1269 & n1270 ;
  assign n1272 = ( ~x733 & x734 ) | ( ~x733 & x735 ) | ( x734 & x735 ) ;
  assign n1273 = ( x733 & x734 ) | ( x733 & x735 ) | ( x734 & x735 ) ;
  assign n1274 = ( x733 & n1272 ) | ( x733 & ~n1273 ) | ( n1272 & ~n1273 ) ;
  assign n1275 = ( ~x736 & x737 ) | ( ~x736 & x738 ) | ( x737 & x738 ) ;
  assign n1276 = ( x736 & x737 ) | ( x736 & x738 ) | ( x737 & x738 ) ;
  assign n1277 = ( x736 & n1275 ) | ( x736 & ~n1276 ) | ( n1275 & ~n1276 ) ;
  assign n1278 = ( n1271 & n1274 ) | ( n1271 & n1277 ) | ( n1274 & n1277 ) ;
  assign n1279 = ( ~n1271 & n1274 ) | ( ~n1271 & n1277 ) | ( n1274 & n1277 ) ;
  assign n1280 = ( n1271 & ~n1278 ) | ( n1271 & n1279 ) | ( ~n1278 & n1279 ) ;
  assign n1281 = n1262 & n1280 ;
  assign n1282 = n1262 | n1280 ;
  assign n1283 = ~n1281 & n1282 ;
  assign n1284 = ( x715 & x716 ) | ( x715 & x717 ) | ( x716 & x717 ) ;
  assign n1285 = ( ~x715 & x716 ) | ( ~x715 & x717 ) | ( x716 & x717 ) ;
  assign n1286 = ( x715 & ~n1284 ) | ( x715 & n1285 ) | ( ~n1284 & n1285 ) ;
  assign n1287 = ( x718 & x719 ) | ( x718 & x720 ) | ( x719 & x720 ) ;
  assign n1288 = ( ~x718 & x719 ) | ( ~x718 & x720 ) | ( x719 & x720 ) ;
  assign n1289 = ( x718 & ~n1287 ) | ( x718 & n1288 ) | ( ~n1287 & n1288 ) ;
  assign n1290 = n1286 & n1289 ;
  assign n1291 = n1286 | n1289 ;
  assign n1292 = ~n1290 & n1291 ;
  assign n1293 = ( x724 & x725 ) | ( x724 & x726 ) | ( x725 & x726 ) ;
  assign n1294 = ( ~x724 & x725 ) | ( ~x724 & x726 ) | ( x725 & x726 ) ;
  assign n1295 = ( x724 & ~n1293 ) | ( x724 & n1294 ) | ( ~n1293 & n1294 ) ;
  assign n1296 = ( x721 & x722 ) | ( x721 & x723 ) | ( x722 & x723 ) ;
  assign n1297 = ( ~x721 & x722 ) | ( ~x721 & x723 ) | ( x722 & x723 ) ;
  assign n1298 = ( x721 & ~n1296 ) | ( x721 & n1297 ) | ( ~n1296 & n1297 ) ;
  assign n1299 = ( n1292 & n1295 ) | ( n1292 & n1298 ) | ( n1295 & n1298 ) ;
  assign n1300 = ( ~n1292 & n1295 ) | ( ~n1292 & n1298 ) | ( n1295 & n1298 ) ;
  assign n1301 = ( n1292 & ~n1299 ) | ( n1292 & n1300 ) | ( ~n1299 & n1300 ) ;
  assign n1302 = ( x709 & x710 ) | ( x709 & x711 ) | ( x710 & x711 ) ;
  assign n1303 = ( ~x709 & x710 ) | ( ~x709 & x711 ) | ( x710 & x711 ) ;
  assign n1304 = ( x709 & ~n1302 ) | ( x709 & n1303 ) | ( ~n1302 & n1303 ) ;
  assign n1305 = ( x712 & x713 ) | ( x712 & x714 ) | ( x713 & x714 ) ;
  assign n1306 = ( ~x712 & x713 ) | ( ~x712 & x714 ) | ( x713 & x714 ) ;
  assign n1307 = ( x712 & ~n1305 ) | ( x712 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1308 = ( x706 & x707 ) | ( x706 & x708 ) | ( x707 & x708 ) ;
  assign n1309 = ( ~x706 & x707 ) | ( ~x706 & x708 ) | ( x707 & x708 ) ;
  assign n1310 = ( x706 & ~n1308 ) | ( x706 & n1309 ) | ( ~n1308 & n1309 ) ;
  assign n1311 = ( x703 & x704 ) | ( x703 & x705 ) | ( x704 & x705 ) ;
  assign n1312 = ( ~x703 & x704 ) | ( ~x703 & x705 ) | ( x704 & x705 ) ;
  assign n1313 = ( x703 & ~n1311 ) | ( x703 & n1312 ) | ( ~n1311 & n1312 ) ;
  assign n1314 = n1310 & n1313 ;
  assign n1315 = n1310 | n1313 ;
  assign n1316 = ~n1314 & n1315 ;
  assign n1317 = ( n1304 & n1307 ) | ( n1304 & n1316 ) | ( n1307 & n1316 ) ;
  assign n1318 = ( ~n1304 & n1307 ) | ( ~n1304 & n1316 ) | ( n1307 & n1316 ) ;
  assign n1319 = ( n1304 & ~n1317 ) | ( n1304 & n1318 ) | ( ~n1317 & n1318 ) ;
  assign n1320 = n1301 & n1319 ;
  assign n1321 = n1301 | n1319 ;
  assign n1322 = ~n1320 & n1321 ;
  assign n1323 = n1283 & n1322 ;
  assign n1324 = n1283 | n1322 ;
  assign n1325 = ~n1323 & n1324 ;
  assign n1326 = n1244 & n1325 ;
  assign n1327 = n1244 | n1325 ;
  assign n1328 = ~n1326 & n1327 ;
  assign n1329 = n1163 & n1328 ;
  assign n1330 = ( n1002 & n1005 ) | ( n1002 & n1008 ) | ( n1005 & n1008 ) ;
  assign n1331 = ( ~n1002 & n1005 ) | ( ~n1002 & n1008 ) | ( n1005 & n1008 ) ;
  assign n1332 = ( n1002 & ~n1330 ) | ( n1002 & n1331 ) | ( ~n1330 & n1331 ) ;
  assign n1333 = n1011 & n1014 ;
  assign n1334 = n1011 | n1014 ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1336 = ( n1017 & n1332 ) | ( n1017 & n1335 ) | ( n1332 & n1335 ) ;
  assign n1337 = ( ~n1017 & n1332 ) | ( ~n1017 & n1335 ) | ( n1332 & n1335 ) ;
  assign n1338 = ( n1017 & ~n1336 ) | ( n1017 & n1337 ) | ( ~n1336 & n1337 ) ;
  assign n1339 = n1022 & n1025 ;
  assign n1340 = n1020 & n1023 ;
  assign n1341 = n1020 | n1023 ;
  assign n1342 = ~n1340 & n1341 ;
  assign n1343 = ~n1339 & n1342 ;
  assign n1344 = ( n1026 & n1029 ) | ( n1026 & n1032 ) | ( n1029 & n1032 ) ;
  assign n1345 = ( ~n1026 & n1029 ) | ( ~n1026 & n1032 ) | ( n1029 & n1032 ) ;
  assign n1346 = ( n1026 & ~n1344 ) | ( n1026 & n1345 ) | ( ~n1344 & n1345 ) ;
  assign n1347 = ( n1035 & ~n1342 ) | ( n1035 & n1343 ) | ( ~n1342 & n1343 ) ;
  assign n1348 = ( n1343 & n1346 ) | ( n1343 & n1347 ) | ( n1346 & n1347 ) ;
  assign n1349 = ( n1035 & ~n1342 ) | ( n1035 & n1346 ) | ( ~n1342 & n1346 ) ;
  assign n1350 = ( n1343 & ~n1348 ) | ( n1343 & n1349 ) | ( ~n1348 & n1349 ) ;
  assign n1351 = ( n1038 & n1338 ) | ( n1038 & n1350 ) | ( n1338 & n1350 ) ;
  assign n1352 = ( ~n1038 & n1338 ) | ( ~n1038 & n1350 ) | ( n1338 & n1350 ) ;
  assign n1353 = ( n1038 & ~n1351 ) | ( n1038 & n1352 ) | ( ~n1351 & n1352 ) ;
  assign n1354 = ( n1041 & n1044 ) | ( n1041 & n1047 ) | ( n1044 & n1047 ) ;
  assign n1355 = ( ~n1041 & n1044 ) | ( ~n1041 & n1047 ) | ( n1044 & n1047 ) ;
  assign n1356 = ( n1041 & ~n1354 ) | ( n1041 & n1355 ) | ( ~n1354 & n1355 ) ;
  assign n1357 = n1050 & n1053 ;
  assign n1358 = n1050 | n1053 ;
  assign n1359 = ~n1357 & n1358 ;
  assign n1360 = ( n1056 & n1356 ) | ( n1056 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1361 = ( ~n1056 & n1356 ) | ( ~n1056 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1362 = ( n1056 & ~n1360 ) | ( n1056 & n1361 ) | ( ~n1360 & n1361 ) ;
  assign n1363 = ( n1059 & n1062 ) | ( n1059 & n1065 ) | ( n1062 & n1065 ) ;
  assign n1364 = ( ~n1059 & n1062 ) | ( ~n1059 & n1065 ) | ( n1062 & n1065 ) ;
  assign n1365 = ( n1059 & ~n1363 ) | ( n1059 & n1364 ) | ( ~n1363 & n1364 ) ;
  assign n1366 = n1068 & n1071 ;
  assign n1367 = n1068 | n1071 ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = ( n1074 & n1365 ) | ( n1074 & n1368 ) | ( n1365 & n1368 ) ;
  assign n1370 = ( n1074 & ~n1365 ) | ( n1074 & n1368 ) | ( ~n1365 & n1368 ) ;
  assign n1371 = ( n1365 & ~n1369 ) | ( n1365 & n1370 ) | ( ~n1369 & n1370 ) ;
  assign n1372 = ( n1077 & n1362 ) | ( n1077 & n1371 ) | ( n1362 & n1371 ) ;
  assign n1373 = ( n1077 & ~n1362 ) | ( n1077 & n1371 ) | ( ~n1362 & n1371 ) ;
  assign n1374 = ( n1362 & ~n1372 ) | ( n1362 & n1373 ) | ( ~n1372 & n1373 ) ;
  assign n1375 = n1353 | n1374 ;
  assign n1376 = n1353 & n1374 ;
  assign n1377 = n1375 & ~n1376 ;
  assign n1378 = ( n1125 & n1128 ) | ( n1125 & n1131 ) | ( n1128 & n1131 ) ;
  assign n1379 = ( ~n1125 & n1128 ) | ( ~n1125 & n1131 ) | ( n1128 & n1131 ) ;
  assign n1380 = ( n1125 & ~n1378 ) | ( n1125 & n1379 ) | ( ~n1378 & n1379 ) ;
  assign n1381 = n1120 & n1123 ;
  assign n1382 = n1120 | n1123 ;
  assign n1383 = ~n1381 & n1382 ;
  assign n1384 = ( n1134 & n1380 ) | ( n1134 & n1383 ) | ( n1380 & n1383 ) ;
  assign n1385 = ( ~n1134 & n1380 ) | ( ~n1134 & n1383 ) | ( n1380 & n1383 ) ;
  assign n1386 = ( n1134 & ~n1384 ) | ( n1134 & n1385 ) | ( ~n1384 & n1385 ) ;
  assign n1387 = ( n1137 & n1140 ) | ( n1137 & n1143 ) | ( n1140 & n1143 ) ;
  assign n1388 = ( ~n1137 & n1140 ) | ( ~n1137 & n1143 ) | ( n1140 & n1143 ) ;
  assign n1389 = ( n1137 & ~n1387 ) | ( n1137 & n1388 ) | ( ~n1387 & n1388 ) ;
  assign n1390 = n1146 & n1149 ;
  assign n1391 = n1146 | n1149 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = ( n1152 & n1389 ) | ( n1152 & n1392 ) | ( n1389 & n1392 ) ;
  assign n1394 = ( ~n1152 & n1389 ) | ( ~n1152 & n1392 ) | ( n1389 & n1392 ) ;
  assign n1395 = ( n1152 & ~n1393 ) | ( n1152 & n1394 ) | ( ~n1393 & n1394 ) ;
  assign n1396 = ( n1155 & n1386 ) | ( n1155 & n1395 ) | ( n1386 & n1395 ) ;
  assign n1397 = ( ~n1155 & n1386 ) | ( ~n1155 & n1395 ) | ( n1386 & n1395 ) ;
  assign n1398 = ( n1155 & ~n1396 ) | ( n1155 & n1397 ) | ( ~n1396 & n1397 ) ;
  assign n1399 = ( n1080 & n1083 ) | ( n1080 & n1086 ) | ( n1083 & n1086 ) ;
  assign n1400 = ( ~n1080 & n1083 ) | ( ~n1080 & n1086 ) | ( n1083 & n1086 ) ;
  assign n1401 = ( n1080 & ~n1399 ) | ( n1080 & n1400 ) | ( ~n1399 & n1400 ) ;
  assign n1402 = n1095 & n1401 ;
  assign n1403 = n1095 | n1401 ;
  assign n1404 = ~n1402 & n1403 ;
  assign n1405 = ( n1090 & n1093 ) | ( n1090 & n1404 ) | ( n1093 & n1404 ) ;
  assign n1406 = ( n1090 & n1093 ) | ( n1090 & ~n1404 ) | ( n1093 & ~n1404 ) ;
  assign n1407 = ( n1404 & ~n1405 ) | ( n1404 & n1406 ) | ( ~n1405 & n1406 ) ;
  assign n1408 = n1100 & n1103 ;
  assign n1409 = n1098 & n1101 ;
  assign n1410 = n1098 | n1101 ;
  assign n1411 = ~n1409 & n1410 ;
  assign n1412 = ~n1408 & n1411 ;
  assign n1413 = ( n1104 & n1107 ) | ( n1104 & n1110 ) | ( n1107 & n1110 ) ;
  assign n1414 = ( ~n1104 & n1107 ) | ( ~n1104 & n1110 ) | ( n1107 & n1110 ) ;
  assign n1415 = ( n1104 & ~n1413 ) | ( n1104 & n1414 ) | ( ~n1413 & n1414 ) ;
  assign n1416 = ( n1113 & ~n1411 ) | ( n1113 & n1412 ) | ( ~n1411 & n1412 ) ;
  assign n1417 = ( n1412 & n1415 ) | ( n1412 & n1416 ) | ( n1415 & n1416 ) ;
  assign n1418 = ( n1113 & ~n1411 ) | ( n1113 & n1415 ) | ( ~n1411 & n1415 ) ;
  assign n1419 = ( n1412 & ~n1417 ) | ( n1412 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = ( n1116 & n1407 ) | ( n1116 & n1419 ) | ( n1407 & n1419 ) ;
  assign n1421 = ( n1116 & ~n1407 ) | ( n1116 & n1419 ) | ( ~n1407 & n1419 ) ;
  assign n1422 = ( n1407 & ~n1420 ) | ( n1407 & n1421 ) | ( ~n1420 & n1421 ) ;
  assign n1423 = ( n1158 & n1398 ) | ( n1158 & n1422 ) | ( n1398 & n1422 ) ;
  assign n1424 = ( ~n1158 & n1398 ) | ( ~n1158 & n1422 ) | ( n1398 & n1422 ) ;
  assign n1425 = ( n1158 & ~n1423 ) | ( n1158 & n1424 ) | ( ~n1423 & n1424 ) ;
  assign n1426 = ( n1161 & n1377 ) | ( n1161 & n1425 ) | ( n1377 & n1425 ) ;
  assign n1427 = ( n1161 & ~n1377 ) | ( n1161 & n1425 ) | ( ~n1377 & n1425 ) ;
  assign n1428 = ( n1377 & ~n1426 ) | ( n1377 & n1427 ) | ( ~n1426 & n1427 ) ;
  assign n1429 = ( n1263 & n1266 ) | ( n1263 & n1269 ) | ( n1266 & n1269 ) ;
  assign n1430 = ( ~n1263 & n1266 ) | ( ~n1263 & n1269 ) | ( n1266 & n1269 ) ;
  assign n1431 = ( n1263 & ~n1429 ) | ( n1263 & n1430 ) | ( ~n1429 & n1430 ) ;
  assign n1432 = n1273 & n1276 ;
  assign n1433 = n1273 | n1276 ;
  assign n1434 = ~n1432 & n1433 ;
  assign n1435 = ( n1278 & n1431 ) | ( n1278 & n1434 ) | ( n1431 & n1434 ) ;
  assign n1436 = ( n1278 & ~n1431 ) | ( n1278 & n1434 ) | ( ~n1431 & n1434 ) ;
  assign n1437 = ( n1431 & ~n1435 ) | ( n1431 & n1436 ) | ( ~n1435 & n1436 ) ;
  assign n1438 = ( n1245 & n1248 ) | ( n1245 & n1251 ) | ( n1248 & n1251 ) ;
  assign n1439 = ( ~n1245 & n1248 ) | ( ~n1245 & n1251 ) | ( n1248 & n1251 ) ;
  assign n1440 = ( n1245 & ~n1438 ) | ( n1245 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1441 = n1254 & n1257 ;
  assign n1442 = n1254 | n1257 ;
  assign n1443 = ~n1441 & n1442 ;
  assign n1444 = ( n1260 & n1440 ) | ( n1260 & n1443 ) | ( n1440 & n1443 ) ;
  assign n1445 = ( ~n1260 & n1440 ) | ( ~n1260 & n1443 ) | ( n1440 & n1443 ) ;
  assign n1446 = ( n1260 & ~n1444 ) | ( n1260 & n1445 ) | ( ~n1444 & n1445 ) ;
  assign n1447 = ( n1281 & n1437 ) | ( n1281 & n1446 ) | ( n1437 & n1446 ) ;
  assign n1448 = ( n1281 & ~n1437 ) | ( n1281 & n1446 ) | ( ~n1437 & n1446 ) ;
  assign n1449 = ( n1437 & ~n1447 ) | ( n1437 & n1448 ) | ( ~n1447 & n1448 ) ;
  assign n1450 = ( n1284 & n1287 ) | ( n1284 & n1290 ) | ( n1287 & n1290 ) ;
  assign n1451 = ( ~n1284 & n1287 ) | ( ~n1284 & n1290 ) | ( n1287 & n1290 ) ;
  assign n1452 = ( n1284 & ~n1450 ) | ( n1284 & n1451 ) | ( ~n1450 & n1451 ) ;
  assign n1453 = n1293 & n1296 ;
  assign n1454 = n1293 | n1296 ;
  assign n1455 = ~n1453 & n1454 ;
  assign n1456 = ( n1299 & n1452 ) | ( n1299 & n1455 ) | ( n1452 & n1455 ) ;
  assign n1457 = ( ~n1299 & n1452 ) | ( ~n1299 & n1455 ) | ( n1452 & n1455 ) ;
  assign n1458 = ( n1299 & ~n1456 ) | ( n1299 & n1457 ) | ( ~n1456 & n1457 ) ;
  assign n1459 = ( n1308 & n1311 ) | ( n1308 & n1314 ) | ( n1311 & n1314 ) ;
  assign n1460 = ( ~n1308 & n1311 ) | ( ~n1308 & n1314 ) | ( n1311 & n1314 ) ;
  assign n1461 = ( n1308 & ~n1459 ) | ( n1308 & n1460 ) | ( ~n1459 & n1460 ) ;
  assign n1462 = n1302 & n1305 ;
  assign n1463 = n1302 | n1305 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = ( n1317 & n1461 ) | ( n1317 & n1464 ) | ( n1461 & n1464 ) ;
  assign n1466 = ( ~n1317 & n1461 ) | ( ~n1317 & n1464 ) | ( n1461 & n1464 ) ;
  assign n1467 = ( n1317 & ~n1465 ) | ( n1317 & n1466 ) | ( ~n1465 & n1466 ) ;
  assign n1468 = ( n1320 & n1458 ) | ( n1320 & n1467 ) | ( n1458 & n1467 ) ;
  assign n1469 = ( n1320 & ~n1458 ) | ( n1320 & n1467 ) | ( ~n1458 & n1467 ) ;
  assign n1470 = ( n1458 & ~n1468 ) | ( n1458 & n1469 ) | ( ~n1468 & n1469 ) ;
  assign n1471 = ( n1323 & n1449 ) | ( n1323 & n1470 ) | ( n1449 & n1470 ) ;
  assign n1472 = ( ~n1323 & n1449 ) | ( ~n1323 & n1470 ) | ( n1449 & n1470 ) ;
  assign n1473 = ( n1323 & ~n1471 ) | ( n1323 & n1472 ) | ( ~n1471 & n1472 ) ;
  assign n1474 = ( n1170 & n1173 ) | ( n1170 & n1176 ) | ( n1173 & n1176 ) ;
  assign n1475 = ( ~n1170 & n1173 ) | ( ~n1170 & n1176 ) | ( n1173 & n1176 ) ;
  assign n1476 = ( n1170 & ~n1474 ) | ( n1170 & n1475 ) | ( ~n1474 & n1475 ) ;
  assign n1477 = n1165 & n1168 ;
  assign n1478 = n1165 | n1168 ;
  assign n1479 = ~n1477 & n1478 ;
  assign n1480 = ( n1179 & n1476 ) | ( n1179 & n1479 ) | ( n1476 & n1479 ) ;
  assign n1481 = ( ~n1179 & n1476 ) | ( ~n1179 & n1479 ) | ( n1476 & n1479 ) ;
  assign n1482 = ( n1179 & ~n1480 ) | ( n1179 & n1481 ) | ( ~n1480 & n1481 ) ;
  assign n1483 = ( n1182 & n1185 ) | ( n1182 & n1188 ) | ( n1185 & n1188 ) ;
  assign n1484 = ( ~n1182 & n1185 ) | ( ~n1182 & n1188 ) | ( n1185 & n1188 ) ;
  assign n1485 = ( n1182 & ~n1483 ) | ( n1182 & n1484 ) | ( ~n1483 & n1484 ) ;
  assign n1486 = n1191 & n1194 ;
  assign n1487 = n1191 | n1194 ;
  assign n1488 = ~n1486 & n1487 ;
  assign n1489 = ( n1197 & n1485 ) | ( n1197 & n1488 ) | ( n1485 & n1488 ) ;
  assign n1490 = ( ~n1197 & n1485 ) | ( ~n1197 & n1488 ) | ( n1485 & n1488 ) ;
  assign n1491 = ( n1197 & ~n1489 ) | ( n1197 & n1490 ) | ( ~n1489 & n1490 ) ;
  assign n1492 = ( n1200 & n1482 ) | ( n1200 & n1491 ) | ( n1482 & n1491 ) ;
  assign n1493 = ( ~n1200 & n1482 ) | ( ~n1200 & n1491 ) | ( n1482 & n1491 ) ;
  assign n1494 = ( n1200 & ~n1492 ) | ( n1200 & n1493 ) | ( ~n1492 & n1493 ) ;
  assign n1495 = ( n1221 & n1224 ) | ( n1221 & n1227 ) | ( n1224 & n1227 ) ;
  assign n1496 = ( ~n1221 & n1224 ) | ( ~n1221 & n1227 ) | ( n1224 & n1227 ) ;
  assign n1497 = ( n1221 & ~n1495 ) | ( n1221 & n1496 ) | ( ~n1495 & n1496 ) ;
  assign n1498 = n1236 & n1497 ;
  assign n1499 = n1236 | n1497 ;
  assign n1500 = ~n1498 & n1499 ;
  assign n1501 = ( n1231 & n1234 ) | ( n1231 & n1500 ) | ( n1234 & n1500 ) ;
  assign n1502 = ( n1231 & n1234 ) | ( n1231 & ~n1500 ) | ( n1234 & ~n1500 ) ;
  assign n1503 = ( n1500 & ~n1501 ) | ( n1500 & n1502 ) | ( ~n1501 & n1502 ) ;
  assign n1504 = ( n1209 & n1212 ) | ( n1209 & n1215 ) | ( n1212 & n1215 ) ;
  assign n1505 = ( ~n1209 & n1212 ) | ( ~n1209 & n1215 ) | ( n1212 & n1215 ) ;
  assign n1506 = ( n1209 & ~n1504 ) | ( n1209 & n1505 ) | ( ~n1504 & n1505 ) ;
  assign n1507 = n1204 & n1207 ;
  assign n1508 = n1204 | n1207 ;
  assign n1509 = ~n1507 & n1508 ;
  assign n1510 = ( n1218 & n1506 ) | ( n1218 & n1509 ) | ( n1506 & n1509 ) ;
  assign n1511 = ( ~n1218 & n1506 ) | ( ~n1218 & n1509 ) | ( n1506 & n1509 ) ;
  assign n1512 = ( n1218 & ~n1510 ) | ( n1218 & n1511 ) | ( ~n1510 & n1511 ) ;
  assign n1513 = ( n1239 & n1503 ) | ( n1239 & n1512 ) | ( n1503 & n1512 ) ;
  assign n1514 = ( n1239 & ~n1503 ) | ( n1239 & n1512 ) | ( ~n1503 & n1512 ) ;
  assign n1515 = ( n1503 & ~n1513 ) | ( n1503 & n1514 ) | ( ~n1513 & n1514 ) ;
  assign n1516 = ( n1242 & n1494 ) | ( n1242 & n1515 ) | ( n1494 & n1515 ) ;
  assign n1517 = ( n1242 & ~n1494 ) | ( n1242 & n1515 ) | ( ~n1494 & n1515 ) ;
  assign n1518 = ( n1494 & ~n1516 ) | ( n1494 & n1517 ) | ( ~n1516 & n1517 ) ;
  assign n1519 = ( n1326 & n1473 ) | ( n1326 & n1518 ) | ( n1473 & n1518 ) ;
  assign n1520 = ( n1326 & ~n1473 ) | ( n1326 & n1518 ) | ( ~n1473 & n1518 ) ;
  assign n1521 = ( n1473 & ~n1519 ) | ( n1473 & n1520 ) | ( ~n1519 & n1520 ) ;
  assign n1522 = ( n1329 & n1428 ) | ( n1329 & n1521 ) | ( n1428 & n1521 ) ;
  assign n1523 = n1040 & n1079 ;
  assign n1524 = n1377 & n1523 ;
  assign n1525 = n1426 & ~n1524 ;
  assign n1526 = ( n1020 & n1023 ) | ( n1020 & n1339 ) | ( n1023 & n1339 ) ;
  assign n1527 = ( n1344 & n1348 ) | ( n1344 & n1526 ) | ( n1348 & n1526 ) ;
  assign n1528 = ( ~n1344 & n1348 ) | ( ~n1344 & n1526 ) | ( n1348 & n1526 ) ;
  assign n1529 = ( n1344 & ~n1527 ) | ( n1344 & n1528 ) | ( ~n1527 & n1528 ) ;
  assign n1530 = ( n1330 & n1333 ) | ( n1330 & n1336 ) | ( n1333 & n1336 ) ;
  assign n1531 = ( n1330 & n1333 ) | ( n1330 & ~n1336 ) | ( n1333 & ~n1336 ) ;
  assign n1532 = ( n1336 & ~n1530 ) | ( n1336 & n1531 ) | ( ~n1530 & n1531 ) ;
  assign n1533 = ( n1351 & n1529 ) | ( n1351 & n1532 ) | ( n1529 & n1532 ) ;
  assign n1534 = ( ~n1351 & n1529 ) | ( ~n1351 & n1532 ) | ( n1529 & n1532 ) ;
  assign n1535 = ( n1351 & ~n1533 ) | ( n1351 & n1534 ) | ( ~n1533 & n1534 ) ;
  assign n1536 = ( n1353 & n1374 ) | ( n1353 & n1523 ) | ( n1374 & n1523 ) ;
  assign n1537 = ( n1354 & n1357 ) | ( n1354 & n1360 ) | ( n1357 & n1360 ) ;
  assign n1538 = ( n1354 & n1357 ) | ( n1354 & ~n1360 ) | ( n1357 & ~n1360 ) ;
  assign n1539 = ( n1360 & ~n1537 ) | ( n1360 & n1538 ) | ( ~n1537 & n1538 ) ;
  assign n1540 = ( n1363 & n1366 ) | ( n1363 & n1369 ) | ( n1366 & n1369 ) ;
  assign n1541 = ( n1363 & n1366 ) | ( n1363 & ~n1369 ) | ( n1366 & ~n1369 ) ;
  assign n1542 = ( n1369 & ~n1540 ) | ( n1369 & n1541 ) | ( ~n1540 & n1541 ) ;
  assign n1543 = ( n1372 & n1539 ) | ( n1372 & n1542 ) | ( n1539 & n1542 ) ;
  assign n1544 = ( ~n1372 & n1539 ) | ( ~n1372 & n1542 ) | ( n1539 & n1542 ) ;
  assign n1545 = ( n1372 & ~n1543 ) | ( n1372 & n1544 ) | ( ~n1543 & n1544 ) ;
  assign n1546 = ( n1535 & n1536 ) | ( n1535 & n1545 ) | ( n1536 & n1545 ) ;
  assign n1547 = ( ~n1535 & n1536 ) | ( ~n1535 & n1545 ) | ( n1536 & n1545 ) ;
  assign n1548 = ( n1535 & ~n1546 ) | ( n1535 & n1547 ) | ( ~n1546 & n1547 ) ;
  assign n1549 = ( n1098 & n1101 ) | ( n1098 & n1408 ) | ( n1101 & n1408 ) ;
  assign n1550 = ( n1413 & n1417 ) | ( n1413 & n1549 ) | ( n1417 & n1549 ) ;
  assign n1551 = ( ~n1413 & n1417 ) | ( ~n1413 & n1549 ) | ( n1417 & n1549 ) ;
  assign n1552 = ( n1413 & ~n1550 ) | ( n1413 & n1551 ) | ( ~n1550 & n1551 ) ;
  assign n1553 = ( n1399 & n1402 ) | ( n1399 & n1405 ) | ( n1402 & n1405 ) ;
  assign n1554 = ( n1399 & n1402 ) | ( n1399 & ~n1405 ) | ( n1402 & ~n1405 ) ;
  assign n1555 = ( n1405 & ~n1553 ) | ( n1405 & n1554 ) | ( ~n1553 & n1554 ) ;
  assign n1556 = ( n1420 & n1552 ) | ( n1420 & n1555 ) | ( n1552 & n1555 ) ;
  assign n1557 = ( ~n1420 & n1552 ) | ( ~n1420 & n1555 ) | ( n1552 & n1555 ) ;
  assign n1558 = ( n1420 & ~n1556 ) | ( n1420 & n1557 ) | ( ~n1556 & n1557 ) ;
  assign n1559 = ( n1387 & n1390 ) | ( n1387 & n1393 ) | ( n1390 & n1393 ) ;
  assign n1560 = ( n1387 & n1390 ) | ( n1387 & ~n1393 ) | ( n1390 & ~n1393 ) ;
  assign n1561 = ( n1393 & ~n1559 ) | ( n1393 & n1560 ) | ( ~n1559 & n1560 ) ;
  assign n1562 = n1133 & ~n1136 ;
  assign n1563 = ( n1380 & ~n1386 ) | ( n1380 & n1562 ) | ( ~n1386 & n1562 ) ;
  assign n1564 = n1121 & n1124 ;
  assign n1565 = ( n1120 & n1123 ) | ( n1120 & n1564 ) | ( n1123 & n1564 ) ;
  assign n1566 = ( n1378 & n1563 ) | ( n1378 & n1565 ) | ( n1563 & n1565 ) ;
  assign n1567 = ( n1378 & ~n1563 ) | ( n1378 & n1565 ) | ( ~n1563 & n1565 ) ;
  assign n1568 = ( n1563 & ~n1566 ) | ( n1563 & n1567 ) | ( ~n1566 & n1567 ) ;
  assign n1569 = ( n1396 & n1561 ) | ( n1396 & n1568 ) | ( n1561 & n1568 ) ;
  assign n1570 = ( ~n1396 & n1561 ) | ( ~n1396 & n1568 ) | ( n1561 & n1568 ) ;
  assign n1571 = ( n1396 & ~n1569 ) | ( n1396 & n1570 ) | ( ~n1569 & n1570 ) ;
  assign n1572 = ( n1423 & n1558 ) | ( n1423 & n1571 ) | ( n1558 & n1571 ) ;
  assign n1573 = ( ~n1423 & n1558 ) | ( ~n1423 & n1571 ) | ( n1558 & n1571 ) ;
  assign n1574 = ( n1423 & ~n1572 ) | ( n1423 & n1573 ) | ( ~n1572 & n1573 ) ;
  assign n1575 = ( n1525 & n1548 ) | ( n1525 & n1574 ) | ( n1548 & n1574 ) ;
  assign n1576 = ( ~n1525 & n1548 ) | ( ~n1525 & n1574 ) | ( n1548 & n1574 ) ;
  assign n1577 = ( n1525 & ~n1575 ) | ( n1525 & n1576 ) | ( ~n1575 & n1576 ) ;
  assign n1578 = ( n1438 & n1441 ) | ( n1438 & n1444 ) | ( n1441 & n1444 ) ;
  assign n1579 = ( n1438 & n1441 ) | ( n1438 & ~n1444 ) | ( n1441 & ~n1444 ) ;
  assign n1580 = ( n1444 & ~n1578 ) | ( n1444 & n1579 ) | ( ~n1578 & n1579 ) ;
  assign n1581 = n1279 & ~n1436 ;
  assign n1582 = ( ~n1279 & n1435 ) | ( ~n1279 & n1581 ) | ( n1435 & n1581 ) ;
  assign n1583 = n1274 & n1277 ;
  assign n1584 = ( n1273 & n1276 ) | ( n1273 & n1583 ) | ( n1276 & n1583 ) ;
  assign n1585 = ( n1429 & n1582 ) | ( n1429 & n1584 ) | ( n1582 & n1584 ) ;
  assign n1586 = ( n1429 & ~n1582 ) | ( n1429 & n1584 ) | ( ~n1582 & n1584 ) ;
  assign n1587 = ( n1582 & ~n1585 ) | ( n1582 & n1586 ) | ( ~n1585 & n1586 ) ;
  assign n1588 = ( n1447 & n1580 ) | ( n1447 & n1587 ) | ( n1580 & n1587 ) ;
  assign n1589 = ( ~n1447 & n1580 ) | ( ~n1447 & n1587 ) | ( n1580 & n1587 ) ;
  assign n1590 = ( n1447 & ~n1588 ) | ( n1447 & n1589 ) | ( ~n1588 & n1589 ) ;
  assign n1591 = n1304 & n1307 ;
  assign n1592 = n1464 & ~n1591 ;
  assign n1593 = ( n1461 & ~n1467 ) | ( n1461 & n1592 ) | ( ~n1467 & n1592 ) ;
  assign n1594 = ( n1302 & n1305 ) | ( n1302 & n1591 ) | ( n1305 & n1591 ) ;
  assign n1595 = ( n1459 & n1593 ) | ( n1459 & n1594 ) | ( n1593 & n1594 ) ;
  assign n1596 = ( n1459 & ~n1593 ) | ( n1459 & n1594 ) | ( ~n1593 & n1594 ) ;
  assign n1597 = ( n1593 & ~n1595 ) | ( n1593 & n1596 ) | ( ~n1595 & n1596 ) ;
  assign n1598 = ( n1450 & n1453 ) | ( n1450 & n1456 ) | ( n1453 & n1456 ) ;
  assign n1599 = ( n1450 & n1453 ) | ( n1450 & ~n1456 ) | ( n1453 & ~n1456 ) ;
  assign n1600 = ( n1456 & ~n1598 ) | ( n1456 & n1599 ) | ( ~n1598 & n1599 ) ;
  assign n1601 = ( n1468 & n1597 ) | ( n1468 & n1600 ) | ( n1597 & n1600 ) ;
  assign n1602 = ( n1468 & ~n1597 ) | ( n1468 & n1600 ) | ( ~n1597 & n1600 ) ;
  assign n1603 = ( n1597 & ~n1601 ) | ( n1597 & n1602 ) | ( ~n1601 & n1602 ) ;
  assign n1604 = ( n1471 & n1590 ) | ( n1471 & n1603 ) | ( n1590 & n1603 ) ;
  assign n1605 = ( ~n1471 & n1590 ) | ( ~n1471 & n1603 ) | ( n1590 & n1603 ) ;
  assign n1606 = ( n1471 & ~n1604 ) | ( n1471 & n1605 ) | ( ~n1604 & n1605 ) ;
  assign n1607 = n1178 & ~n1181 ;
  assign n1608 = ( n1476 & ~n1482 ) | ( n1476 & n1607 ) | ( ~n1482 & n1607 ) ;
  assign n1609 = n1166 & n1169 ;
  assign n1610 = ( n1165 & n1168 ) | ( n1165 & n1609 ) | ( n1168 & n1609 ) ;
  assign n1611 = ( n1474 & n1608 ) | ( n1474 & n1610 ) | ( n1608 & n1610 ) ;
  assign n1612 = ( n1474 & ~n1608 ) | ( n1474 & n1610 ) | ( ~n1608 & n1610 ) ;
  assign n1613 = ( n1608 & ~n1611 ) | ( n1608 & n1612 ) | ( ~n1611 & n1612 ) ;
  assign n1614 = ( n1483 & n1486 ) | ( n1483 & n1489 ) | ( n1486 & n1489 ) ;
  assign n1615 = ( n1483 & n1486 ) | ( n1483 & ~n1489 ) | ( n1486 & ~n1489 ) ;
  assign n1616 = ( n1489 & ~n1614 ) | ( n1489 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = ( n1492 & n1613 ) | ( n1492 & n1616 ) | ( n1613 & n1616 ) ;
  assign n1618 = ( ~n1492 & n1613 ) | ( ~n1492 & n1616 ) | ( n1613 & n1616 ) ;
  assign n1619 = ( n1492 & ~n1617 ) | ( n1492 & n1618 ) | ( ~n1617 & n1618 ) ;
  assign n1620 = n1217 & ~n1220 ;
  assign n1621 = ( n1506 & ~n1512 ) | ( n1506 & n1620 ) | ( ~n1512 & n1620 ) ;
  assign n1622 = n1205 & n1208 ;
  assign n1623 = ( n1204 & n1207 ) | ( n1204 & n1622 ) | ( n1207 & n1622 ) ;
  assign n1624 = ( n1504 & n1621 ) | ( n1504 & n1623 ) | ( n1621 & n1623 ) ;
  assign n1625 = ( n1504 & ~n1621 ) | ( n1504 & n1623 ) | ( ~n1621 & n1623 ) ;
  assign n1626 = ( n1621 & ~n1624 ) | ( n1621 & n1625 ) | ( ~n1624 & n1625 ) ;
  assign n1627 = ( n1495 & n1498 ) | ( n1495 & n1501 ) | ( n1498 & n1501 ) ;
  assign n1628 = ( n1495 & n1498 ) | ( n1495 & ~n1501 ) | ( n1498 & ~n1501 ) ;
  assign n1629 = ( n1501 & ~n1627 ) | ( n1501 & n1628 ) | ( ~n1627 & n1628 ) ;
  assign n1630 = ( n1513 & n1626 ) | ( n1513 & n1629 ) | ( n1626 & n1629 ) ;
  assign n1631 = ( n1513 & ~n1626 ) | ( n1513 & n1629 ) | ( ~n1626 & n1629 ) ;
  assign n1632 = ( n1626 & ~n1630 ) | ( n1626 & n1631 ) | ( ~n1630 & n1631 ) ;
  assign n1633 = ( n1516 & n1619 ) | ( n1516 & n1632 ) | ( n1619 & n1632 ) ;
  assign n1634 = ( ~n1516 & n1619 ) | ( ~n1516 & n1632 ) | ( n1619 & n1632 ) ;
  assign n1635 = ( n1516 & ~n1633 ) | ( n1516 & n1634 ) | ( ~n1633 & n1634 ) ;
  assign n1636 = ( n1519 & n1606 ) | ( n1519 & n1635 ) | ( n1606 & n1635 ) ;
  assign n1637 = ( ~n1519 & n1606 ) | ( ~n1519 & n1635 ) | ( n1606 & n1635 ) ;
  assign n1638 = ( n1519 & ~n1636 ) | ( n1519 & n1637 ) | ( ~n1636 & n1637 ) ;
  assign n1639 = ( n1522 & n1577 ) | ( n1522 & n1638 ) | ( n1577 & n1638 ) ;
  assign n1640 = ( n1550 & n1553 ) | ( n1550 & n1556 ) | ( n1553 & n1556 ) ;
  assign n1641 = ( n1550 & n1553 ) | ( n1550 & ~n1556 ) | ( n1553 & ~n1556 ) ;
  assign n1642 = ( n1556 & ~n1640 ) | ( n1556 & n1641 ) | ( ~n1640 & n1641 ) ;
  assign n1643 = ( n1559 & n1566 ) | ( n1559 & n1569 ) | ( n1566 & n1569 ) ;
  assign n1644 = ( n1559 & n1566 ) | ( n1559 & ~n1569 ) | ( n1566 & ~n1569 ) ;
  assign n1645 = ( n1569 & ~n1643 ) | ( n1569 & n1644 ) | ( ~n1643 & n1644 ) ;
  assign n1646 = ( n1572 & n1642 ) | ( n1572 & n1645 ) | ( n1642 & n1645 ) ;
  assign n1647 = ( ~n1572 & n1642 ) | ( ~n1572 & n1645 ) | ( n1642 & n1645 ) ;
  assign n1648 = ( n1572 & ~n1646 ) | ( n1572 & n1647 ) | ( ~n1646 & n1647 ) ;
  assign n1649 = ( n1527 & n1530 ) | ( n1527 & n1533 ) | ( n1530 & n1533 ) ;
  assign n1650 = ( n1527 & n1530 ) | ( n1527 & ~n1533 ) | ( n1530 & ~n1533 ) ;
  assign n1651 = ( n1533 & ~n1649 ) | ( n1533 & n1650 ) | ( ~n1649 & n1650 ) ;
  assign n1652 = ( n1537 & n1540 ) | ( n1537 & n1543 ) | ( n1540 & n1543 ) ;
  assign n1653 = ( ~n1537 & n1540 ) | ( ~n1537 & n1543 ) | ( n1540 & n1543 ) ;
  assign n1654 = ( n1537 & ~n1652 ) | ( n1537 & n1653 ) | ( ~n1652 & n1653 ) ;
  assign n1655 = ( n1546 & n1651 ) | ( n1546 & n1654 ) | ( n1651 & n1654 ) ;
  assign n1656 = ( ~n1546 & n1651 ) | ( ~n1546 & n1654 ) | ( n1651 & n1654 ) ;
  assign n1657 = ( n1546 & ~n1655 ) | ( n1546 & n1656 ) | ( ~n1655 & n1656 ) ;
  assign n1658 = ( n1575 & n1648 ) | ( n1575 & n1657 ) | ( n1648 & n1657 ) ;
  assign n1659 = ( ~n1575 & n1648 ) | ( ~n1575 & n1657 ) | ( n1648 & n1657 ) ;
  assign n1660 = ( n1575 & ~n1658 ) | ( n1575 & n1659 ) | ( ~n1658 & n1659 ) ;
  assign n1661 = ( n1624 & n1627 ) | ( n1624 & n1630 ) | ( n1627 & n1630 ) ;
  assign n1662 = ( ~n1624 & n1627 ) | ( ~n1624 & n1630 ) | ( n1627 & n1630 ) ;
  assign n1663 = ( n1624 & ~n1661 ) | ( n1624 & n1662 ) | ( ~n1661 & n1662 ) ;
  assign n1664 = ( n1611 & n1614 ) | ( n1611 & n1617 ) | ( n1614 & n1617 ) ;
  assign n1665 = ( n1611 & n1614 ) | ( n1611 & ~n1617 ) | ( n1614 & ~n1617 ) ;
  assign n1666 = ( n1617 & ~n1664 ) | ( n1617 & n1665 ) | ( ~n1664 & n1665 ) ;
  assign n1667 = ( n1633 & n1663 ) | ( n1633 & n1666 ) | ( n1663 & n1666 ) ;
  assign n1668 = ( ~n1633 & n1663 ) | ( ~n1633 & n1666 ) | ( n1663 & n1666 ) ;
  assign n1669 = ( n1633 & ~n1667 ) | ( n1633 & n1668 ) | ( ~n1667 & n1668 ) ;
  assign n1670 = ( n1595 & n1598 ) | ( n1595 & n1601 ) | ( n1598 & n1601 ) ;
  assign n1671 = ( n1595 & n1598 ) | ( n1595 & ~n1601 ) | ( n1598 & ~n1601 ) ;
  assign n1672 = ( n1601 & ~n1670 ) | ( n1601 & n1671 ) | ( ~n1670 & n1671 ) ;
  assign n1673 = ( n1578 & n1585 ) | ( n1578 & n1588 ) | ( n1585 & n1588 ) ;
  assign n1674 = ( n1578 & n1585 ) | ( n1578 & ~n1588 ) | ( n1585 & ~n1588 ) ;
  assign n1675 = ( n1588 & ~n1673 ) | ( n1588 & n1674 ) | ( ~n1673 & n1674 ) ;
  assign n1676 = ( n1604 & n1672 ) | ( n1604 & n1675 ) | ( n1672 & n1675 ) ;
  assign n1677 = ( ~n1604 & n1672 ) | ( ~n1604 & n1675 ) | ( n1672 & n1675 ) ;
  assign n1678 = ( n1604 & ~n1676 ) | ( n1604 & n1677 ) | ( ~n1676 & n1677 ) ;
  assign n1679 = ( n1636 & n1669 ) | ( n1636 & n1678 ) | ( n1669 & n1678 ) ;
  assign n1680 = ( ~n1636 & n1669 ) | ( ~n1636 & n1678 ) | ( n1669 & n1678 ) ;
  assign n1681 = ( n1636 & ~n1679 ) | ( n1636 & n1680 ) | ( ~n1679 & n1680 ) ;
  assign n1682 = ( n1639 & n1660 ) | ( n1639 & n1681 ) | ( n1660 & n1681 ) ;
  assign n1683 = ( n1640 & n1643 ) | ( n1640 & n1646 ) | ( n1643 & n1646 ) ;
  assign n1684 = ( n1640 & n1643 ) | ( n1640 & ~n1646 ) | ( n1643 & ~n1646 ) ;
  assign n1685 = ( n1646 & ~n1683 ) | ( n1646 & n1684 ) | ( ~n1683 & n1684 ) ;
  assign n1686 = ( n1649 & n1652 ) | ( n1649 & n1655 ) | ( n1652 & n1655 ) ;
  assign n1687 = ( n1649 & n1652 ) | ( n1649 & ~n1655 ) | ( n1652 & ~n1655 ) ;
  assign n1688 = ( n1655 & ~n1686 ) | ( n1655 & n1687 ) | ( ~n1686 & n1687 ) ;
  assign n1689 = ( n1658 & n1685 ) | ( n1658 & n1688 ) | ( n1685 & n1688 ) ;
  assign n1690 = ( ~n1658 & n1685 ) | ( ~n1658 & n1688 ) | ( n1685 & n1688 ) ;
  assign n1691 = ( n1658 & ~n1689 ) | ( n1658 & n1690 ) | ( ~n1689 & n1690 ) ;
  assign n1692 = ( n1661 & n1664 ) | ( n1661 & n1667 ) | ( n1664 & n1667 ) ;
  assign n1693 = ( n1661 & n1664 ) | ( n1661 & ~n1667 ) | ( n1664 & ~n1667 ) ;
  assign n1694 = ( n1667 & ~n1692 ) | ( n1667 & n1693 ) | ( ~n1692 & n1693 ) ;
  assign n1695 = ( n1670 & n1673 ) | ( n1670 & n1676 ) | ( n1673 & n1676 ) ;
  assign n1696 = ( n1670 & n1673 ) | ( n1670 & ~n1676 ) | ( n1673 & ~n1676 ) ;
  assign n1697 = ( n1676 & ~n1695 ) | ( n1676 & n1696 ) | ( ~n1695 & n1696 ) ;
  assign n1698 = ( n1679 & n1694 ) | ( n1679 & n1697 ) | ( n1694 & n1697 ) ;
  assign n1699 = ( ~n1679 & n1694 ) | ( ~n1679 & n1697 ) | ( n1694 & n1697 ) ;
  assign n1700 = ( n1679 & ~n1698 ) | ( n1679 & n1699 ) | ( ~n1698 & n1699 ) ;
  assign n1701 = ( n1682 & n1691 ) | ( n1682 & n1700 ) | ( n1691 & n1700 ) ;
  assign n1702 = ( n1692 & n1695 ) | ( n1692 & n1698 ) | ( n1695 & n1698 ) ;
  assign n1703 = ( n1692 & n1695 ) | ( n1692 & ~n1698 ) | ( n1695 & ~n1698 ) ;
  assign n1704 = ( n1698 & ~n1702 ) | ( n1698 & n1703 ) | ( ~n1702 & n1703 ) ;
  assign n1705 = ( n1683 & n1686 ) | ( n1683 & n1689 ) | ( n1686 & n1689 ) ;
  assign n1706 = ( n1683 & n1686 ) | ( n1683 & ~n1689 ) | ( n1686 & ~n1689 ) ;
  assign n1707 = ( n1689 & ~n1705 ) | ( n1689 & n1706 ) | ( ~n1705 & n1706 ) ;
  assign n1708 = ( n1701 & n1704 ) | ( n1701 & n1707 ) | ( n1704 & n1707 ) ;
  assign n1709 = ( n1702 & n1705 ) | ( n1702 & n1708 ) | ( n1705 & n1708 ) ;
  assign n1710 = ( n1702 & n1705 ) | ( n1702 & ~n1708 ) | ( n1705 & ~n1708 ) ;
  assign n1711 = ( n1708 & ~n1709 ) | ( n1708 & n1710 ) | ( ~n1709 & n1710 ) ;
  assign n1712 = ( x502 & x503 ) | ( x502 & x504 ) | ( x503 & x504 ) ;
  assign n1713 = ( ~x502 & x503 ) | ( ~x502 & x504 ) | ( x503 & x504 ) ;
  assign n1714 = ( x502 & ~n1712 ) | ( x502 & n1713 ) | ( ~n1712 & n1713 ) ;
  assign n1715 = ( x499 & x500 ) | ( x499 & x501 ) | ( x500 & x501 ) ;
  assign n1716 = ( ~x499 & x500 ) | ( ~x499 & x501 ) | ( x500 & x501 ) ;
  assign n1717 = ( x499 & ~n1715 ) | ( x499 & n1716 ) | ( ~n1715 & n1716 ) ;
  assign n1718 = n1714 & n1717 ;
  assign n1719 = n1714 | n1717 ;
  assign n1720 = ~n1718 & n1719 ;
  assign n1721 = ( x505 & x506 ) | ( x505 & x507 ) | ( x506 & x507 ) ;
  assign n1722 = ( ~x505 & x506 ) | ( ~x505 & x507 ) | ( x506 & x507 ) ;
  assign n1723 = ( x505 & ~n1721 ) | ( x505 & n1722 ) | ( ~n1721 & n1722 ) ;
  assign n1724 = ( x508 & x509 ) | ( x508 & x510 ) | ( x509 & x510 ) ;
  assign n1725 = ( ~x508 & x509 ) | ( ~x508 & x510 ) | ( x509 & x510 ) ;
  assign n1726 = ( x508 & ~n1724 ) | ( x508 & n1725 ) | ( ~n1724 & n1725 ) ;
  assign n1727 = ( n1720 & n1723 ) | ( n1720 & n1726 ) | ( n1723 & n1726 ) ;
  assign n1728 = ( ~n1720 & n1723 ) | ( ~n1720 & n1726 ) | ( n1723 & n1726 ) ;
  assign n1729 = ( n1720 & ~n1727 ) | ( n1720 & n1728 ) | ( ~n1727 & n1728 ) ;
  assign n1730 = ( x490 & x491 ) | ( x490 & x492 ) | ( x491 & x492 ) ;
  assign n1731 = ( ~x490 & x491 ) | ( ~x490 & x492 ) | ( x491 & x492 ) ;
  assign n1732 = ( x490 & ~n1730 ) | ( x490 & n1731 ) | ( ~n1730 & n1731 ) ;
  assign n1733 = ( x487 & x488 ) | ( x487 & x489 ) | ( x488 & x489 ) ;
  assign n1734 = ( ~x487 & x488 ) | ( ~x487 & x489 ) | ( x488 & x489 ) ;
  assign n1735 = ( x487 & ~n1733 ) | ( x487 & n1734 ) | ( ~n1733 & n1734 ) ;
  assign n1736 = n1732 & n1735 ;
  assign n1737 = n1732 | n1735 ;
  assign n1738 = ~n1736 & n1737 ;
  assign n1739 = ( x493 & x494 ) | ( x493 & x495 ) | ( x494 & x495 ) ;
  assign n1740 = ( ~x493 & x494 ) | ( ~x493 & x495 ) | ( x494 & x495 ) ;
  assign n1741 = ( x493 & ~n1739 ) | ( x493 & n1740 ) | ( ~n1739 & n1740 ) ;
  assign n1742 = ( x496 & x497 ) | ( x496 & x498 ) | ( x497 & x498 ) ;
  assign n1743 = ( ~x496 & x497 ) | ( ~x496 & x498 ) | ( x497 & x498 ) ;
  assign n1744 = ( x496 & ~n1742 ) | ( x496 & n1743 ) | ( ~n1742 & n1743 ) ;
  assign n1745 = ( n1738 & n1741 ) | ( n1738 & n1744 ) | ( n1741 & n1744 ) ;
  assign n1746 = ( ~n1738 & n1741 ) | ( ~n1738 & n1744 ) | ( n1741 & n1744 ) ;
  assign n1747 = ( n1738 & ~n1745 ) | ( n1738 & n1746 ) | ( ~n1745 & n1746 ) ;
  assign n1748 = n1729 & n1747 ;
  assign n1749 = n1729 | n1747 ;
  assign n1750 = ~n1748 & n1749 ;
  assign n1751 = ( x466 & x467 ) | ( x466 & x468 ) | ( x467 & x468 ) ;
  assign n1752 = ( ~x466 & x467 ) | ( ~x466 & x468 ) | ( x467 & x468 ) ;
  assign n1753 = ( x466 & ~n1751 ) | ( x466 & n1752 ) | ( ~n1751 & n1752 ) ;
  assign n1754 = ( x463 & x464 ) | ( x463 & x465 ) | ( x464 & x465 ) ;
  assign n1755 = ( ~x463 & x464 ) | ( ~x463 & x465 ) | ( x464 & x465 ) ;
  assign n1756 = ( x463 & ~n1754 ) | ( x463 & n1755 ) | ( ~n1754 & n1755 ) ;
  assign n1757 = n1753 & n1756 ;
  assign n1758 = n1753 | n1756 ;
  assign n1759 = ~n1757 & n1758 ;
  assign n1760 = ( x469 & x470 ) | ( x469 & x471 ) | ( x470 & x471 ) ;
  assign n1761 = ( ~x469 & x470 ) | ( ~x469 & x471 ) | ( x470 & x471 ) ;
  assign n1762 = ( x469 & ~n1760 ) | ( x469 & n1761 ) | ( ~n1760 & n1761 ) ;
  assign n1763 = ( x472 & x473 ) | ( x472 & x474 ) | ( x473 & x474 ) ;
  assign n1764 = ( ~x472 & x473 ) | ( ~x472 & x474 ) | ( x473 & x474 ) ;
  assign n1765 = ( x472 & ~n1763 ) | ( x472 & n1764 ) | ( ~n1763 & n1764 ) ;
  assign n1766 = ( n1759 & n1762 ) | ( n1759 & n1765 ) | ( n1762 & n1765 ) ;
  assign n1767 = ( ~n1759 & n1762 ) | ( ~n1759 & n1765 ) | ( n1762 & n1765 ) ;
  assign n1768 = ( n1759 & ~n1766 ) | ( n1759 & n1767 ) | ( ~n1766 & n1767 ) ;
  assign n1769 = ( x475 & x476 ) | ( x475 & x477 ) | ( x476 & x477 ) ;
  assign n1770 = ( ~x475 & x476 ) | ( ~x475 & x477 ) | ( x476 & x477 ) ;
  assign n1771 = ( x475 & ~n1769 ) | ( x475 & n1770 ) | ( ~n1769 & n1770 ) ;
  assign n1772 = ( x478 & x479 ) | ( x478 & x480 ) | ( x479 & x480 ) ;
  assign n1773 = ( ~x478 & x479 ) | ( ~x478 & x480 ) | ( x479 & x480 ) ;
  assign n1774 = ( x478 & ~n1772 ) | ( x478 & n1773 ) | ( ~n1772 & n1773 ) ;
  assign n1775 = n1771 & n1774 ;
  assign n1776 = n1771 | n1774 ;
  assign n1777 = ~n1775 & n1776 ;
  assign n1778 = ( x484 & x485 ) | ( x484 & x486 ) | ( x485 & x486 ) ;
  assign n1779 = ( ~x484 & x485 ) | ( ~x484 & x486 ) | ( x485 & x486 ) ;
  assign n1780 = ( x484 & ~n1778 ) | ( x484 & n1779 ) | ( ~n1778 & n1779 ) ;
  assign n1781 = ( x481 & x482 ) | ( x481 & x483 ) | ( x482 & x483 ) ;
  assign n1782 = ( ~x481 & x482 ) | ( ~x481 & x483 ) | ( x482 & x483 ) ;
  assign n1783 = ( x481 & ~n1781 ) | ( x481 & n1782 ) | ( ~n1781 & n1782 ) ;
  assign n1784 = ( n1777 & n1780 ) | ( n1777 & n1783 ) | ( n1780 & n1783 ) ;
  assign n1785 = ( ~n1777 & n1780 ) | ( ~n1777 & n1783 ) | ( n1780 & n1783 ) ;
  assign n1786 = ( n1777 & ~n1784 ) | ( n1777 & n1785 ) | ( ~n1784 & n1785 ) ;
  assign n1787 = n1768 & n1786 ;
  assign n1788 = n1768 | n1786 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = n1750 & n1789 ;
  assign n1791 = n1750 | n1789 ;
  assign n1792 = ~n1790 & n1791 ;
  assign n1793 = ( x547 & x548 ) | ( x547 & x549 ) | ( x548 & x549 ) ;
  assign n1794 = ( ~x547 & x548 ) | ( ~x547 & x549 ) | ( x548 & x549 ) ;
  assign n1795 = ( x547 & ~n1793 ) | ( x547 & n1794 ) | ( ~n1793 & n1794 ) ;
  assign n1796 = x551 & x552 ;
  assign n1797 = x551 | x552 ;
  assign n1798 = ~n1796 & n1797 ;
  assign n1799 = ( x550 & n1795 ) | ( x550 & n1798 ) | ( n1795 & n1798 ) ;
  assign n1800 = ( ~x550 & n1795 ) | ( ~x550 & n1798 ) | ( n1795 & n1798 ) ;
  assign n1801 = ( x550 & ~n1799 ) | ( x550 & n1800 ) | ( ~n1799 & n1800 ) ;
  assign n1802 = ( x553 & x554 ) | ( x553 & x555 ) | ( x554 & x555 ) ;
  assign n1803 = ( ~x553 & x554 ) | ( ~x553 & x555 ) | ( x554 & x555 ) ;
  assign n1804 = ( x553 & ~n1802 ) | ( x553 & n1803 ) | ( ~n1802 & n1803 ) ;
  assign n1805 = ( x556 & x557 ) | ( x556 & x558 ) | ( x557 & x558 ) ;
  assign n1806 = ( ~x556 & x557 ) | ( ~x556 & x558 ) | ( x557 & x558 ) ;
  assign n1807 = ( x556 & ~n1805 ) | ( x556 & n1806 ) | ( ~n1805 & n1806 ) ;
  assign n1808 = ( n1801 & n1804 ) | ( n1801 & n1807 ) | ( n1804 & n1807 ) ;
  assign n1809 = ( ~n1801 & n1804 ) | ( ~n1801 & n1807 ) | ( n1804 & n1807 ) ;
  assign n1810 = ( n1801 & ~n1808 ) | ( n1801 & n1809 ) | ( ~n1808 & n1809 ) ;
  assign n1811 = ( x535 & x536 ) | ( x535 & x537 ) | ( x536 & x537 ) ;
  assign n1812 = ( ~x535 & x536 ) | ( ~x535 & x537 ) | ( x536 & x537 ) ;
  assign n1813 = ( x535 & ~n1811 ) | ( x535 & n1812 ) | ( ~n1811 & n1812 ) ;
  assign n1814 = ( x538 & x539 ) | ( x538 & x540 ) | ( x539 & x540 ) ;
  assign n1815 = ( ~x538 & x539 ) | ( ~x538 & x540 ) | ( x539 & x540 ) ;
  assign n1816 = ( x538 & ~n1814 ) | ( x538 & n1815 ) | ( ~n1814 & n1815 ) ;
  assign n1817 = n1813 & n1816 ;
  assign n1818 = n1813 | n1816 ;
  assign n1819 = ~n1817 & n1818 ;
  assign n1820 = ( x541 & x542 ) | ( x541 & x543 ) | ( x542 & x543 ) ;
  assign n1821 = ( ~x541 & x542 ) | ( ~x541 & x543 ) | ( x542 & x543 ) ;
  assign n1822 = ( x541 & ~n1820 ) | ( x541 & n1821 ) | ( ~n1820 & n1821 ) ;
  assign n1823 = ( x544 & x545 ) | ( x544 & x546 ) | ( x545 & x546 ) ;
  assign n1824 = ( ~x544 & x545 ) | ( ~x544 & x546 ) | ( x545 & x546 ) ;
  assign n1825 = ( x544 & ~n1823 ) | ( x544 & n1824 ) | ( ~n1823 & n1824 ) ;
  assign n1826 = ( n1819 & n1822 ) | ( n1819 & n1825 ) | ( n1822 & n1825 ) ;
  assign n1827 = ( ~n1819 & n1822 ) | ( ~n1819 & n1825 ) | ( n1822 & n1825 ) ;
  assign n1828 = ( n1819 & ~n1826 ) | ( n1819 & n1827 ) | ( ~n1826 & n1827 ) ;
  assign n1829 = n1810 & n1828 ;
  assign n1830 = n1810 | n1828 ;
  assign n1831 = ~n1829 & n1830 ;
  assign n1832 = ( ~x529 & x530 ) | ( ~x529 & x531 ) | ( x530 & x531 ) ;
  assign n1833 = ( x529 & x530 ) | ( x529 & x531 ) | ( x530 & x531 ) ;
  assign n1834 = ( x529 & n1832 ) | ( x529 & ~n1833 ) | ( n1832 & ~n1833 ) ;
  assign n1835 = ( ~x532 & x533 ) | ( ~x532 & x534 ) | ( x533 & x534 ) ;
  assign n1836 = ( x532 & x533 ) | ( x532 & x534 ) | ( x533 & x534 ) ;
  assign n1837 = ( x532 & n1835 ) | ( x532 & ~n1836 ) | ( n1835 & ~n1836 ) ;
  assign n1838 = ( x526 & x527 ) | ( x526 & x528 ) | ( x527 & x528 ) ;
  assign n1839 = ( ~x526 & x527 ) | ( ~x526 & x528 ) | ( x527 & x528 ) ;
  assign n1840 = ( x526 & ~n1838 ) | ( x526 & n1839 ) | ( ~n1838 & n1839 ) ;
  assign n1841 = ( x523 & x524 ) | ( x523 & x525 ) | ( x524 & x525 ) ;
  assign n1842 = ( ~x523 & x524 ) | ( ~x523 & x525 ) | ( x524 & x525 ) ;
  assign n1843 = ( x523 & ~n1841 ) | ( x523 & n1842 ) | ( ~n1841 & n1842 ) ;
  assign n1844 = n1840 & n1843 ;
  assign n1845 = n1840 | n1843 ;
  assign n1846 = ~n1844 & n1845 ;
  assign n1847 = ( n1834 & n1837 ) | ( n1834 & n1846 ) | ( n1837 & n1846 ) ;
  assign n1848 = ( ~n1834 & n1837 ) | ( ~n1834 & n1846 ) | ( n1837 & n1846 ) ;
  assign n1849 = ( n1834 & ~n1847 ) | ( n1834 & n1848 ) | ( ~n1847 & n1848 ) ;
  assign n1850 = ( x517 & x518 ) | ( x517 & x519 ) | ( x518 & x519 ) ;
  assign n1851 = ( ~x517 & x518 ) | ( ~x517 & x519 ) | ( x518 & x519 ) ;
  assign n1852 = ( x517 & ~n1850 ) | ( x517 & n1851 ) | ( ~n1850 & n1851 ) ;
  assign n1853 = ( x520 & x521 ) | ( x520 & x522 ) | ( x521 & x522 ) ;
  assign n1854 = ( ~x520 & x521 ) | ( ~x520 & x522 ) | ( x521 & x522 ) ;
  assign n1855 = ( x520 & ~n1853 ) | ( x520 & n1854 ) | ( ~n1853 & n1854 ) ;
  assign n1856 = ( x514 & x515 ) | ( x514 & x516 ) | ( x515 & x516 ) ;
  assign n1857 = ( ~x514 & x515 ) | ( ~x514 & x516 ) | ( x515 & x516 ) ;
  assign n1858 = ( x514 & ~n1856 ) | ( x514 & n1857 ) | ( ~n1856 & n1857 ) ;
  assign n1859 = ( x511 & x512 ) | ( x511 & x513 ) | ( x512 & x513 ) ;
  assign n1860 = ( ~x511 & x512 ) | ( ~x511 & x513 ) | ( x512 & x513 ) ;
  assign n1861 = ( x511 & ~n1859 ) | ( x511 & n1860 ) | ( ~n1859 & n1860 ) ;
  assign n1862 = n1858 & n1861 ;
  assign n1863 = n1858 | n1861 ;
  assign n1864 = ~n1862 & n1863 ;
  assign n1865 = ( n1852 & n1855 ) | ( n1852 & n1864 ) | ( n1855 & n1864 ) ;
  assign n1866 = ( ~n1852 & n1855 ) | ( ~n1852 & n1864 ) | ( n1855 & n1864 ) ;
  assign n1867 = ( n1852 & ~n1865 ) | ( n1852 & n1866 ) | ( ~n1865 & n1866 ) ;
  assign n1868 = n1849 & n1867 ;
  assign n1869 = n1849 | n1867 ;
  assign n1870 = ~n1868 & n1869 ;
  assign n1871 = n1831 & n1870 ;
  assign n1872 = n1831 | n1870 ;
  assign n1873 = ~n1871 & n1872 ;
  assign n1874 = n1792 & n1873 ;
  assign n1875 = n1792 | n1873 ;
  assign n1876 = ~n1874 & n1875 ;
  assign n1877 = ( x631 & x632 ) | ( x631 & x633 ) | ( x632 & x633 ) ;
  assign n1878 = ( ~x631 & x632 ) | ( ~x631 & x633 ) | ( x632 & x633 ) ;
  assign n1879 = ( x631 & ~n1877 ) | ( x631 & n1878 ) | ( ~n1877 & n1878 ) ;
  assign n1880 = ( x634 & x635 ) | ( x634 & x636 ) | ( x635 & x636 ) ;
  assign n1881 = ( ~x634 & x635 ) | ( ~x634 & x636 ) | ( x635 & x636 ) ;
  assign n1882 = ( x634 & ~n1880 ) | ( x634 & n1881 ) | ( ~n1880 & n1881 ) ;
  assign n1883 = n1879 & n1882 ;
  assign n1884 = n1879 | n1882 ;
  assign n1885 = ~n1883 & n1884 ;
  assign n1886 = ( x640 & x641 ) | ( x640 & x642 ) | ( x641 & x642 ) ;
  assign n1887 = ( ~x640 & x641 ) | ( ~x640 & x642 ) | ( x641 & x642 ) ;
  assign n1888 = ( x640 & ~n1886 ) | ( x640 & n1887 ) | ( ~n1886 & n1887 ) ;
  assign n1889 = ( x637 & x638 ) | ( x637 & x639 ) | ( x638 & x639 ) ;
  assign n1890 = ( ~x637 & x638 ) | ( ~x637 & x639 ) | ( x638 & x639 ) ;
  assign n1891 = ( x637 & ~n1889 ) | ( x637 & n1890 ) | ( ~n1889 & n1890 ) ;
  assign n1892 = ( n1885 & n1888 ) | ( n1885 & n1891 ) | ( n1888 & n1891 ) ;
  assign n1893 = ( ~n1885 & n1888 ) | ( ~n1885 & n1891 ) | ( n1888 & n1891 ) ;
  assign n1894 = ( n1885 & ~n1892 ) | ( n1885 & n1893 ) | ( ~n1892 & n1893 ) ;
  assign n1895 = ( x643 & x644 ) | ( x643 & x645 ) | ( x644 & x645 ) ;
  assign n1896 = ( ~x643 & x644 ) | ( ~x643 & x645 ) | ( x644 & x645 ) ;
  assign n1897 = ( x643 & ~n1895 ) | ( x643 & n1896 ) | ( ~n1895 & n1896 ) ;
  assign n1898 = ( x646 & x647 ) | ( x646 & x648 ) | ( x647 & x648 ) ;
  assign n1899 = ( ~x646 & x647 ) | ( ~x646 & x648 ) | ( x647 & x648 ) ;
  assign n1900 = ( x646 & ~n1898 ) | ( x646 & n1899 ) | ( ~n1898 & n1899 ) ;
  assign n1901 = n1897 & n1900 ;
  assign n1902 = n1897 | n1900 ;
  assign n1903 = ~n1901 & n1902 ;
  assign n1904 = ( x649 & x650 ) | ( x649 & x651 ) | ( x650 & x651 ) ;
  assign n1905 = ( ~x649 & x650 ) | ( ~x649 & x651 ) | ( x650 & x651 ) ;
  assign n1906 = ( x649 & ~n1904 ) | ( x649 & n1905 ) | ( ~n1904 & n1905 ) ;
  assign n1907 = ( x652 & x653 ) | ( x652 & x654 ) | ( x653 & x654 ) ;
  assign n1908 = ( ~x652 & x653 ) | ( ~x652 & x654 ) | ( x653 & x654 ) ;
  assign n1909 = ( x652 & ~n1907 ) | ( x652 & n1908 ) | ( ~n1907 & n1908 ) ;
  assign n1910 = ( n1903 & n1906 ) | ( n1903 & n1909 ) | ( n1906 & n1909 ) ;
  assign n1911 = ( ~n1903 & n1906 ) | ( ~n1903 & n1909 ) | ( n1906 & n1909 ) ;
  assign n1912 = ( n1903 & ~n1910 ) | ( n1903 & n1911 ) | ( ~n1910 & n1911 ) ;
  assign n1913 = n1894 & n1912 ;
  assign n1914 = n1894 | n1912 ;
  assign n1915 = ~n1913 & n1914 ;
  assign n1916 = ( x619 & x620 ) | ( x619 & x621 ) | ( x620 & x621 ) ;
  assign n1917 = ( ~x619 & x620 ) | ( ~x619 & x621 ) | ( x620 & x621 ) ;
  assign n1918 = ( x619 & ~n1916 ) | ( x619 & n1917 ) | ( ~n1916 & n1917 ) ;
  assign n1919 = ( x622 & x623 ) | ( x622 & x624 ) | ( x623 & x624 ) ;
  assign n1920 = ( ~x622 & x623 ) | ( ~x622 & x624 ) | ( x623 & x624 ) ;
  assign n1921 = ( x622 & ~n1919 ) | ( x622 & n1920 ) | ( ~n1919 & n1920 ) ;
  assign n1922 = n1918 & n1921 ;
  assign n1923 = n1918 | n1921 ;
  assign n1924 = ~n1922 & n1923 ;
  assign n1925 = ( x625 & x626 ) | ( x625 & x627 ) | ( x626 & x627 ) ;
  assign n1926 = ( ~x625 & x626 ) | ( ~x625 & x627 ) | ( x626 & x627 ) ;
  assign n1927 = ( x625 & ~n1925 ) | ( x625 & n1926 ) | ( ~n1925 & n1926 ) ;
  assign n1928 = ( x628 & x629 ) | ( x628 & x630 ) | ( x629 & x630 ) ;
  assign n1929 = ( ~x628 & x629 ) | ( ~x628 & x630 ) | ( x629 & x630 ) ;
  assign n1930 = ( x628 & ~n1928 ) | ( x628 & n1929 ) | ( ~n1928 & n1929 ) ;
  assign n1931 = ( n1924 & n1927 ) | ( n1924 & n1930 ) | ( n1927 & n1930 ) ;
  assign n1932 = ( ~n1924 & n1927 ) | ( ~n1924 & n1930 ) | ( n1927 & n1930 ) ;
  assign n1933 = ( n1924 & ~n1931 ) | ( n1924 & n1932 ) | ( ~n1931 & n1932 ) ;
  assign n1934 = ( x607 & x608 ) | ( x607 & x609 ) | ( x608 & x609 ) ;
  assign n1935 = ( ~x607 & x608 ) | ( ~x607 & x609 ) | ( x608 & x609 ) ;
  assign n1936 = ( x607 & ~n1934 ) | ( x607 & n1935 ) | ( ~n1934 & n1935 ) ;
  assign n1937 = ( x610 & x611 ) | ( x610 & x612 ) | ( x611 & x612 ) ;
  assign n1938 = ( ~x610 & x611 ) | ( ~x610 & x612 ) | ( x611 & x612 ) ;
  assign n1939 = ( x610 & ~n1937 ) | ( x610 & n1938 ) | ( ~n1937 & n1938 ) ;
  assign n1940 = n1936 & n1939 ;
  assign n1941 = n1936 | n1939 ;
  assign n1942 = ~n1940 & n1941 ;
  assign n1943 = ( ~x613 & x614 ) | ( ~x613 & x615 ) | ( x614 & x615 ) ;
  assign n1944 = ( x613 & x614 ) | ( x613 & x615 ) | ( x614 & x615 ) ;
  assign n1945 = ( x613 & n1943 ) | ( x613 & ~n1944 ) | ( n1943 & ~n1944 ) ;
  assign n1946 = ( ~x616 & x617 ) | ( ~x616 & x618 ) | ( x617 & x618 ) ;
  assign n1947 = ( x616 & x617 ) | ( x616 & x618 ) | ( x617 & x618 ) ;
  assign n1948 = ( x616 & n1946 ) | ( x616 & ~n1947 ) | ( n1946 & ~n1947 ) ;
  assign n1949 = ( n1942 & n1945 ) | ( n1942 & n1948 ) | ( n1945 & n1948 ) ;
  assign n1950 = ( ~n1942 & n1945 ) | ( ~n1942 & n1948 ) | ( n1945 & n1948 ) ;
  assign n1951 = ( n1942 & ~n1949 ) | ( n1942 & n1950 ) | ( ~n1949 & n1950 ) ;
  assign n1952 = n1933 & n1951 ;
  assign n1953 = n1933 | n1951 ;
  assign n1954 = ~n1952 & n1953 ;
  assign n1955 = n1915 & n1954 ;
  assign n1956 = n1915 | n1954 ;
  assign n1957 = ~n1955 & n1956 ;
  assign n1958 = ( x562 & x563 ) | ( x562 & x564 ) | ( x563 & x564 ) ;
  assign n1959 = ( ~x562 & x563 ) | ( ~x562 & x564 ) | ( x563 & x564 ) ;
  assign n1960 = ( x562 & ~n1958 ) | ( x562 & n1959 ) | ( ~n1958 & n1959 ) ;
  assign n1961 = ( x559 & x560 ) | ( x559 & x561 ) | ( x560 & x561 ) ;
  assign n1962 = ( ~x559 & x560 ) | ( ~x559 & x561 ) | ( x560 & x561 ) ;
  assign n1963 = ( x559 & ~n1961 ) | ( x559 & n1962 ) | ( ~n1961 & n1962 ) ;
  assign n1964 = n1960 & n1963 ;
  assign n1965 = n1960 | n1963 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1967 = ( x565 & x566 ) | ( x565 & x567 ) | ( x566 & x567 ) ;
  assign n1968 = ( ~x565 & x566 ) | ( ~x565 & x567 ) | ( x566 & x567 ) ;
  assign n1969 = ( x565 & ~n1967 ) | ( x565 & n1968 ) | ( ~n1967 & n1968 ) ;
  assign n1970 = ( x568 & x569 ) | ( x568 & x570 ) | ( x569 & x570 ) ;
  assign n1971 = ( ~x568 & x569 ) | ( ~x568 & x570 ) | ( x569 & x570 ) ;
  assign n1972 = ( x568 & ~n1970 ) | ( x568 & n1971 ) | ( ~n1970 & n1971 ) ;
  assign n1973 = ( n1966 & n1969 ) | ( n1966 & n1972 ) | ( n1969 & n1972 ) ;
  assign n1974 = ( ~n1966 & n1969 ) | ( ~n1966 & n1972 ) | ( n1969 & n1972 ) ;
  assign n1975 = ( n1966 & ~n1973 ) | ( n1966 & n1974 ) | ( ~n1973 & n1974 ) ;
  assign n1976 = ( x574 & x575 ) | ( x574 & x576 ) | ( x575 & x576 ) ;
  assign n1977 = ( ~x574 & x575 ) | ( ~x574 & x576 ) | ( x575 & x576 ) ;
  assign n1978 = ( x574 & ~n1976 ) | ( x574 & n1977 ) | ( ~n1976 & n1977 ) ;
  assign n1979 = ( x571 & x572 ) | ( x571 & x573 ) | ( x572 & x573 ) ;
  assign n1980 = ( ~x571 & x572 ) | ( ~x571 & x573 ) | ( x572 & x573 ) ;
  assign n1981 = ( x571 & ~n1979 ) | ( x571 & n1980 ) | ( ~n1979 & n1980 ) ;
  assign n1982 = n1978 & n1981 ;
  assign n1983 = n1978 | n1981 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = ( x580 & x581 ) | ( x580 & x582 ) | ( x581 & x582 ) ;
  assign n1986 = ( ~x580 & x581 ) | ( ~x580 & x582 ) | ( x581 & x582 ) ;
  assign n1987 = ( x580 & ~n1985 ) | ( x580 & n1986 ) | ( ~n1985 & n1986 ) ;
  assign n1988 = ( x577 & x578 ) | ( x577 & x579 ) | ( x578 & x579 ) ;
  assign n1989 = ( ~x577 & x578 ) | ( ~x577 & x579 ) | ( x578 & x579 ) ;
  assign n1990 = ( x577 & ~n1988 ) | ( x577 & n1989 ) | ( ~n1988 & n1989 ) ;
  assign n1991 = ( n1984 & n1987 ) | ( n1984 & n1990 ) | ( n1987 & n1990 ) ;
  assign n1992 = ( ~n1984 & n1987 ) | ( ~n1984 & n1990 ) | ( n1987 & n1990 ) ;
  assign n1993 = ( n1984 & ~n1991 ) | ( n1984 & n1992 ) | ( ~n1991 & n1992 ) ;
  assign n1994 = n1975 & n1993 ;
  assign n1995 = n1975 | n1993 ;
  assign n1996 = ~n1994 & n1995 ;
  assign n1997 = ( x595 & x596 ) | ( x595 & x597 ) | ( x596 & x597 ) ;
  assign n1998 = ( ~x595 & x596 ) | ( ~x595 & x597 ) | ( x596 & x597 ) ;
  assign n1999 = ( x595 & ~n1997 ) | ( x595 & n1998 ) | ( ~n1997 & n1998 ) ;
  assign n2000 = ( x598 & x599 ) | ( x598 & x600 ) | ( x599 & x600 ) ;
  assign n2001 = ( ~x598 & x599 ) | ( ~x598 & x600 ) | ( x599 & x600 ) ;
  assign n2002 = ( x598 & ~n2000 ) | ( x598 & n2001 ) | ( ~n2000 & n2001 ) ;
  assign n2003 = n1999 & n2002 ;
  assign n2004 = n1999 | n2002 ;
  assign n2005 = ~n2003 & n2004 ;
  assign n2006 = ( x601 & x602 ) | ( x601 & x603 ) | ( x602 & x603 ) ;
  assign n2007 = ( ~x601 & x602 ) | ( ~x601 & x603 ) | ( x602 & x603 ) ;
  assign n2008 = ( x601 & ~n2006 ) | ( x601 & n2007 ) | ( ~n2006 & n2007 ) ;
  assign n2009 = ( x604 & x605 ) | ( x604 & x606 ) | ( x605 & x606 ) ;
  assign n2010 = ( ~x604 & x605 ) | ( ~x604 & x606 ) | ( x605 & x606 ) ;
  assign n2011 = ( x604 & ~n2009 ) | ( x604 & n2010 ) | ( ~n2009 & n2010 ) ;
  assign n2012 = ( n2005 & n2008 ) | ( n2005 & n2011 ) | ( n2008 & n2011 ) ;
  assign n2013 = ( ~n2005 & n2008 ) | ( ~n2005 & n2011 ) | ( n2008 & n2011 ) ;
  assign n2014 = ( n2005 & ~n2012 ) | ( n2005 & n2013 ) | ( ~n2012 & n2013 ) ;
  assign n2015 = ( x583 & x584 ) | ( x583 & x585 ) | ( x584 & x585 ) ;
  assign n2016 = ( ~x583 & x584 ) | ( ~x583 & x585 ) | ( x584 & x585 ) ;
  assign n2017 = ( x583 & ~n2015 ) | ( x583 & n2016 ) | ( ~n2015 & n2016 ) ;
  assign n2018 = ( x586 & x587 ) | ( x586 & x588 ) | ( x587 & x588 ) ;
  assign n2019 = ( ~x586 & x587 ) | ( ~x586 & x588 ) | ( x587 & x588 ) ;
  assign n2020 = ( x586 & ~n2018 ) | ( x586 & n2019 ) | ( ~n2018 & n2019 ) ;
  assign n2021 = n2017 & n2020 ;
  assign n2022 = n2017 | n2020 ;
  assign n2023 = ~n2021 & n2022 ;
  assign n2024 = ( x589 & x590 ) | ( x589 & x591 ) | ( x590 & x591 ) ;
  assign n2025 = ( ~x589 & x590 ) | ( ~x589 & x591 ) | ( x590 & x591 ) ;
  assign n2026 = ( x589 & ~n2024 ) | ( x589 & n2025 ) | ( ~n2024 & n2025 ) ;
  assign n2027 = ( x592 & x593 ) | ( x592 & x594 ) | ( x593 & x594 ) ;
  assign n2028 = ( ~x592 & x593 ) | ( ~x592 & x594 ) | ( x593 & x594 ) ;
  assign n2029 = ( x592 & ~n2027 ) | ( x592 & n2028 ) | ( ~n2027 & n2028 ) ;
  assign n2030 = ( n2023 & n2026 ) | ( n2023 & n2029 ) | ( n2026 & n2029 ) ;
  assign n2031 = ( ~n2023 & n2026 ) | ( ~n2023 & n2029 ) | ( n2026 & n2029 ) ;
  assign n2032 = ( n2023 & ~n2030 ) | ( n2023 & n2031 ) | ( ~n2030 & n2031 ) ;
  assign n2033 = n2014 & n2032 ;
  assign n2034 = n2014 | n2032 ;
  assign n2035 = ~n2033 & n2034 ;
  assign n2036 = n1996 & n2035 ;
  assign n2037 = n1996 | n2035 ;
  assign n2038 = ~n2036 & n2037 ;
  assign n2039 = n1957 & n2038 ;
  assign n2040 = n1957 | n2038 ;
  assign n2041 = ~n2039 & n2040 ;
  assign n2042 = n1876 & n2041 ;
  assign n2043 = n1876 | n2041 ;
  assign n2044 = ~n2042 & n2043 ;
  assign n2045 = n1163 | n1328 ;
  assign n2046 = ~n1329 & n2045 ;
  assign n2047 = n2044 & n2046 ;
  assign n2048 = ( n1769 & n1772 ) | ( n1769 & n1775 ) | ( n1772 & n1775 ) ;
  assign n2049 = ( ~n1769 & n1772 ) | ( ~n1769 & n1775 ) | ( n1772 & n1775 ) ;
  assign n2050 = ( n1769 & ~n2048 ) | ( n1769 & n2049 ) | ( ~n2048 & n2049 ) ;
  assign n2051 = n1778 & n1781 ;
  assign n2052 = n1778 | n1781 ;
  assign n2053 = ~n2051 & n2052 ;
  assign n2054 = ( n1784 & n2050 ) | ( n1784 & n2053 ) | ( n2050 & n2053 ) ;
  assign n2055 = ( ~n1784 & n2050 ) | ( ~n1784 & n2053 ) | ( n2050 & n2053 ) ;
  assign n2056 = ( n1784 & ~n2054 ) | ( n1784 & n2055 ) | ( ~n2054 & n2055 ) ;
  assign n2057 = ( n1751 & n1754 ) | ( n1751 & n1757 ) | ( n1754 & n1757 ) ;
  assign n2058 = ( ~n1751 & n1754 ) | ( ~n1751 & n1757 ) | ( n1754 & n1757 ) ;
  assign n2059 = ( n1751 & ~n2057 ) | ( n1751 & n2058 ) | ( ~n2057 & n2058 ) ;
  assign n2060 = n1760 & n1763 ;
  assign n2061 = n1760 | n1763 ;
  assign n2062 = ~n2060 & n2061 ;
  assign n2063 = ( n1766 & n2059 ) | ( n1766 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2064 = ( ~n1766 & n2059 ) | ( ~n1766 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2065 = ( n1766 & ~n2063 ) | ( n1766 & n2064 ) | ( ~n2063 & n2064 ) ;
  assign n2066 = ( n1787 & n2056 ) | ( n1787 & n2065 ) | ( n2056 & n2065 ) ;
  assign n2067 = ( n1787 & ~n2056 ) | ( n1787 & n2065 ) | ( ~n2056 & n2065 ) ;
  assign n2068 = ( n2056 & ~n2066 ) | ( n2056 & n2067 ) | ( ~n2066 & n2067 ) ;
  assign n2069 = ( n1712 & n1715 ) | ( n1712 & n1718 ) | ( n1715 & n1718 ) ;
  assign n2070 = ( ~n1712 & n1715 ) | ( ~n1712 & n1718 ) | ( n1715 & n1718 ) ;
  assign n2071 = ( n1712 & ~n2069 ) | ( n1712 & n2070 ) | ( ~n2069 & n2070 ) ;
  assign n2072 = n1721 & n1724 ;
  assign n2073 = n1721 | n1724 ;
  assign n2074 = ~n2072 & n2073 ;
  assign n2075 = ( n1727 & n2071 ) | ( n1727 & n2074 ) | ( n2071 & n2074 ) ;
  assign n2076 = ( ~n1727 & n2071 ) | ( ~n1727 & n2074 ) | ( n2071 & n2074 ) ;
  assign n2077 = ( n1727 & ~n2075 ) | ( n1727 & n2076 ) | ( ~n2075 & n2076 ) ;
  assign n2078 = ( n1730 & n1733 ) | ( n1730 & n1736 ) | ( n1733 & n1736 ) ;
  assign n2079 = ( ~n1730 & n1733 ) | ( ~n1730 & n1736 ) | ( n1733 & n1736 ) ;
  assign n2080 = ( n1730 & ~n2078 ) | ( n1730 & n2079 ) | ( ~n2078 & n2079 ) ;
  assign n2081 = n1739 & n1742 ;
  assign n2082 = n1739 | n1742 ;
  assign n2083 = ~n2081 & n2082 ;
  assign n2084 = ( n1745 & n2080 ) | ( n1745 & n2083 ) | ( n2080 & n2083 ) ;
  assign n2085 = ( ~n1745 & n2080 ) | ( ~n1745 & n2083 ) | ( n2080 & n2083 ) ;
  assign n2086 = ( n1745 & ~n2084 ) | ( n1745 & n2085 ) | ( ~n2084 & n2085 ) ;
  assign n2087 = ( n1748 & n2077 ) | ( n1748 & n2086 ) | ( n2077 & n2086 ) ;
  assign n2088 = ( n1748 & ~n2077 ) | ( n1748 & n2086 ) | ( ~n2077 & n2086 ) ;
  assign n2089 = ( n2077 & ~n2087 ) | ( n2077 & n2088 ) | ( ~n2087 & n2088 ) ;
  assign n2090 = ( n1790 & n2068 ) | ( n1790 & n2089 ) | ( n2068 & n2089 ) ;
  assign n2091 = ( ~n1790 & n2068 ) | ( ~n1790 & n2089 ) | ( n2068 & n2089 ) ;
  assign n2092 = ( n1790 & ~n2090 ) | ( n1790 & n2091 ) | ( ~n2090 & n2091 ) ;
  assign n2093 = ( n1838 & n1841 ) | ( n1838 & n1844 ) | ( n1841 & n1844 ) ;
  assign n2094 = ( ~n1838 & n1841 ) | ( ~n1838 & n1844 ) | ( n1841 & n1844 ) ;
  assign n2095 = ( n1838 & ~n2093 ) | ( n1838 & n2094 ) | ( ~n2093 & n2094 ) ;
  assign n2096 = n1833 & n1836 ;
  assign n2097 = n1833 | n1836 ;
  assign n2098 = ~n2096 & n2097 ;
  assign n2099 = ( n1847 & n2095 ) | ( n1847 & n2098 ) | ( n2095 & n2098 ) ;
  assign n2100 = ( ~n1847 & n2095 ) | ( ~n1847 & n2098 ) | ( n2095 & n2098 ) ;
  assign n2101 = ( n1847 & ~n2099 ) | ( n1847 & n2100 ) | ( ~n2099 & n2100 ) ;
  assign n2102 = ( n1856 & n1859 ) | ( n1856 & n1862 ) | ( n1859 & n1862 ) ;
  assign n2103 = ( ~n1856 & n1859 ) | ( ~n1856 & n1862 ) | ( n1859 & n1862 ) ;
  assign n2104 = ( n1856 & ~n2102 ) | ( n1856 & n2103 ) | ( ~n2102 & n2103 ) ;
  assign n2105 = n1850 & n1853 ;
  assign n2106 = n1850 | n1853 ;
  assign n2107 = ~n2105 & n2106 ;
  assign n2108 = ( ~n1865 & n2104 ) | ( ~n1865 & n2107 ) | ( n2104 & n2107 ) ;
  assign n2109 = ( n1865 & n2104 ) | ( n1865 & n2107 ) | ( n2104 & n2107 ) ;
  assign n2110 = ( n1865 & n2108 ) | ( n1865 & ~n2109 ) | ( n2108 & ~n2109 ) ;
  assign n2111 = ( n1868 & n2101 ) | ( n1868 & n2110 ) | ( n2101 & n2110 ) ;
  assign n2112 = ( n1868 & ~n2101 ) | ( n1868 & n2110 ) | ( ~n2101 & n2110 ) ;
  assign n2113 = ( n2101 & ~n2111 ) | ( n2101 & n2112 ) | ( ~n2111 & n2112 ) ;
  assign n2114 = ( n1811 & n1814 ) | ( n1811 & n1817 ) | ( n1814 & n1817 ) ;
  assign n2115 = ( ~n1811 & n1814 ) | ( ~n1811 & n1817 ) | ( n1814 & n1817 ) ;
  assign n2116 = ( n1811 & ~n2114 ) | ( n1811 & n2115 ) | ( ~n2114 & n2115 ) ;
  assign n2117 = n1820 & n1823 ;
  assign n2118 = n1820 | n1823 ;
  assign n2119 = ~n2117 & n2118 ;
  assign n2120 = ( n1826 & n2116 ) | ( n1826 & n2119 ) | ( n2116 & n2119 ) ;
  assign n2121 = ( ~n1826 & n2116 ) | ( ~n1826 & n2119 ) | ( n2116 & n2119 ) ;
  assign n2122 = ( n1826 & ~n2120 ) | ( n1826 & n2121 ) | ( ~n2120 & n2121 ) ;
  assign n2123 = n1802 & n1805 ;
  assign n2124 = n1802 | n1805 ;
  assign n2125 = ~n2123 & n2124 ;
  assign n2126 = n1804 & n1807 ;
  assign n2127 = n2125 & ~n2126 ;
  assign n2128 = ( n1808 & ~n2125 ) | ( n1808 & n2127 ) | ( ~n2125 & n2127 ) ;
  assign n2129 = ( n1793 & n1796 ) | ( n1793 & n1799 ) | ( n1796 & n1799 ) ;
  assign n2130 = ( n1793 & n1796 ) | ( n1793 & ~n1799 ) | ( n1796 & ~n1799 ) ;
  assign n2131 = ( n1799 & ~n2129 ) | ( n1799 & n2130 ) | ( ~n2129 & n2130 ) ;
  assign n2132 = ( n2127 & n2128 ) | ( n2127 & n2131 ) | ( n2128 & n2131 ) ;
  assign n2133 = ( n2127 & ~n2128 ) | ( n2127 & n2131 ) | ( ~n2128 & n2131 ) ;
  assign n2134 = ( n2128 & ~n2132 ) | ( n2128 & n2133 ) | ( ~n2132 & n2133 ) ;
  assign n2135 = ( n1829 & n2122 ) | ( n1829 & n2134 ) | ( n2122 & n2134 ) ;
  assign n2136 = ( ~n1829 & n2122 ) | ( ~n1829 & n2134 ) | ( n2122 & n2134 ) ;
  assign n2137 = ( n1829 & ~n2135 ) | ( n1829 & n2136 ) | ( ~n2135 & n2136 ) ;
  assign n2138 = ( n1871 & n2113 ) | ( n1871 & n2137 ) | ( n2113 & n2137 ) ;
  assign n2139 = ( n1871 & ~n2113 ) | ( n1871 & n2137 ) | ( ~n2113 & n2137 ) ;
  assign n2140 = ( n2113 & ~n2138 ) | ( n2113 & n2139 ) | ( ~n2138 & n2139 ) ;
  assign n2141 = ( n1874 & n2092 ) | ( n1874 & n2140 ) | ( n2092 & n2140 ) ;
  assign n2142 = ( n1874 & ~n2092 ) | ( n1874 & n2140 ) | ( ~n2092 & n2140 ) ;
  assign n2143 = ( n2092 & ~n2141 ) | ( n2092 & n2142 ) | ( ~n2141 & n2142 ) ;
  assign n2144 = ( n2015 & n2018 ) | ( n2015 & n2021 ) | ( n2018 & n2021 ) ;
  assign n2145 = ( ~n2015 & n2018 ) | ( ~n2015 & n2021 ) | ( n2018 & n2021 ) ;
  assign n2146 = ( n2015 & ~n2144 ) | ( n2015 & n2145 ) | ( ~n2144 & n2145 ) ;
  assign n2147 = n2024 & n2027 ;
  assign n2148 = n2024 | n2027 ;
  assign n2149 = ~n2147 & n2148 ;
  assign n2150 = ( n2030 & n2146 ) | ( n2030 & n2149 ) | ( n2146 & n2149 ) ;
  assign n2151 = ( ~n2030 & n2146 ) | ( ~n2030 & n2149 ) | ( n2146 & n2149 ) ;
  assign n2152 = ( n2030 & ~n2150 ) | ( n2030 & n2151 ) | ( ~n2150 & n2151 ) ;
  assign n2153 = ( n1997 & n2000 ) | ( n1997 & n2003 ) | ( n2000 & n2003 ) ;
  assign n2154 = ( ~n1997 & n2000 ) | ( ~n1997 & n2003 ) | ( n2000 & n2003 ) ;
  assign n2155 = ( n1997 & ~n2153 ) | ( n1997 & n2154 ) | ( ~n2153 & n2154 ) ;
  assign n2156 = n2006 & n2009 ;
  assign n2157 = n2006 | n2009 ;
  assign n2158 = ~n2156 & n2157 ;
  assign n2159 = ( n2012 & n2155 ) | ( n2012 & n2158 ) | ( n2155 & n2158 ) ;
  assign n2160 = ( ~n2012 & n2155 ) | ( ~n2012 & n2158 ) | ( n2155 & n2158 ) ;
  assign n2161 = ( n2012 & ~n2159 ) | ( n2012 & n2160 ) | ( ~n2159 & n2160 ) ;
  assign n2162 = ( n2033 & n2152 ) | ( n2033 & n2161 ) | ( n2152 & n2161 ) ;
  assign n2163 = ( n2033 & ~n2152 ) | ( n2033 & n2161 ) | ( ~n2152 & n2161 ) ;
  assign n2164 = ( n2152 & ~n2162 ) | ( n2152 & n2163 ) | ( ~n2162 & n2163 ) ;
  assign n2165 = ( n1958 & n1961 ) | ( n1958 & n1964 ) | ( n1961 & n1964 ) ;
  assign n2166 = ( ~n1958 & n1961 ) | ( ~n1958 & n1964 ) | ( n1961 & n1964 ) ;
  assign n2167 = ( n1958 & ~n2165 ) | ( n1958 & n2166 ) | ( ~n2165 & n2166 ) ;
  assign n2168 = n1967 & n1970 ;
  assign n2169 = n1967 | n1970 ;
  assign n2170 = ~n2168 & n2169 ;
  assign n2171 = ( n1973 & n2167 ) | ( n1973 & n2170 ) | ( n2167 & n2170 ) ;
  assign n2172 = ( ~n1973 & n2167 ) | ( ~n1973 & n2170 ) | ( n2167 & n2170 ) ;
  assign n2173 = ( n1973 & ~n2171 ) | ( n1973 & n2172 ) | ( ~n2171 & n2172 ) ;
  assign n2174 = ( n1976 & n1979 ) | ( n1976 & n1982 ) | ( n1979 & n1982 ) ;
  assign n2175 = ( ~n1976 & n1979 ) | ( ~n1976 & n1982 ) | ( n1979 & n1982 ) ;
  assign n2176 = ( n1976 & ~n2174 ) | ( n1976 & n2175 ) | ( ~n2174 & n2175 ) ;
  assign n2177 = n1985 & n1988 ;
  assign n2178 = n1985 | n1988 ;
  assign n2179 = ~n2177 & n2178 ;
  assign n2180 = ( n1991 & n2176 ) | ( n1991 & n2179 ) | ( n2176 & n2179 ) ;
  assign n2181 = ( ~n1991 & n2176 ) | ( ~n1991 & n2179 ) | ( n2176 & n2179 ) ;
  assign n2182 = ( n1991 & ~n2180 ) | ( n1991 & n2181 ) | ( ~n2180 & n2181 ) ;
  assign n2183 = ( n1994 & n2173 ) | ( n1994 & n2182 ) | ( n2173 & n2182 ) ;
  assign n2184 = ( n1994 & ~n2173 ) | ( n1994 & n2182 ) | ( ~n2173 & n2182 ) ;
  assign n2185 = ( n2173 & ~n2183 ) | ( n2173 & n2184 ) | ( ~n2183 & n2184 ) ;
  assign n2186 = ( n2036 & n2164 ) | ( n2036 & n2185 ) | ( n2164 & n2185 ) ;
  assign n2187 = ( n2036 & ~n2164 ) | ( n2036 & n2185 ) | ( ~n2164 & n2185 ) ;
  assign n2188 = ( n2164 & ~n2186 ) | ( n2164 & n2187 ) | ( ~n2186 & n2187 ) ;
  assign n2189 = ( n1934 & n1937 ) | ( n1934 & n1940 ) | ( n1937 & n1940 ) ;
  assign n2190 = ( ~n1934 & n1937 ) | ( ~n1934 & n1940 ) | ( n1937 & n1940 ) ;
  assign n2191 = ( n1934 & ~n2189 ) | ( n1934 & n2190 ) | ( ~n2189 & n2190 ) ;
  assign n2192 = n1944 | n1947 ;
  assign n2193 = n1944 & n1947 ;
  assign n2194 = n2192 & ~n2193 ;
  assign n2195 = ( n1949 & n2191 ) | ( n1949 & n2194 ) | ( n2191 & n2194 ) ;
  assign n2196 = ( n1949 & ~n2191 ) | ( n1949 & n2194 ) | ( ~n2191 & n2194 ) ;
  assign n2197 = ( n2191 & ~n2195 ) | ( n2191 & n2196 ) | ( ~n2195 & n2196 ) ;
  assign n2198 = ( n1916 & n1919 ) | ( n1916 & n1922 ) | ( n1919 & n1922 ) ;
  assign n2199 = ( ~n1916 & n1919 ) | ( ~n1916 & n1922 ) | ( n1919 & n1922 ) ;
  assign n2200 = ( n1916 & ~n2198 ) | ( n1916 & n2199 ) | ( ~n2198 & n2199 ) ;
  assign n2201 = n1925 & n1928 ;
  assign n2202 = n1925 | n1928 ;
  assign n2203 = ~n2201 & n2202 ;
  assign n2204 = ( n1931 & n2200 ) | ( n1931 & n2203 ) | ( n2200 & n2203 ) ;
  assign n2205 = ( ~n1931 & n2200 ) | ( ~n1931 & n2203 ) | ( n2200 & n2203 ) ;
  assign n2206 = ( n1931 & ~n2204 ) | ( n1931 & n2205 ) | ( ~n2204 & n2205 ) ;
  assign n2207 = ( n1952 & n2197 ) | ( n1952 & n2206 ) | ( n2197 & n2206 ) ;
  assign n2208 = ( n1952 & ~n2197 ) | ( n1952 & n2206 ) | ( ~n2197 & n2206 ) ;
  assign n2209 = ( n2197 & ~n2207 ) | ( n2197 & n2208 ) | ( ~n2207 & n2208 ) ;
  assign n2210 = ( n1895 & n1898 ) | ( n1895 & n1901 ) | ( n1898 & n1901 ) ;
  assign n2211 = ( ~n1895 & n1898 ) | ( ~n1895 & n1901 ) | ( n1898 & n1901 ) ;
  assign n2212 = ( n1895 & ~n2210 ) | ( n1895 & n2211 ) | ( ~n2210 & n2211 ) ;
  assign n2213 = n1904 & n1907 ;
  assign n2214 = n1904 | n1907 ;
  assign n2215 = ~n2213 & n2214 ;
  assign n2216 = ( n1910 & n2212 ) | ( n1910 & n2215 ) | ( n2212 & n2215 ) ;
  assign n2217 = ( ~n1910 & n2212 ) | ( ~n1910 & n2215 ) | ( n2212 & n2215 ) ;
  assign n2218 = ( n1910 & ~n2216 ) | ( n1910 & n2217 ) | ( ~n2216 & n2217 ) ;
  assign n2219 = ( n1877 & n1880 ) | ( n1877 & n1883 ) | ( n1880 & n1883 ) ;
  assign n2220 = ( ~n1877 & n1880 ) | ( ~n1877 & n1883 ) | ( n1880 & n1883 ) ;
  assign n2221 = ( n1877 & ~n2219 ) | ( n1877 & n2220 ) | ( ~n2219 & n2220 ) ;
  assign n2222 = n1886 & n1889 ;
  assign n2223 = n1886 | n1889 ;
  assign n2224 = ~n2222 & n2223 ;
  assign n2225 = ( n1892 & n2221 ) | ( n1892 & n2224 ) | ( n2221 & n2224 ) ;
  assign n2226 = ( ~n1892 & n2221 ) | ( ~n1892 & n2224 ) | ( n2221 & n2224 ) ;
  assign n2227 = ( n1892 & ~n2225 ) | ( n1892 & n2226 ) | ( ~n2225 & n2226 ) ;
  assign n2228 = ( n1913 & n2218 ) | ( n1913 & n2227 ) | ( n2218 & n2227 ) ;
  assign n2229 = ( n1913 & ~n2218 ) | ( n1913 & n2227 ) | ( ~n2218 & n2227 ) ;
  assign n2230 = ( n2218 & ~n2228 ) | ( n2218 & n2229 ) | ( ~n2228 & n2229 ) ;
  assign n2231 = ( n1955 & n2209 ) | ( n1955 & n2230 ) | ( n2209 & n2230 ) ;
  assign n2232 = ( n1955 & ~n2209 ) | ( n1955 & n2230 ) | ( ~n2209 & n2230 ) ;
  assign n2233 = ( n2209 & ~n2231 ) | ( n2209 & n2232 ) | ( ~n2231 & n2232 ) ;
  assign n2234 = ( n2039 & n2188 ) | ( n2039 & n2233 ) | ( n2188 & n2233 ) ;
  assign n2235 = ( ~n2039 & n2188 ) | ( ~n2039 & n2233 ) | ( n2188 & n2233 ) ;
  assign n2236 = ( n2039 & ~n2234 ) | ( n2039 & n2235 ) | ( ~n2234 & n2235 ) ;
  assign n2237 = ( n2042 & n2143 ) | ( n2042 & n2236 ) | ( n2143 & n2236 ) ;
  assign n2238 = ( ~n2042 & n2143 ) | ( ~n2042 & n2236 ) | ( n2143 & n2236 ) ;
  assign n2239 = ( n2042 & ~n2237 ) | ( n2042 & n2238 ) | ( ~n2237 & n2238 ) ;
  assign n2240 = ( n1329 & ~n1428 ) | ( n1329 & n1521 ) | ( ~n1428 & n1521 ) ;
  assign n2241 = ( n1428 & ~n1522 ) | ( n1428 & n2240 ) | ( ~n1522 & n2240 ) ;
  assign n2242 = ( n2047 & n2239 ) | ( n2047 & n2241 ) | ( n2239 & n2241 ) ;
  assign n2243 = ( ~n1522 & n1577 ) | ( ~n1522 & n1638 ) | ( n1577 & n1638 ) ;
  assign n2244 = ( n1522 & ~n1639 ) | ( n1522 & n2243 ) | ( ~n1639 & n2243 ) ;
  assign n2245 = ( n2210 & n2213 ) | ( n2210 & n2216 ) | ( n2213 & n2216 ) ;
  assign n2246 = ( n2210 & n2213 ) | ( n2210 & ~n2216 ) | ( n2213 & ~n2216 ) ;
  assign n2247 = ( n2216 & ~n2245 ) | ( n2216 & n2246 ) | ( ~n2245 & n2246 ) ;
  assign n2248 = ( n2219 & n2222 ) | ( n2219 & n2225 ) | ( n2222 & n2225 ) ;
  assign n2249 = ( n2219 & n2222 ) | ( n2219 & ~n2225 ) | ( n2222 & ~n2225 ) ;
  assign n2250 = ( n2225 & ~n2248 ) | ( n2225 & n2249 ) | ( ~n2248 & n2249 ) ;
  assign n2251 = ( n2228 & n2247 ) | ( n2228 & n2250 ) | ( n2247 & n2250 ) ;
  assign n2252 = ( n2228 & ~n2247 ) | ( n2228 & n2250 ) | ( ~n2247 & n2250 ) ;
  assign n2253 = ( n2247 & ~n2251 ) | ( n2247 & n2252 ) | ( ~n2251 & n2252 ) ;
  assign n2254 = ( n2198 & n2201 ) | ( n2198 & n2204 ) | ( n2201 & n2204 ) ;
  assign n2255 = ( n2198 & n2201 ) | ( n2198 & ~n2204 ) | ( n2201 & ~n2204 ) ;
  assign n2256 = ( n2204 & ~n2254 ) | ( n2204 & n2255 ) | ( ~n2254 & n2255 ) ;
  assign n2257 = n1950 & ~n2196 ;
  assign n2258 = ( ~n1950 & n2195 ) | ( ~n1950 & n2257 ) | ( n2195 & n2257 ) ;
  assign n2259 = n1945 & n1948 ;
  assign n2260 = ( n1944 & n1947 ) | ( n1944 & n2259 ) | ( n1947 & n2259 ) ;
  assign n2261 = ( n2189 & n2258 ) | ( n2189 & n2260 ) | ( n2258 & n2260 ) ;
  assign n2262 = ( n2189 & ~n2258 ) | ( n2189 & n2260 ) | ( ~n2258 & n2260 ) ;
  assign n2263 = ( n2258 & ~n2261 ) | ( n2258 & n2262 ) | ( ~n2261 & n2262 ) ;
  assign n2264 = ( n2207 & n2256 ) | ( n2207 & n2263 ) | ( n2256 & n2263 ) ;
  assign n2265 = ( ~n2207 & n2256 ) | ( ~n2207 & n2263 ) | ( n2256 & n2263 ) ;
  assign n2266 = ( n2207 & ~n2264 ) | ( n2207 & n2265 ) | ( ~n2264 & n2265 ) ;
  assign n2267 = ( n2231 & n2253 ) | ( n2231 & n2266 ) | ( n2253 & n2266 ) ;
  assign n2268 = ( ~n2231 & n2253 ) | ( ~n2231 & n2266 ) | ( n2253 & n2266 ) ;
  assign n2269 = ( n2231 & ~n2267 ) | ( n2231 & n2268 ) | ( ~n2267 & n2268 ) ;
  assign n2270 = ( n2153 & n2156 ) | ( n2153 & n2159 ) | ( n2156 & n2159 ) ;
  assign n2271 = ( n2153 & n2156 ) | ( n2153 & ~n2159 ) | ( n2156 & ~n2159 ) ;
  assign n2272 = ( n2159 & ~n2270 ) | ( n2159 & n2271 ) | ( ~n2270 & n2271 ) ;
  assign n2273 = ( n2144 & n2147 ) | ( n2144 & n2150 ) | ( n2147 & n2150 ) ;
  assign n2274 = ( n2144 & n2147 ) | ( n2144 & ~n2150 ) | ( n2147 & ~n2150 ) ;
  assign n2275 = ( n2150 & ~n2273 ) | ( n2150 & n2274 ) | ( ~n2273 & n2274 ) ;
  assign n2276 = ( n2162 & n2272 ) | ( n2162 & n2275 ) | ( n2272 & n2275 ) ;
  assign n2277 = ( ~n2162 & n2272 ) | ( ~n2162 & n2275 ) | ( n2272 & n2275 ) ;
  assign n2278 = ( n2162 & ~n2276 ) | ( n2162 & n2277 ) | ( ~n2276 & n2277 ) ;
  assign n2279 = ( n2165 & n2168 ) | ( n2165 & n2171 ) | ( n2168 & n2171 ) ;
  assign n2280 = ( n2165 & n2168 ) | ( n2165 & ~n2171 ) | ( n2168 & ~n2171 ) ;
  assign n2281 = ( n2171 & ~n2279 ) | ( n2171 & n2280 ) | ( ~n2279 & n2280 ) ;
  assign n2282 = ( n2174 & n2177 ) | ( n2174 & n2180 ) | ( n2177 & n2180 ) ;
  assign n2283 = ( n2174 & n2177 ) | ( n2174 & ~n2180 ) | ( n2177 & ~n2180 ) ;
  assign n2284 = ( n2180 & ~n2282 ) | ( n2180 & n2283 ) | ( ~n2282 & n2283 ) ;
  assign n2285 = ( n2183 & n2281 ) | ( n2183 & n2284 ) | ( n2281 & n2284 ) ;
  assign n2286 = ( ~n2183 & n2281 ) | ( ~n2183 & n2284 ) | ( n2281 & n2284 ) ;
  assign n2287 = ( n2183 & ~n2285 ) | ( n2183 & n2286 ) | ( ~n2285 & n2286 ) ;
  assign n2288 = ( n2186 & n2278 ) | ( n2186 & n2287 ) | ( n2278 & n2287 ) ;
  assign n2289 = ( ~n2186 & n2278 ) | ( ~n2186 & n2287 ) | ( n2278 & n2287 ) ;
  assign n2290 = ( n2186 & ~n2288 ) | ( n2186 & n2289 ) | ( ~n2288 & n2289 ) ;
  assign n2291 = ( n2234 & n2269 ) | ( n2234 & n2290 ) | ( n2269 & n2290 ) ;
  assign n2292 = ( ~n2234 & n2269 ) | ( ~n2234 & n2290 ) | ( n2269 & n2290 ) ;
  assign n2293 = ( n2234 & ~n2291 ) | ( n2234 & n2292 ) | ( ~n2291 & n2292 ) ;
  assign n2294 = ( n2069 & n2072 ) | ( n2069 & n2075 ) | ( n2072 & n2075 ) ;
  assign n2295 = ( n2069 & n2072 ) | ( n2069 & ~n2075 ) | ( n2072 & ~n2075 ) ;
  assign n2296 = ( n2075 & ~n2294 ) | ( n2075 & n2295 ) | ( ~n2294 & n2295 ) ;
  assign n2297 = ( n2078 & n2081 ) | ( n2078 & n2084 ) | ( n2081 & n2084 ) ;
  assign n2298 = ( n2078 & n2081 ) | ( n2078 & ~n2084 ) | ( n2081 & ~n2084 ) ;
  assign n2299 = ( n2084 & ~n2297 ) | ( n2084 & n2298 ) | ( ~n2297 & n2298 ) ;
  assign n2300 = ( n2087 & n2296 ) | ( n2087 & n2299 ) | ( n2296 & n2299 ) ;
  assign n2301 = ( ~n2087 & n2296 ) | ( ~n2087 & n2299 ) | ( n2296 & n2299 ) ;
  assign n2302 = ( n2087 & ~n2300 ) | ( n2087 & n2301 ) | ( ~n2300 & n2301 ) ;
  assign n2303 = ( n2048 & n2051 ) | ( n2048 & n2054 ) | ( n2051 & n2054 ) ;
  assign n2304 = ( n2048 & n2051 ) | ( n2048 & ~n2054 ) | ( n2051 & ~n2054 ) ;
  assign n2305 = ( n2054 & ~n2303 ) | ( n2054 & n2304 ) | ( ~n2303 & n2304 ) ;
  assign n2306 = ( n2057 & n2060 ) | ( n2057 & n2063 ) | ( n2060 & n2063 ) ;
  assign n2307 = ( n2057 & n2060 ) | ( n2057 & ~n2063 ) | ( n2060 & ~n2063 ) ;
  assign n2308 = ( n2063 & ~n2306 ) | ( n2063 & n2307 ) | ( ~n2306 & n2307 ) ;
  assign n2309 = ( n2066 & n2305 ) | ( n2066 & n2308 ) | ( n2305 & n2308 ) ;
  assign n2310 = ( ~n2066 & n2305 ) | ( ~n2066 & n2308 ) | ( n2305 & n2308 ) ;
  assign n2311 = ( n2066 & ~n2309 ) | ( n2066 & n2310 ) | ( ~n2309 & n2310 ) ;
  assign n2312 = ( n2090 & n2302 ) | ( n2090 & n2311 ) | ( n2302 & n2311 ) ;
  assign n2313 = ( ~n2090 & n2302 ) | ( ~n2090 & n2311 ) | ( n2302 & n2311 ) ;
  assign n2314 = ( n2090 & ~n2312 ) | ( n2090 & n2313 ) | ( ~n2312 & n2313 ) ;
  assign n2315 = n1852 & n1855 ;
  assign n2316 = ( n1850 & n1853 ) | ( n1850 & n2315 ) | ( n1853 & n2315 ) ;
  assign n2317 = n2107 & ~n2315 ;
  assign n2318 = ( n2104 & ~n2108 ) | ( n2104 & n2317 ) | ( ~n2108 & n2317 ) ;
  assign n2319 = ( n2102 & n2316 ) | ( n2102 & n2318 ) | ( n2316 & n2318 ) ;
  assign n2320 = ( ~n2102 & n2316 ) | ( ~n2102 & n2318 ) | ( n2316 & n2318 ) ;
  assign n2321 = ( n2102 & ~n2319 ) | ( n2102 & n2320 ) | ( ~n2319 & n2320 ) ;
  assign n2322 = n1846 & ~n1849 ;
  assign n2323 = ( n2095 & ~n2101 ) | ( n2095 & n2322 ) | ( ~n2101 & n2322 ) ;
  assign n2324 = n1834 & n1837 ;
  assign n2325 = ( n1833 & n1836 ) | ( n1833 & n2324 ) | ( n1836 & n2324 ) ;
  assign n2326 = ( n2093 & n2323 ) | ( n2093 & n2325 ) | ( n2323 & n2325 ) ;
  assign n2327 = ( n2093 & ~n2323 ) | ( n2093 & n2325 ) | ( ~n2323 & n2325 ) ;
  assign n2328 = ( n2323 & ~n2326 ) | ( n2323 & n2327 ) | ( ~n2326 & n2327 ) ;
  assign n2329 = ( n2111 & n2321 ) | ( n2111 & n2328 ) | ( n2321 & n2328 ) ;
  assign n2330 = ( ~n2111 & n2321 ) | ( ~n2111 & n2328 ) | ( n2321 & n2328 ) ;
  assign n2331 = ( n2111 & ~n2329 ) | ( n2111 & n2330 ) | ( ~n2329 & n2330 ) ;
  assign n2332 = ( n2114 & n2117 ) | ( n2114 & n2120 ) | ( n2117 & n2120 ) ;
  assign n2333 = ( n2114 & n2117 ) | ( n2114 & ~n2120 ) | ( n2117 & ~n2120 ) ;
  assign n2334 = ( n2120 & ~n2332 ) | ( n2120 & n2333 ) | ( ~n2332 & n2333 ) ;
  assign n2335 = ( n1802 & n1805 ) | ( n1802 & n2126 ) | ( n1805 & n2126 ) ;
  assign n2336 = ( n2129 & n2132 ) | ( n2129 & n2335 ) | ( n2132 & n2335 ) ;
  assign n2337 = ( n2129 & ~n2132 ) | ( n2129 & n2335 ) | ( ~n2132 & n2335 ) ;
  assign n2338 = ( n2132 & ~n2336 ) | ( n2132 & n2337 ) | ( ~n2336 & n2337 ) ;
  assign n2339 = ( n2135 & n2334 ) | ( n2135 & n2338 ) | ( n2334 & n2338 ) ;
  assign n2340 = ( ~n2135 & n2334 ) | ( ~n2135 & n2338 ) | ( n2334 & n2338 ) ;
  assign n2341 = ( n2135 & ~n2339 ) | ( n2135 & n2340 ) | ( ~n2339 & n2340 ) ;
  assign n2342 = ( n2138 & n2331 ) | ( n2138 & n2341 ) | ( n2331 & n2341 ) ;
  assign n2343 = ( n2138 & ~n2331 ) | ( n2138 & n2341 ) | ( ~n2331 & n2341 ) ;
  assign n2344 = ( n2331 & ~n2342 ) | ( n2331 & n2343 ) | ( ~n2342 & n2343 ) ;
  assign n2345 = ( n2141 & n2314 ) | ( n2141 & n2344 ) | ( n2314 & n2344 ) ;
  assign n2346 = ( ~n2141 & n2314 ) | ( ~n2141 & n2344 ) | ( n2314 & n2344 ) ;
  assign n2347 = ( n2141 & ~n2345 ) | ( n2141 & n2346 ) | ( ~n2345 & n2346 ) ;
  assign n2348 = ( n2237 & n2293 ) | ( n2237 & n2347 ) | ( n2293 & n2347 ) ;
  assign n2349 = ( ~n2237 & n2293 ) | ( ~n2237 & n2347 ) | ( n2293 & n2347 ) ;
  assign n2350 = ( n2237 & ~n2348 ) | ( n2237 & n2349 ) | ( ~n2348 & n2349 ) ;
  assign n2351 = ( n2242 & n2244 ) | ( n2242 & n2350 ) | ( n2244 & n2350 ) ;
  assign n2352 = ( n2245 & n2248 ) | ( n2245 & n2251 ) | ( n2248 & n2251 ) ;
  assign n2353 = ( n2245 & n2248 ) | ( n2245 & ~n2251 ) | ( n2248 & ~n2251 ) ;
  assign n2354 = ( n2251 & ~n2352 ) | ( n2251 & n2353 ) | ( ~n2352 & n2353 ) ;
  assign n2355 = ( n2254 & n2261 ) | ( n2254 & n2264 ) | ( n2261 & n2264 ) ;
  assign n2356 = ( ~n2254 & n2261 ) | ( ~n2254 & n2264 ) | ( n2261 & n2264 ) ;
  assign n2357 = ( n2254 & ~n2355 ) | ( n2254 & n2356 ) | ( ~n2355 & n2356 ) ;
  assign n2358 = ( n2267 & n2354 ) | ( n2267 & n2357 ) | ( n2354 & n2357 ) ;
  assign n2359 = ( ~n2267 & n2354 ) | ( ~n2267 & n2357 ) | ( n2354 & n2357 ) ;
  assign n2360 = ( n2267 & ~n2358 ) | ( n2267 & n2359 ) | ( ~n2358 & n2359 ) ;
  assign n2361 = ( n2279 & n2282 ) | ( n2279 & n2285 ) | ( n2282 & n2285 ) ;
  assign n2362 = ( n2279 & n2282 ) | ( n2279 & ~n2285 ) | ( n2282 & ~n2285 ) ;
  assign n2363 = ( n2285 & ~n2361 ) | ( n2285 & n2362 ) | ( ~n2361 & n2362 ) ;
  assign n2364 = ( n2270 & n2273 ) | ( n2270 & n2276 ) | ( n2273 & n2276 ) ;
  assign n2365 = ( n2270 & n2273 ) | ( n2270 & ~n2276 ) | ( n2273 & ~n2276 ) ;
  assign n2366 = ( n2276 & ~n2364 ) | ( n2276 & n2365 ) | ( ~n2364 & n2365 ) ;
  assign n2367 = ( n2288 & n2363 ) | ( n2288 & n2366 ) | ( n2363 & n2366 ) ;
  assign n2368 = ( ~n2288 & n2363 ) | ( ~n2288 & n2366 ) | ( n2363 & n2366 ) ;
  assign n2369 = ( n2288 & ~n2367 ) | ( n2288 & n2368 ) | ( ~n2367 & n2368 ) ;
  assign n2370 = ( n2291 & n2360 ) | ( n2291 & n2369 ) | ( n2360 & n2369 ) ;
  assign n2371 = ( ~n2291 & n2360 ) | ( ~n2291 & n2369 ) | ( n2360 & n2369 ) ;
  assign n2372 = ( n2291 & ~n2370 ) | ( n2291 & n2371 ) | ( ~n2370 & n2371 ) ;
  assign n2373 = ( n2294 & n2297 ) | ( n2294 & n2300 ) | ( n2297 & n2300 ) ;
  assign n2374 = ( n2294 & n2297 ) | ( n2294 & ~n2300 ) | ( n2297 & ~n2300 ) ;
  assign n2375 = ( n2300 & ~n2373 ) | ( n2300 & n2374 ) | ( ~n2373 & n2374 ) ;
  assign n2376 = ( n2303 & n2306 ) | ( n2303 & n2309 ) | ( n2306 & n2309 ) ;
  assign n2377 = ( n2303 & n2306 ) | ( n2303 & ~n2309 ) | ( n2306 & ~n2309 ) ;
  assign n2378 = ( n2309 & ~n2376 ) | ( n2309 & n2377 ) | ( ~n2376 & n2377 ) ;
  assign n2379 = ( n2312 & n2375 ) | ( n2312 & n2378 ) | ( n2375 & n2378 ) ;
  assign n2380 = ( ~n2312 & n2375 ) | ( ~n2312 & n2378 ) | ( n2375 & n2378 ) ;
  assign n2381 = ( n2312 & ~n2379 ) | ( n2312 & n2380 ) | ( ~n2379 & n2380 ) ;
  assign n2382 = ( n2319 & n2326 ) | ( n2319 & n2329 ) | ( n2326 & n2329 ) ;
  assign n2383 = ( n2319 & n2326 ) | ( n2319 & ~n2329 ) | ( n2326 & ~n2329 ) ;
  assign n2384 = ( n2329 & ~n2382 ) | ( n2329 & n2383 ) | ( ~n2382 & n2383 ) ;
  assign n2385 = ( n2332 & n2336 ) | ( n2332 & n2339 ) | ( n2336 & n2339 ) ;
  assign n2386 = ( n2332 & ~n2336 ) | ( n2332 & n2339 ) | ( ~n2336 & n2339 ) ;
  assign n2387 = ( n2336 & ~n2385 ) | ( n2336 & n2386 ) | ( ~n2385 & n2386 ) ;
  assign n2388 = ( n2342 & n2384 ) | ( n2342 & n2387 ) | ( n2384 & n2387 ) ;
  assign n2389 = ( ~n2342 & n2384 ) | ( ~n2342 & n2387 ) | ( n2384 & n2387 ) ;
  assign n2390 = ( n2342 & ~n2388 ) | ( n2342 & n2389 ) | ( ~n2388 & n2389 ) ;
  assign n2391 = ( n2345 & n2381 ) | ( n2345 & n2390 ) | ( n2381 & n2390 ) ;
  assign n2392 = ( ~n2345 & n2381 ) | ( ~n2345 & n2390 ) | ( n2381 & n2390 ) ;
  assign n2393 = ( n2345 & ~n2391 ) | ( n2345 & n2392 ) | ( ~n2391 & n2392 ) ;
  assign n2394 = ( n2348 & n2372 ) | ( n2348 & n2393 ) | ( n2372 & n2393 ) ;
  assign n2395 = ( ~n2348 & n2372 ) | ( ~n2348 & n2393 ) | ( n2372 & n2393 ) ;
  assign n2396 = ( n2348 & ~n2394 ) | ( n2348 & n2395 ) | ( ~n2394 & n2395 ) ;
  assign n2397 = ( ~n1639 & n1660 ) | ( ~n1639 & n1681 ) | ( n1660 & n1681 ) ;
  assign n2398 = ( n1639 & ~n1682 ) | ( n1639 & n2397 ) | ( ~n1682 & n2397 ) ;
  assign n2399 = ( n2351 & n2396 ) | ( n2351 & n2398 ) | ( n2396 & n2398 ) ;
  assign n2400 = ( ~n1682 & n1691 ) | ( ~n1682 & n1700 ) | ( n1691 & n1700 ) ;
  assign n2401 = ( n1682 & ~n1701 ) | ( n1682 & n2400 ) | ( ~n1701 & n2400 ) ;
  assign n2402 = ( n2373 & n2376 ) | ( n2373 & n2379 ) | ( n2376 & n2379 ) ;
  assign n2403 = ( n2373 & n2376 ) | ( n2373 & ~n2379 ) | ( n2376 & ~n2379 ) ;
  assign n2404 = ( n2379 & ~n2402 ) | ( n2379 & n2403 ) | ( ~n2402 & n2403 ) ;
  assign n2405 = ( n2382 & n2385 ) | ( n2382 & n2388 ) | ( n2385 & n2388 ) ;
  assign n2406 = ( n2382 & n2385 ) | ( n2382 & ~n2388 ) | ( n2385 & ~n2388 ) ;
  assign n2407 = ( n2388 & ~n2405 ) | ( n2388 & n2406 ) | ( ~n2405 & n2406 ) ;
  assign n2408 = ( n2391 & n2404 ) | ( n2391 & n2407 ) | ( n2404 & n2407 ) ;
  assign n2409 = ( ~n2391 & n2404 ) | ( ~n2391 & n2407 ) | ( n2404 & n2407 ) ;
  assign n2410 = ( n2391 & ~n2408 ) | ( n2391 & n2409 ) | ( ~n2408 & n2409 ) ;
  assign n2411 = ( n2361 & n2364 ) | ( n2361 & n2367 ) | ( n2364 & n2367 ) ;
  assign n2412 = ( n2361 & n2364 ) | ( n2361 & ~n2367 ) | ( n2364 & ~n2367 ) ;
  assign n2413 = ( n2367 & ~n2411 ) | ( n2367 & n2412 ) | ( ~n2411 & n2412 ) ;
  assign n2414 = ( n2352 & n2355 ) | ( n2352 & n2358 ) | ( n2355 & n2358 ) ;
  assign n2415 = ( n2352 & n2355 ) | ( n2352 & ~n2358 ) | ( n2355 & ~n2358 ) ;
  assign n2416 = ( n2358 & ~n2414 ) | ( n2358 & n2415 ) | ( ~n2414 & n2415 ) ;
  assign n2417 = ( n2370 & n2413 ) | ( n2370 & n2416 ) | ( n2413 & n2416 ) ;
  assign n2418 = ( ~n2370 & n2413 ) | ( ~n2370 & n2416 ) | ( n2413 & n2416 ) ;
  assign n2419 = ( n2370 & ~n2417 ) | ( n2370 & n2418 ) | ( ~n2417 & n2418 ) ;
  assign n2420 = ( n2394 & n2410 ) | ( n2394 & n2419 ) | ( n2410 & n2419 ) ;
  assign n2421 = ( ~n2394 & n2410 ) | ( ~n2394 & n2419 ) | ( n2410 & n2419 ) ;
  assign n2422 = ( n2394 & ~n2420 ) | ( n2394 & n2421 ) | ( ~n2420 & n2421 ) ;
  assign n2423 = ( n2399 & n2401 ) | ( n2399 & n2422 ) | ( n2401 & n2422 ) ;
  assign n2424 = ( ~n1701 & n1704 ) | ( ~n1701 & n1707 ) | ( n1704 & n1707 ) ;
  assign n2425 = ( n1701 & ~n1708 ) | ( n1701 & n2424 ) | ( ~n1708 & n2424 ) ;
  assign n2426 = ( n2402 & n2405 ) | ( n2402 & n2408 ) | ( n2405 & n2408 ) ;
  assign n2427 = ( n2402 & n2405 ) | ( n2402 & ~n2408 ) | ( n2405 & ~n2408 ) ;
  assign n2428 = ( n2408 & ~n2426 ) | ( n2408 & n2427 ) | ( ~n2426 & n2427 ) ;
  assign n2429 = ( n2411 & n2414 ) | ( n2411 & n2417 ) | ( n2414 & n2417 ) ;
  assign n2430 = ( ~n2411 & n2414 ) | ( ~n2411 & n2417 ) | ( n2414 & n2417 ) ;
  assign n2431 = ( n2411 & ~n2429 ) | ( n2411 & n2430 ) | ( ~n2429 & n2430 ) ;
  assign n2432 = ( n2420 & n2428 ) | ( n2420 & n2431 ) | ( n2428 & n2431 ) ;
  assign n2433 = ( ~n2420 & n2428 ) | ( ~n2420 & n2431 ) | ( n2428 & n2431 ) ;
  assign n2434 = ( n2420 & ~n2432 ) | ( n2420 & n2433 ) | ( ~n2432 & n2433 ) ;
  assign n2435 = ( n2423 & n2425 ) | ( n2423 & n2434 ) | ( n2425 & n2434 ) ;
  assign n2436 = ( n2426 & n2429 ) | ( n2426 & n2432 ) | ( n2429 & n2432 ) ;
  assign n2437 = ( n2426 & n2429 ) | ( n2426 & ~n2432 ) | ( n2429 & ~n2432 ) ;
  assign n2438 = ( n2432 & ~n2436 ) | ( n2432 & n2437 ) | ( ~n2436 & n2437 ) ;
  assign n2439 = ( n1711 & n2435 ) | ( n1711 & n2438 ) | ( n2435 & n2438 ) ;
  assign n2440 = ( n1709 & n2436 ) | ( n1709 & n2439 ) | ( n2436 & n2439 ) ;
  assign n2441 = ( n1709 & n2436 ) | ( n1709 & ~n2439 ) | ( n2436 & ~n2439 ) ;
  assign n2442 = ( n2439 & ~n2440 ) | ( n2439 & n2441 ) | ( ~n2440 & n2441 ) ;
  assign n2443 = ( x85 & x86 ) | ( x85 & x87 ) | ( x86 & x87 ) ;
  assign n2444 = ( x88 & x89 ) | ( x88 & x90 ) | ( x89 & x90 ) ;
  assign n2445 = ( ~x85 & x86 ) | ( ~x85 & x87 ) | ( x86 & x87 ) ;
  assign n2446 = ( x85 & ~n2443 ) | ( x85 & n2445 ) | ( ~n2443 & n2445 ) ;
  assign n2447 = ( ~x88 & x89 ) | ( ~x88 & x90 ) | ( x89 & x90 ) ;
  assign n2448 = ( x88 & ~n2444 ) | ( x88 & n2447 ) | ( ~n2444 & n2447 ) ;
  assign n2449 = n2446 & n2448 ;
  assign n2450 = ( n2443 & n2444 ) | ( n2443 & n2449 ) | ( n2444 & n2449 ) ;
  assign n2451 = ( x79 & x80 ) | ( x79 & x81 ) | ( x80 & x81 ) ;
  assign n2452 = ( x82 & x83 ) | ( x82 & x84 ) | ( x83 & x84 ) ;
  assign n2453 = ( ~x79 & x80 ) | ( ~x79 & x81 ) | ( x80 & x81 ) ;
  assign n2454 = ( x79 & ~n2451 ) | ( x79 & n2453 ) | ( ~n2451 & n2453 ) ;
  assign n2455 = ( ~x82 & x83 ) | ( ~x82 & x84 ) | ( x83 & x84 ) ;
  assign n2456 = ( x82 & ~n2452 ) | ( x82 & n2455 ) | ( ~n2452 & n2455 ) ;
  assign n2457 = n2454 & n2456 ;
  assign n2458 = ( n2451 & n2452 ) | ( n2451 & n2457 ) | ( n2452 & n2457 ) ;
  assign n2459 = n2443 | n2444 ;
  assign n2460 = n2443 & n2444 ;
  assign n2461 = n2459 & ~n2460 ;
  assign n2462 = ~n2449 & n2461 ;
  assign n2463 = n2454 | n2456 ;
  assign n2464 = ~n2457 & n2463 ;
  assign n2465 = ( n2446 & n2448 ) | ( n2446 & n2464 ) | ( n2448 & n2464 ) ;
  assign n2466 = ( ~n2451 & n2452 ) | ( ~n2451 & n2457 ) | ( n2452 & n2457 ) ;
  assign n2467 = ( n2451 & ~n2458 ) | ( n2451 & n2466 ) | ( ~n2458 & n2466 ) ;
  assign n2468 = ( n2461 & n2465 ) | ( n2461 & n2467 ) | ( n2465 & n2467 ) ;
  assign n2469 = ( ~n2461 & n2462 ) | ( ~n2461 & n2468 ) | ( n2462 & n2468 ) ;
  assign n2470 = ( n2450 & n2458 ) | ( n2450 & n2469 ) | ( n2458 & n2469 ) ;
  assign n2471 = x91 | x92 ;
  assign n2472 = ~x91 & x92 ;
  assign n2473 = ( ~x92 & n2471 ) | ( ~x92 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2474 = ( x93 & x96 ) | ( x93 & ~n2473 ) | ( x96 & ~n2473 ) ;
  assign n2475 = ( x93 & x96 ) | ( x93 & n2473 ) | ( x96 & n2473 ) ;
  assign n2476 = ( n2473 & n2474 ) | ( n2473 & ~n2475 ) | ( n2474 & ~n2475 ) ;
  assign n2477 = ( x94 & x95 ) | ( x94 & n2476 ) | ( x95 & n2476 ) ;
  assign n2478 = ( x92 & x93 ) | ( x92 & x96 ) | ( x93 & x96 ) ;
  assign n2479 = x91 & ~n2476 ;
  assign n2480 = ( n2477 & n2478 ) | ( n2477 & n2479 ) | ( n2478 & n2479 ) ;
  assign n2481 = ( x97 & x98 ) | ( x97 & x99 ) | ( x98 & x99 ) ;
  assign n2482 = ( x100 & x101 ) | ( x100 & x102 ) | ( x101 & x102 ) ;
  assign n2483 = ( ~n2477 & n2478 ) | ( ~n2477 & n2479 ) | ( n2478 & n2479 ) ;
  assign n2484 = ( n2477 & ~n2480 ) | ( n2477 & n2483 ) | ( ~n2480 & n2483 ) ;
  assign n2485 = ( n2481 & n2482 ) | ( n2481 & n2484 ) | ( n2482 & n2484 ) ;
  assign n2486 = ( ~x94 & x95 ) | ( ~x94 & n2476 ) | ( x95 & n2476 ) ;
  assign n2487 = ( x94 & ~n2477 ) | ( x94 & n2486 ) | ( ~n2477 & n2486 ) ;
  assign n2488 = ( ~x97 & x98 ) | ( ~x97 & x99 ) | ( x98 & x99 ) ;
  assign n2489 = ( x97 & ~n2481 ) | ( x97 & n2488 ) | ( ~n2481 & n2488 ) ;
  assign n2490 = ( ~x100 & x101 ) | ( ~x100 & x102 ) | ( x101 & x102 ) ;
  assign n2491 = ( x100 & ~n2482 ) | ( x100 & n2490 ) | ( ~n2482 & n2490 ) ;
  assign n2492 = ( n2487 & n2489 ) | ( n2487 & n2491 ) | ( n2489 & n2491 ) ;
  assign n2493 = ( n2481 & n2482 ) | ( n2481 & ~n2484 ) | ( n2482 & ~n2484 ) ;
  assign n2494 = ( n2484 & ~n2485 ) | ( n2484 & n2493 ) | ( ~n2485 & n2493 ) ;
  assign n2495 = n2492 & n2494 ;
  assign n2496 = ( n2480 & n2485 ) | ( n2480 & n2495 ) | ( n2485 & n2495 ) ;
  assign n2497 = n2492 | n2494 ;
  assign n2498 = ~n2495 & n2497 ;
  assign n2499 = ( ~n2487 & n2489 ) | ( ~n2487 & n2491 ) | ( n2489 & n2491 ) ;
  assign n2500 = ( n2487 & ~n2492 ) | ( n2487 & n2499 ) | ( ~n2492 & n2499 ) ;
  assign n2501 = ( n2446 & n2448 ) | ( n2446 & ~n2464 ) | ( n2448 & ~n2464 ) ;
  assign n2502 = ( n2464 & ~n2465 ) | ( n2464 & n2501 ) | ( ~n2465 & n2501 ) ;
  assign n2503 = n2500 & n2502 ;
  assign n2504 = ( ~n2461 & n2465 ) | ( ~n2461 & n2467 ) | ( n2465 & n2467 ) ;
  assign n2505 = ( n2462 & ~n2469 ) | ( n2462 & n2504 ) | ( ~n2469 & n2504 ) ;
  assign n2506 = ( n2498 & n2503 ) | ( n2498 & n2505 ) | ( n2503 & n2505 ) ;
  assign n2507 = ( n2450 & ~n2458 ) | ( n2450 & n2469 ) | ( ~n2458 & n2469 ) ;
  assign n2508 = ( n2458 & ~n2470 ) | ( n2458 & n2507 ) | ( ~n2470 & n2507 ) ;
  assign n2509 = ( ~n2480 & n2485 ) | ( ~n2480 & n2495 ) | ( n2485 & n2495 ) ;
  assign n2510 = ( n2480 & ~n2496 ) | ( n2480 & n2509 ) | ( ~n2496 & n2509 ) ;
  assign n2511 = ( n2506 & n2508 ) | ( n2506 & n2510 ) | ( n2508 & n2510 ) ;
  assign n2512 = ( n2470 & n2496 ) | ( n2470 & n2511 ) | ( n2496 & n2511 ) ;
  assign n2513 = ( x118 & x119 ) | ( x118 & x120 ) | ( x119 & x120 ) ;
  assign n2514 = ( x115 & x116 ) | ( x115 & x117 ) | ( x116 & x117 ) ;
  assign n2515 = ( ~x118 & x119 ) | ( ~x118 & x120 ) | ( x119 & x120 ) ;
  assign n2516 = ( x118 & ~n2513 ) | ( x118 & n2515 ) | ( ~n2513 & n2515 ) ;
  assign n2517 = ( ~x115 & x116 ) | ( ~x115 & x117 ) | ( x116 & x117 ) ;
  assign n2518 = ( x115 & ~n2514 ) | ( x115 & n2517 ) | ( ~n2514 & n2517 ) ;
  assign n2519 = n2516 & n2518 ;
  assign n2520 = ( n2513 & n2514 ) | ( n2513 & n2519 ) | ( n2514 & n2519 ) ;
  assign n2521 = ( x124 & x125 ) | ( x124 & x126 ) | ( x125 & x126 ) ;
  assign n2522 = ( x121 & x122 ) | ( x121 & x123 ) | ( x122 & x123 ) ;
  assign n2523 = n2521 & n2522 ;
  assign n2524 = n2516 | n2518 ;
  assign n2525 = ~n2519 & n2524 ;
  assign n2526 = ( ~x124 & x125 ) | ( ~x124 & x126 ) | ( x125 & x126 ) ;
  assign n2527 = ( x124 & ~n2521 ) | ( x124 & n2526 ) | ( ~n2521 & n2526 ) ;
  assign n2528 = ( ~x121 & x122 ) | ( ~x121 & x123 ) | ( x122 & x123 ) ;
  assign n2529 = ( x121 & ~n2522 ) | ( x121 & n2528 ) | ( ~n2522 & n2528 ) ;
  assign n2530 = ( n2525 & n2527 ) | ( n2525 & n2529 ) | ( n2527 & n2529 ) ;
  assign n2531 = ( ~n2513 & n2514 ) | ( ~n2513 & n2519 ) | ( n2514 & n2519 ) ;
  assign n2532 = ( n2513 & ~n2520 ) | ( n2513 & n2531 ) | ( ~n2520 & n2531 ) ;
  assign n2533 = n2521 | n2522 ;
  assign n2534 = ~n2523 & n2533 ;
  assign n2535 = ( n2530 & n2532 ) | ( n2530 & n2534 ) | ( n2532 & n2534 ) ;
  assign n2536 = ( n2520 & n2523 ) | ( n2520 & n2535 ) | ( n2523 & n2535 ) ;
  assign n2537 = ( x106 & x107 ) | ( x106 & x108 ) | ( x107 & x108 ) ;
  assign n2538 = ( x103 & x104 ) | ( x103 & x105 ) | ( x104 & x105 ) ;
  assign n2539 = ( ~x106 & x107 ) | ( ~x106 & x108 ) | ( x107 & x108 ) ;
  assign n2540 = ( x106 & ~n2537 ) | ( x106 & n2539 ) | ( ~n2537 & n2539 ) ;
  assign n2541 = ( ~x103 & x104 ) | ( ~x103 & x105 ) | ( x104 & x105 ) ;
  assign n2542 = ( x103 & ~n2538 ) | ( x103 & n2541 ) | ( ~n2538 & n2541 ) ;
  assign n2543 = n2540 & n2542 ;
  assign n2544 = ( n2537 & n2538 ) | ( n2537 & n2543 ) | ( n2538 & n2543 ) ;
  assign n2545 = ( x112 & x113 ) | ( x112 & x114 ) | ( x113 & x114 ) ;
  assign n2546 = ( x109 & x110 ) | ( x109 & x111 ) | ( x110 & x111 ) ;
  assign n2547 = n2545 & n2546 ;
  assign n2548 = n2540 | n2542 ;
  assign n2549 = ~n2543 & n2548 ;
  assign n2550 = ( ~x112 & x113 ) | ( ~x112 & x114 ) | ( x113 & x114 ) ;
  assign n2551 = ( x112 & ~n2545 ) | ( x112 & n2550 ) | ( ~n2545 & n2550 ) ;
  assign n2552 = ( ~x109 & x110 ) | ( ~x109 & x111 ) | ( x110 & x111 ) ;
  assign n2553 = ( x109 & ~n2546 ) | ( x109 & n2552 ) | ( ~n2546 & n2552 ) ;
  assign n2554 = ( n2549 & n2551 ) | ( n2549 & n2553 ) | ( n2551 & n2553 ) ;
  assign n2555 = ( ~n2537 & n2538 ) | ( ~n2537 & n2543 ) | ( n2538 & n2543 ) ;
  assign n2556 = ( n2537 & ~n2544 ) | ( n2537 & n2555 ) | ( ~n2544 & n2555 ) ;
  assign n2557 = n2545 | n2546 ;
  assign n2558 = ~n2547 & n2557 ;
  assign n2559 = ( n2554 & n2556 ) | ( n2554 & n2558 ) | ( n2556 & n2558 ) ;
  assign n2560 = ( n2544 & n2547 ) | ( n2544 & n2559 ) | ( n2547 & n2559 ) ;
  assign n2561 = ( ~n2525 & n2527 ) | ( ~n2525 & n2529 ) | ( n2527 & n2529 ) ;
  assign n2562 = ( n2525 & ~n2530 ) | ( n2525 & n2561 ) | ( ~n2530 & n2561 ) ;
  assign n2563 = ( ~n2549 & n2551 ) | ( ~n2549 & n2553 ) | ( n2551 & n2553 ) ;
  assign n2564 = ( n2549 & ~n2554 ) | ( n2549 & n2563 ) | ( ~n2554 & n2563 ) ;
  assign n2565 = n2562 & n2564 ;
  assign n2566 = ( ~n2530 & n2532 ) | ( ~n2530 & n2534 ) | ( n2532 & n2534 ) ;
  assign n2567 = ( n2530 & ~n2535 ) | ( n2530 & n2566 ) | ( ~n2535 & n2566 ) ;
  assign n2568 = ( ~n2554 & n2556 ) | ( ~n2554 & n2558 ) | ( n2556 & n2558 ) ;
  assign n2569 = ( n2554 & ~n2559 ) | ( n2554 & n2568 ) | ( ~n2559 & n2568 ) ;
  assign n2570 = ( n2565 & n2567 ) | ( n2565 & n2569 ) | ( n2567 & n2569 ) ;
  assign n2571 = ( n2520 & n2523 ) | ( n2520 & ~n2535 ) | ( n2523 & ~n2535 ) ;
  assign n2572 = ( n2535 & ~n2536 ) | ( n2535 & n2571 ) | ( ~n2536 & n2571 ) ;
  assign n2573 = ( n2544 & n2547 ) | ( n2544 & ~n2559 ) | ( n2547 & ~n2559 ) ;
  assign n2574 = ( n2559 & ~n2560 ) | ( n2559 & n2573 ) | ( ~n2560 & n2573 ) ;
  assign n2575 = ( n2570 & n2572 ) | ( n2570 & n2574 ) | ( n2572 & n2574 ) ;
  assign n2576 = ( n2536 & n2560 ) | ( n2536 & n2575 ) | ( n2560 & n2575 ) ;
  assign n2577 = ( ~n2498 & n2503 ) | ( ~n2498 & n2505 ) | ( n2503 & n2505 ) ;
  assign n2578 = ( n2498 & ~n2506 ) | ( n2498 & n2577 ) | ( ~n2506 & n2577 ) ;
  assign n2579 = ( ~n2565 & n2567 ) | ( ~n2565 & n2569 ) | ( n2567 & n2569 ) ;
  assign n2580 = ( n2565 & ~n2570 ) | ( n2565 & n2579 ) | ( ~n2570 & n2579 ) ;
  assign n2581 = n2562 | n2564 ;
  assign n2582 = ~n2565 & n2581 ;
  assign n2583 = ( n2500 & n2502 ) | ( n2500 & n2582 ) | ( n2502 & n2582 ) ;
  assign n2584 = ~n2503 & n2583 ;
  assign n2585 = ( n2578 & n2580 ) | ( n2578 & n2584 ) | ( n2580 & n2584 ) ;
  assign n2586 = ( ~n2506 & n2508 ) | ( ~n2506 & n2510 ) | ( n2508 & n2510 ) ;
  assign n2587 = ( n2506 & ~n2511 ) | ( n2506 & n2586 ) | ( ~n2511 & n2586 ) ;
  assign n2588 = ( ~n2570 & n2572 ) | ( ~n2570 & n2574 ) | ( n2572 & n2574 ) ;
  assign n2589 = ( n2570 & ~n2575 ) | ( n2570 & n2588 ) | ( ~n2575 & n2588 ) ;
  assign n2590 = ( n2585 & n2587 ) | ( n2585 & n2589 ) | ( n2587 & n2589 ) ;
  assign n2591 = ( n2470 & n2496 ) | ( n2470 & ~n2511 ) | ( n2496 & ~n2511 ) ;
  assign n2592 = ( n2511 & ~n2512 ) | ( n2511 & n2591 ) | ( ~n2512 & n2591 ) ;
  assign n2593 = ( ~n2536 & n2560 ) | ( ~n2536 & n2575 ) | ( n2560 & n2575 ) ;
  assign n2594 = ( n2536 & ~n2576 ) | ( n2536 & n2593 ) | ( ~n2576 & n2593 ) ;
  assign n2595 = ( n2590 & n2592 ) | ( n2590 & n2594 ) | ( n2592 & n2594 ) ;
  assign n2596 = ( n2512 & n2576 ) | ( n2512 & n2595 ) | ( n2576 & n2595 ) ;
  assign n2597 = ( x172 & x173 ) | ( x172 & x174 ) | ( x173 & x174 ) ;
  assign n2598 = ( x169 & x170 ) | ( x169 & x171 ) | ( x170 & x171 ) ;
  assign n2599 = ( ~x163 & x164 ) | ( ~x163 & x165 ) | ( x164 & x165 ) ;
  assign n2600 = ( x163 & x164 ) | ( x163 & x165 ) | ( x164 & x165 ) ;
  assign n2601 = ( x163 & n2599 ) | ( x163 & ~n2600 ) | ( n2599 & ~n2600 ) ;
  assign n2602 = ( ~x166 & x167 ) | ( ~x166 & x168 ) | ( x167 & x168 ) ;
  assign n2603 = ( x166 & x167 ) | ( x166 & x168 ) | ( x167 & x168 ) ;
  assign n2604 = ( x166 & n2602 ) | ( x166 & ~n2603 ) | ( n2602 & ~n2603 ) ;
  assign n2605 = n2601 | n2604 ;
  assign n2606 = n2601 & n2604 ;
  assign n2607 = n2605 & ~n2606 ;
  assign n2608 = ( ~x172 & x173 ) | ( ~x172 & x174 ) | ( x173 & x174 ) ;
  assign n2609 = ( x172 & ~n2597 ) | ( x172 & n2608 ) | ( ~n2597 & n2608 ) ;
  assign n2610 = ( ~x169 & x170 ) | ( ~x169 & x171 ) | ( x170 & x171 ) ;
  assign n2611 = ( x169 & ~n2598 ) | ( x169 & n2610 ) | ( ~n2598 & n2610 ) ;
  assign n2612 = ( n2607 & n2609 ) | ( n2607 & n2611 ) | ( n2609 & n2611 ) ;
  assign n2613 = ( n2597 & n2598 ) | ( n2597 & n2612 ) | ( n2598 & n2612 ) ;
  assign n2614 = ( n2600 & n2603 ) | ( n2600 & n2606 ) | ( n2603 & n2606 ) ;
  assign n2615 = ( n2597 & n2598 ) | ( n2597 & ~n2612 ) | ( n2598 & ~n2612 ) ;
  assign n2616 = ( n2612 & ~n2613 ) | ( n2612 & n2615 ) | ( ~n2613 & n2615 ) ;
  assign n2617 = ( ~n2600 & n2603 ) | ( ~n2600 & n2606 ) | ( n2603 & n2606 ) ;
  assign n2618 = ( n2600 & ~n2614 ) | ( n2600 & n2617 ) | ( ~n2614 & n2617 ) ;
  assign n2619 = n2616 & n2618 ;
  assign n2620 = ( n2613 & n2614 ) | ( n2613 & n2619 ) | ( n2614 & n2619 ) ;
  assign n2621 = ( x151 & x152 ) | ( x151 & x153 ) | ( x152 & x153 ) ;
  assign n2622 = ( x154 & x155 ) | ( x154 & x156 ) | ( x155 & x156 ) ;
  assign n2623 = ( ~x151 & x152 ) | ( ~x151 & x153 ) | ( x152 & x153 ) ;
  assign n2624 = ( x151 & ~n2621 ) | ( x151 & n2623 ) | ( ~n2621 & n2623 ) ;
  assign n2625 = ( ~x154 & x155 ) | ( ~x154 & x156 ) | ( x155 & x156 ) ;
  assign n2626 = ( x154 & ~n2622 ) | ( x154 & n2625 ) | ( ~n2622 & n2625 ) ;
  assign n2627 = n2624 & n2626 ;
  assign n2628 = ( n2621 & n2622 ) | ( n2621 & n2627 ) | ( n2622 & n2627 ) ;
  assign n2629 = ( x157 & x158 ) | ( x157 & x159 ) | ( x158 & x159 ) ;
  assign n2630 = ( x160 & x161 ) | ( x160 & x162 ) | ( x161 & x162 ) ;
  assign n2631 = n2629 & n2630 ;
  assign n2632 = n2624 | n2626 ;
  assign n2633 = ~n2627 & n2632 ;
  assign n2634 = ( ~x157 & x158 ) | ( ~x157 & x159 ) | ( x158 & x159 ) ;
  assign n2635 = ( x157 & ~n2629 ) | ( x157 & n2634 ) | ( ~n2629 & n2634 ) ;
  assign n2636 = ( ~x160 & x161 ) | ( ~x160 & x162 ) | ( x161 & x162 ) ;
  assign n2637 = ( x160 & ~n2630 ) | ( x160 & n2636 ) | ( ~n2630 & n2636 ) ;
  assign n2638 = ( n2633 & n2635 ) | ( n2633 & n2637 ) | ( n2635 & n2637 ) ;
  assign n2639 = ( ~n2621 & n2622 ) | ( ~n2621 & n2627 ) | ( n2622 & n2627 ) ;
  assign n2640 = ( n2621 & ~n2628 ) | ( n2621 & n2639 ) | ( ~n2628 & n2639 ) ;
  assign n2641 = n2629 | n2630 ;
  assign n2642 = ~n2631 & n2641 ;
  assign n2643 = ( n2638 & n2640 ) | ( n2638 & n2642 ) | ( n2640 & n2642 ) ;
  assign n2644 = ( n2628 & n2631 ) | ( n2628 & n2643 ) | ( n2631 & n2643 ) ;
  assign n2645 = ( ~n2633 & n2635 ) | ( ~n2633 & n2637 ) | ( n2635 & n2637 ) ;
  assign n2646 = ( n2633 & ~n2638 ) | ( n2633 & n2645 ) | ( ~n2638 & n2645 ) ;
  assign n2647 = ( ~n2607 & n2609 ) | ( ~n2607 & n2611 ) | ( n2609 & n2611 ) ;
  assign n2648 = ( n2607 & ~n2612 ) | ( n2607 & n2647 ) | ( ~n2612 & n2647 ) ;
  assign n2649 = n2646 & n2648 ;
  assign n2650 = ( ~n2638 & n2640 ) | ( ~n2638 & n2642 ) | ( n2640 & n2642 ) ;
  assign n2651 = ( n2638 & ~n2643 ) | ( n2638 & n2650 ) | ( ~n2643 & n2650 ) ;
  assign n2652 = n2616 | n2618 ;
  assign n2653 = ~n2619 & n2652 ;
  assign n2654 = ( n2649 & n2651 ) | ( n2649 & n2653 ) | ( n2651 & n2653 ) ;
  assign n2655 = ( ~n2613 & n2614 ) | ( ~n2613 & n2619 ) | ( n2614 & n2619 ) ;
  assign n2656 = ( n2613 & ~n2620 ) | ( n2613 & n2655 ) | ( ~n2620 & n2655 ) ;
  assign n2657 = ( n2628 & n2631 ) | ( n2628 & ~n2643 ) | ( n2631 & ~n2643 ) ;
  assign n2658 = ( n2643 & ~n2644 ) | ( n2643 & n2657 ) | ( ~n2644 & n2657 ) ;
  assign n2659 = ( n2654 & n2656 ) | ( n2654 & n2658 ) | ( n2656 & n2658 ) ;
  assign n2660 = ( n2620 & n2644 ) | ( n2620 & n2659 ) | ( n2644 & n2659 ) ;
  assign n2661 = ( x127 & x128 ) | ( x127 & x129 ) | ( x128 & x129 ) ;
  assign n2662 = ( x130 & x131 ) | ( x130 & x132 ) | ( x131 & x132 ) ;
  assign n2663 = ( ~x127 & x128 ) | ( ~x127 & x129 ) | ( x128 & x129 ) ;
  assign n2664 = ( x127 & ~n2661 ) | ( x127 & n2663 ) | ( ~n2661 & n2663 ) ;
  assign n2665 = ( ~x130 & x131 ) | ( ~x130 & x132 ) | ( x131 & x132 ) ;
  assign n2666 = ( x130 & ~n2662 ) | ( x130 & n2665 ) | ( ~n2662 & n2665 ) ;
  assign n2667 = n2664 & n2666 ;
  assign n2668 = ( n2661 & n2662 ) | ( n2661 & n2667 ) | ( n2662 & n2667 ) ;
  assign n2669 = ( x136 & x137 ) | ( x136 & x138 ) | ( x137 & x138 ) ;
  assign n2670 = ( x133 & x134 ) | ( x133 & x135 ) | ( x134 & x135 ) ;
  assign n2671 = n2669 & n2670 ;
  assign n2672 = n2664 | n2666 ;
  assign n2673 = ~n2667 & n2672 ;
  assign n2674 = ( ~x136 & x137 ) | ( ~x136 & x138 ) | ( x137 & x138 ) ;
  assign n2675 = ( x136 & ~n2669 ) | ( x136 & n2674 ) | ( ~n2669 & n2674 ) ;
  assign n2676 = ( ~x133 & x134 ) | ( ~x133 & x135 ) | ( x134 & x135 ) ;
  assign n2677 = ( x133 & ~n2670 ) | ( x133 & n2676 ) | ( ~n2670 & n2676 ) ;
  assign n2678 = ( n2673 & n2675 ) | ( n2673 & n2677 ) | ( n2675 & n2677 ) ;
  assign n2679 = ( ~n2661 & n2662 ) | ( ~n2661 & n2667 ) | ( n2662 & n2667 ) ;
  assign n2680 = ( n2661 & ~n2668 ) | ( n2661 & n2679 ) | ( ~n2668 & n2679 ) ;
  assign n2681 = n2669 | n2670 ;
  assign n2682 = ~n2671 & n2681 ;
  assign n2683 = ( n2678 & n2680 ) | ( n2678 & n2682 ) | ( n2680 & n2682 ) ;
  assign n2684 = ( n2668 & n2671 ) | ( n2668 & n2683 ) | ( n2671 & n2683 ) ;
  assign n2685 = ( x142 & x143 ) | ( x142 & x144 ) | ( x143 & x144 ) ;
  assign n2686 = ( x139 & x140 ) | ( x139 & x141 ) | ( x140 & x141 ) ;
  assign n2687 = ( ~x142 & x143 ) | ( ~x142 & x144 ) | ( x143 & x144 ) ;
  assign n2688 = ( x142 & ~n2685 ) | ( x142 & n2687 ) | ( ~n2685 & n2687 ) ;
  assign n2689 = ( ~x139 & x140 ) | ( ~x139 & x141 ) | ( x140 & x141 ) ;
  assign n2690 = ( x139 & ~n2686 ) | ( x139 & n2689 ) | ( ~n2686 & n2689 ) ;
  assign n2691 = n2688 & n2690 ;
  assign n2692 = ( n2685 & n2686 ) | ( n2685 & n2691 ) | ( n2686 & n2691 ) ;
  assign n2693 = ( x148 & x149 ) | ( x148 & x150 ) | ( x149 & x150 ) ;
  assign n2694 = ( x145 & x146 ) | ( x145 & x147 ) | ( x146 & x147 ) ;
  assign n2695 = n2693 & n2694 ;
  assign n2696 = n2688 | n2690 ;
  assign n2697 = ~n2691 & n2696 ;
  assign n2698 = ( ~x148 & x149 ) | ( ~x148 & x150 ) | ( x149 & x150 ) ;
  assign n2699 = ( x148 & ~n2693 ) | ( x148 & n2698 ) | ( ~n2693 & n2698 ) ;
  assign n2700 = ( ~x145 & x146 ) | ( ~x145 & x147 ) | ( x146 & x147 ) ;
  assign n2701 = ( x145 & ~n2694 ) | ( x145 & n2700 ) | ( ~n2694 & n2700 ) ;
  assign n2702 = ( n2697 & n2699 ) | ( n2697 & n2701 ) | ( n2699 & n2701 ) ;
  assign n2703 = ( ~n2685 & n2686 ) | ( ~n2685 & n2691 ) | ( n2686 & n2691 ) ;
  assign n2704 = ( n2685 & ~n2692 ) | ( n2685 & n2703 ) | ( ~n2692 & n2703 ) ;
  assign n2705 = n2693 | n2694 ;
  assign n2706 = ~n2695 & n2705 ;
  assign n2707 = ( n2702 & n2704 ) | ( n2702 & n2706 ) | ( n2704 & n2706 ) ;
  assign n2708 = ( n2692 & n2695 ) | ( n2692 & n2707 ) | ( n2695 & n2707 ) ;
  assign n2709 = ( ~n2673 & n2675 ) | ( ~n2673 & n2677 ) | ( n2675 & n2677 ) ;
  assign n2710 = ( n2673 & ~n2678 ) | ( n2673 & n2709 ) | ( ~n2678 & n2709 ) ;
  assign n2711 = ( ~n2697 & n2699 ) | ( ~n2697 & n2701 ) | ( n2699 & n2701 ) ;
  assign n2712 = ( n2697 & ~n2702 ) | ( n2697 & n2711 ) | ( ~n2702 & n2711 ) ;
  assign n2713 = n2710 & n2712 ;
  assign n2714 = ( ~n2678 & n2680 ) | ( ~n2678 & n2682 ) | ( n2680 & n2682 ) ;
  assign n2715 = ( n2678 & ~n2683 ) | ( n2678 & n2714 ) | ( ~n2683 & n2714 ) ;
  assign n2716 = ( ~n2702 & n2704 ) | ( ~n2702 & n2706 ) | ( n2704 & n2706 ) ;
  assign n2717 = ( n2702 & ~n2707 ) | ( n2702 & n2716 ) | ( ~n2707 & n2716 ) ;
  assign n2718 = ( n2713 & n2715 ) | ( n2713 & n2717 ) | ( n2715 & n2717 ) ;
  assign n2719 = ( n2668 & n2671 ) | ( n2668 & ~n2683 ) | ( n2671 & ~n2683 ) ;
  assign n2720 = ( n2683 & ~n2684 ) | ( n2683 & n2719 ) | ( ~n2684 & n2719 ) ;
  assign n2721 = ( n2692 & n2695 ) | ( n2692 & ~n2707 ) | ( n2695 & ~n2707 ) ;
  assign n2722 = ( n2707 & ~n2708 ) | ( n2707 & n2721 ) | ( ~n2708 & n2721 ) ;
  assign n2723 = ( n2718 & n2720 ) | ( n2718 & n2722 ) | ( n2720 & n2722 ) ;
  assign n2724 = ( n2684 & n2708 ) | ( n2684 & n2723 ) | ( n2708 & n2723 ) ;
  assign n2725 = n2646 | n2648 ;
  assign n2726 = ~n2649 & n2725 ;
  assign n2727 = n2710 | n2712 ;
  assign n2728 = ~n2713 & n2727 ;
  assign n2729 = n2726 & n2728 ;
  assign n2730 = ( ~n2649 & n2651 ) | ( ~n2649 & n2653 ) | ( n2651 & n2653 ) ;
  assign n2731 = ( n2649 & ~n2654 ) | ( n2649 & n2730 ) | ( ~n2654 & n2730 ) ;
  assign n2732 = ( ~n2713 & n2715 ) | ( ~n2713 & n2717 ) | ( n2715 & n2717 ) ;
  assign n2733 = ( n2713 & ~n2718 ) | ( n2713 & n2732 ) | ( ~n2718 & n2732 ) ;
  assign n2734 = ( n2729 & n2731 ) | ( n2729 & n2733 ) | ( n2731 & n2733 ) ;
  assign n2735 = ( ~n2654 & n2656 ) | ( ~n2654 & n2658 ) | ( n2656 & n2658 ) ;
  assign n2736 = ( n2654 & ~n2659 ) | ( n2654 & n2735 ) | ( ~n2659 & n2735 ) ;
  assign n2737 = ( ~n2718 & n2720 ) | ( ~n2718 & n2722 ) | ( n2720 & n2722 ) ;
  assign n2738 = ( n2718 & ~n2723 ) | ( n2718 & n2737 ) | ( ~n2723 & n2737 ) ;
  assign n2739 = ( n2734 & n2736 ) | ( n2734 & n2738 ) | ( n2736 & n2738 ) ;
  assign n2740 = ( n2620 & n2644 ) | ( n2620 & ~n2659 ) | ( n2644 & ~n2659 ) ;
  assign n2741 = ( n2659 & ~n2660 ) | ( n2659 & n2740 ) | ( ~n2660 & n2740 ) ;
  assign n2742 = ( n2684 & n2708 ) | ( n2684 & ~n2723 ) | ( n2708 & ~n2723 ) ;
  assign n2743 = ( n2723 & ~n2724 ) | ( n2723 & n2742 ) | ( ~n2724 & n2742 ) ;
  assign n2744 = ( n2739 & n2741 ) | ( n2739 & n2743 ) | ( n2741 & n2743 ) ;
  assign n2745 = ( n2660 & n2724 ) | ( n2660 & n2744 ) | ( n2724 & n2744 ) ;
  assign n2746 = ( ~n2500 & n2502 ) | ( ~n2500 & n2582 ) | ( n2502 & n2582 ) ;
  assign n2747 = ( n2500 & ~n2583 ) | ( n2500 & n2746 ) | ( ~n2583 & n2746 ) ;
  assign n2748 = n2726 | n2728 ;
  assign n2749 = ~n2729 & n2748 ;
  assign n2750 = n2747 & n2749 ;
  assign n2751 = ( ~n2578 & n2580 ) | ( ~n2578 & n2584 ) | ( n2580 & n2584 ) ;
  assign n2752 = ( n2578 & ~n2585 ) | ( n2578 & n2751 ) | ( ~n2585 & n2751 ) ;
  assign n2753 = ( n2729 & ~n2731 ) | ( n2729 & n2733 ) | ( ~n2731 & n2733 ) ;
  assign n2754 = ( n2731 & ~n2734 ) | ( n2731 & n2753 ) | ( ~n2734 & n2753 ) ;
  assign n2755 = ( n2750 & n2752 ) | ( n2750 & n2754 ) | ( n2752 & n2754 ) ;
  assign n2756 = ( ~n2585 & n2587 ) | ( ~n2585 & n2589 ) | ( n2587 & n2589 ) ;
  assign n2757 = ( n2585 & ~n2590 ) | ( n2585 & n2756 ) | ( ~n2590 & n2756 ) ;
  assign n2758 = ( n2734 & ~n2736 ) | ( n2734 & n2738 ) | ( ~n2736 & n2738 ) ;
  assign n2759 = ( n2736 & ~n2739 ) | ( n2736 & n2758 ) | ( ~n2739 & n2758 ) ;
  assign n2760 = ( n2755 & n2757 ) | ( n2755 & n2759 ) | ( n2757 & n2759 ) ;
  assign n2761 = ( ~n2739 & n2741 ) | ( ~n2739 & n2743 ) | ( n2741 & n2743 ) ;
  assign n2762 = ( n2739 & ~n2744 ) | ( n2739 & n2761 ) | ( ~n2744 & n2761 ) ;
  assign n2763 = ( ~n2590 & n2592 ) | ( ~n2590 & n2594 ) | ( n2592 & n2594 ) ;
  assign n2764 = ( n2590 & ~n2595 ) | ( n2590 & n2763 ) | ( ~n2595 & n2763 ) ;
  assign n2765 = ( n2760 & n2762 ) | ( n2760 & n2764 ) | ( n2762 & n2764 ) ;
  assign n2766 = ( n2512 & n2576 ) | ( n2512 & ~n2595 ) | ( n2576 & ~n2595 ) ;
  assign n2767 = ( n2595 & ~n2596 ) | ( n2595 & n2766 ) | ( ~n2596 & n2766 ) ;
  assign n2768 = ( n2660 & n2724 ) | ( n2660 & ~n2744 ) | ( n2724 & ~n2744 ) ;
  assign n2769 = ( n2744 & ~n2745 ) | ( n2744 & n2768 ) | ( ~n2745 & n2768 ) ;
  assign n2770 = ( n2765 & n2767 ) | ( n2765 & n2769 ) | ( n2767 & n2769 ) ;
  assign n2771 = ( n2596 & n2745 ) | ( n2596 & n2770 ) | ( n2745 & n2770 ) ;
  assign n2772 = ( x214 & x215 ) | ( x214 & x216 ) | ( x215 & x216 ) ;
  assign n2773 = ( x211 & x212 ) | ( x211 & x213 ) | ( x212 & x213 ) ;
  assign n2774 = ( ~x214 & x215 ) | ( ~x214 & x216 ) | ( x215 & x216 ) ;
  assign n2775 = ( x214 & ~n2772 ) | ( x214 & n2774 ) | ( ~n2772 & n2774 ) ;
  assign n2776 = ( ~x211 & x212 ) | ( ~x211 & x213 ) | ( x212 & x213 ) ;
  assign n2777 = ( x211 & ~n2773 ) | ( x211 & n2776 ) | ( ~n2773 & n2776 ) ;
  assign n2778 = n2775 & n2777 ;
  assign n2779 = ( n2772 & n2773 ) | ( n2772 & n2778 ) | ( n2773 & n2778 ) ;
  assign n2780 = ( x217 & x218 ) | ( x217 & x219 ) | ( x218 & x219 ) ;
  assign n2781 = ( x220 & x221 ) | ( x220 & x222 ) | ( x221 & x222 ) ;
  assign n2782 = n2780 & n2781 ;
  assign n2783 = n2775 | n2777 ;
  assign n2784 = ~n2778 & n2783 ;
  assign n2785 = ( ~x217 & x218 ) | ( ~x217 & x219 ) | ( x218 & x219 ) ;
  assign n2786 = ( x217 & ~n2780 ) | ( x217 & n2785 ) | ( ~n2780 & n2785 ) ;
  assign n2787 = ( ~x220 & x221 ) | ( ~x220 & x222 ) | ( x221 & x222 ) ;
  assign n2788 = ( x220 & ~n2781 ) | ( x220 & n2787 ) | ( ~n2781 & n2787 ) ;
  assign n2789 = ( n2784 & n2786 ) | ( n2784 & n2788 ) | ( n2786 & n2788 ) ;
  assign n2790 = ( ~n2772 & n2773 ) | ( ~n2772 & n2778 ) | ( n2773 & n2778 ) ;
  assign n2791 = ( n2772 & ~n2779 ) | ( n2772 & n2790 ) | ( ~n2779 & n2790 ) ;
  assign n2792 = n2780 | n2781 ;
  assign n2793 = ~n2782 & n2792 ;
  assign n2794 = ( n2789 & n2791 ) | ( n2789 & n2793 ) | ( n2791 & n2793 ) ;
  assign n2795 = ( n2779 & n2782 ) | ( n2779 & n2794 ) | ( n2782 & n2794 ) ;
  assign n2796 = ( ~x199 & x200 ) | ( ~x199 & x201 ) | ( x200 & x201 ) ;
  assign n2797 = ( x199 & x200 ) | ( x199 & x201 ) | ( x200 & x201 ) ;
  assign n2798 = ( x199 & n2796 ) | ( x199 & ~n2797 ) | ( n2796 & ~n2797 ) ;
  assign n2799 = ( ~x202 & x203 ) | ( ~x202 & x204 ) | ( x203 & x204 ) ;
  assign n2800 = ( x202 & x203 ) | ( x202 & x204 ) | ( x203 & x204 ) ;
  assign n2801 = ( x202 & n2799 ) | ( x202 & ~n2800 ) | ( n2799 & ~n2800 ) ;
  assign n2802 = n2798 | n2801 ;
  assign n2803 = n2798 & n2801 ;
  assign n2804 = n2802 & ~n2803 ;
  assign n2805 = ( ~x205 & x206 ) | ( ~x205 & x207 ) | ( x206 & x207 ) ;
  assign n2806 = ( x205 & x206 ) | ( x205 & x207 ) | ( x206 & x207 ) ;
  assign n2807 = ( x205 & n2805 ) | ( x205 & ~n2806 ) | ( n2805 & ~n2806 ) ;
  assign n2808 = ( ~x208 & x209 ) | ( ~x208 & x210 ) | ( x209 & x210 ) ;
  assign n2809 = ( x208 & x209 ) | ( x208 & x210 ) | ( x209 & x210 ) ;
  assign n2810 = ( x208 & n2808 ) | ( x208 & ~n2809 ) | ( n2808 & ~n2809 ) ;
  assign n2811 = ( n2804 & n2807 ) | ( n2804 & n2810 ) | ( n2807 & n2810 ) ;
  assign n2812 = ( ~n2804 & n2807 ) | ( ~n2804 & n2810 ) | ( n2807 & n2810 ) ;
  assign n2813 = ( n2804 & ~n2811 ) | ( n2804 & n2812 ) | ( ~n2811 & n2812 ) ;
  assign n2814 = ( ~n2784 & n2786 ) | ( ~n2784 & n2788 ) | ( n2786 & n2788 ) ;
  assign n2815 = ( n2784 & ~n2789 ) | ( n2784 & n2814 ) | ( ~n2789 & n2814 ) ;
  assign n2816 = n2813 & n2815 ;
  assign n2817 = ( ~n2797 & n2800 ) | ( ~n2797 & n2803 ) | ( n2800 & n2803 ) ;
  assign n2818 = ( n2797 & n2800 ) | ( n2797 & n2803 ) | ( n2800 & n2803 ) ;
  assign n2819 = ( n2797 & n2817 ) | ( n2797 & ~n2818 ) | ( n2817 & ~n2818 ) ;
  assign n2820 = n2806 | n2809 ;
  assign n2821 = ~n2806 & n2809 ;
  assign n2822 = ( ~n2809 & n2820 ) | ( ~n2809 & n2821 ) | ( n2820 & n2821 ) ;
  assign n2823 = ( ~n2811 & n2819 ) | ( ~n2811 & n2822 ) | ( n2819 & n2822 ) ;
  assign n2824 = ( n2811 & n2819 ) | ( n2811 & n2822 ) | ( n2819 & n2822 ) ;
  assign n2825 = ( n2811 & n2823 ) | ( n2811 & ~n2824 ) | ( n2823 & ~n2824 ) ;
  assign n2826 = ( ~n2789 & n2791 ) | ( ~n2789 & n2793 ) | ( n2791 & n2793 ) ;
  assign n2827 = ( n2789 & ~n2794 ) | ( n2789 & n2826 ) | ( ~n2794 & n2826 ) ;
  assign n2828 = ( n2816 & n2825 ) | ( n2816 & n2827 ) | ( n2825 & n2827 ) ;
  assign n2829 = ( n2779 & n2782 ) | ( n2779 & ~n2794 ) | ( n2782 & ~n2794 ) ;
  assign n2830 = ( n2794 & ~n2795 ) | ( n2794 & n2829 ) | ( ~n2795 & n2829 ) ;
  assign n2831 = ( n2811 & n2819 ) | ( n2811 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2832 = ( n2809 & n2811 ) | ( n2809 & n2821 ) | ( n2811 & n2821 ) ;
  assign n2833 = ( n2809 & ~n2819 ) | ( n2809 & n2821 ) | ( ~n2819 & n2821 ) ;
  assign n2834 = ( n2831 & ~n2832 ) | ( n2831 & n2833 ) | ( ~n2832 & n2833 ) ;
  assign n2835 = n2818 | n2834 ;
  assign n2836 = n2818 & n2834 ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2838 = ( n2828 & n2830 ) | ( n2828 & n2837 ) | ( n2830 & n2837 ) ;
  assign n2839 = n2811 & n2819 ;
  assign n2840 = ( n2818 & ~n2837 ) | ( n2818 & n2839 ) | ( ~n2837 & n2839 ) ;
  assign n2841 = ( n2795 & n2838 ) | ( n2795 & n2840 ) | ( n2838 & n2840 ) ;
  assign n2842 = ( x178 & x179 ) | ( x178 & x180 ) | ( x179 & x180 ) ;
  assign n2843 = ( x175 & x176 ) | ( x175 & x177 ) | ( x176 & x177 ) ;
  assign n2844 = ( ~x178 & x179 ) | ( ~x178 & x180 ) | ( x179 & x180 ) ;
  assign n2845 = ( x178 & ~n2842 ) | ( x178 & n2844 ) | ( ~n2842 & n2844 ) ;
  assign n2846 = ( ~x175 & x176 ) | ( ~x175 & x177 ) | ( x176 & x177 ) ;
  assign n2847 = ( x175 & ~n2843 ) | ( x175 & n2846 ) | ( ~n2843 & n2846 ) ;
  assign n2848 = n2845 & n2847 ;
  assign n2849 = ( n2842 & n2843 ) | ( n2842 & n2848 ) | ( n2843 & n2848 ) ;
  assign n2850 = ( x181 & x182 ) | ( x181 & x183 ) | ( x182 & x183 ) ;
  assign n2851 = ( x184 & x185 ) | ( x184 & x186 ) | ( x185 & x186 ) ;
  assign n2852 = n2850 & n2851 ;
  assign n2853 = n2845 | n2847 ;
  assign n2854 = ~n2848 & n2853 ;
  assign n2855 = ( ~x181 & x182 ) | ( ~x181 & x183 ) | ( x182 & x183 ) ;
  assign n2856 = ( x181 & ~n2850 ) | ( x181 & n2855 ) | ( ~n2850 & n2855 ) ;
  assign n2857 = ( ~x184 & x185 ) | ( ~x184 & x186 ) | ( x185 & x186 ) ;
  assign n2858 = ( x184 & ~n2851 ) | ( x184 & n2857 ) | ( ~n2851 & n2857 ) ;
  assign n2859 = ( n2854 & n2856 ) | ( n2854 & n2858 ) | ( n2856 & n2858 ) ;
  assign n2860 = ( ~n2842 & n2843 ) | ( ~n2842 & n2848 ) | ( n2843 & n2848 ) ;
  assign n2861 = ( n2842 & ~n2849 ) | ( n2842 & n2860 ) | ( ~n2849 & n2860 ) ;
  assign n2862 = n2850 | n2851 ;
  assign n2863 = ~n2852 & n2862 ;
  assign n2864 = ( n2859 & n2861 ) | ( n2859 & n2863 ) | ( n2861 & n2863 ) ;
  assign n2865 = ( n2849 & n2852 ) | ( n2849 & n2864 ) | ( n2852 & n2864 ) ;
  assign n2866 = ( x187 & x188 ) | ( x187 & x189 ) | ( x188 & x189 ) ;
  assign n2867 = ( x190 & x191 ) | ( x190 & x192 ) | ( x191 & x192 ) ;
  assign n2868 = ( ~x187 & x188 ) | ( ~x187 & x189 ) | ( x188 & x189 ) ;
  assign n2869 = ( x187 & ~n2866 ) | ( x187 & n2868 ) | ( ~n2866 & n2868 ) ;
  assign n2870 = ( ~x190 & x191 ) | ( ~x190 & x192 ) | ( x191 & x192 ) ;
  assign n2871 = ( x190 & ~n2867 ) | ( x190 & n2870 ) | ( ~n2867 & n2870 ) ;
  assign n2872 = n2869 & n2871 ;
  assign n2873 = ( n2866 & n2867 ) | ( n2866 & n2872 ) | ( n2867 & n2872 ) ;
  assign n2874 = ( x193 & x194 ) | ( x193 & x195 ) | ( x194 & x195 ) ;
  assign n2875 = ( x196 & x197 ) | ( x196 & x198 ) | ( x197 & x198 ) ;
  assign n2876 = n2874 & n2875 ;
  assign n2877 = n2869 | n2871 ;
  assign n2878 = ~n2872 & n2877 ;
  assign n2879 = ( ~x193 & x194 ) | ( ~x193 & x195 ) | ( x194 & x195 ) ;
  assign n2880 = ( x193 & ~n2874 ) | ( x193 & n2879 ) | ( ~n2874 & n2879 ) ;
  assign n2881 = ( ~x196 & x197 ) | ( ~x196 & x198 ) | ( x197 & x198 ) ;
  assign n2882 = ( x196 & ~n2875 ) | ( x196 & n2881 ) | ( ~n2875 & n2881 ) ;
  assign n2883 = ( n2878 & n2880 ) | ( n2878 & n2882 ) | ( n2880 & n2882 ) ;
  assign n2884 = ( ~n2866 & n2867 ) | ( ~n2866 & n2872 ) | ( n2867 & n2872 ) ;
  assign n2885 = ( n2866 & ~n2873 ) | ( n2866 & n2884 ) | ( ~n2873 & n2884 ) ;
  assign n2886 = n2874 | n2875 ;
  assign n2887 = ~n2876 & n2886 ;
  assign n2888 = ( n2883 & n2885 ) | ( n2883 & n2887 ) | ( n2885 & n2887 ) ;
  assign n2889 = ( n2873 & n2876 ) | ( n2873 & n2888 ) | ( n2876 & n2888 ) ;
  assign n2890 = ( ~n2854 & n2856 ) | ( ~n2854 & n2858 ) | ( n2856 & n2858 ) ;
  assign n2891 = ( n2854 & ~n2859 ) | ( n2854 & n2890 ) | ( ~n2859 & n2890 ) ;
  assign n2892 = ( ~n2878 & n2880 ) | ( ~n2878 & n2882 ) | ( n2880 & n2882 ) ;
  assign n2893 = ( n2878 & ~n2883 ) | ( n2878 & n2892 ) | ( ~n2883 & n2892 ) ;
  assign n2894 = n2891 & n2893 ;
  assign n2895 = ( ~n2883 & n2885 ) | ( ~n2883 & n2887 ) | ( n2885 & n2887 ) ;
  assign n2896 = ( n2883 & ~n2888 ) | ( n2883 & n2895 ) | ( ~n2888 & n2895 ) ;
  assign n2897 = ( ~n2859 & n2861 ) | ( ~n2859 & n2863 ) | ( n2861 & n2863 ) ;
  assign n2898 = ( n2859 & ~n2864 ) | ( n2859 & n2897 ) | ( ~n2864 & n2897 ) ;
  assign n2899 = ( n2894 & n2896 ) | ( n2894 & n2898 ) | ( n2896 & n2898 ) ;
  assign n2900 = ( n2849 & n2852 ) | ( n2849 & ~n2864 ) | ( n2852 & ~n2864 ) ;
  assign n2901 = ( n2864 & ~n2865 ) | ( n2864 & n2900 ) | ( ~n2865 & n2900 ) ;
  assign n2902 = ( n2873 & n2876 ) | ( n2873 & ~n2888 ) | ( n2876 & ~n2888 ) ;
  assign n2903 = ( n2888 & ~n2889 ) | ( n2888 & n2902 ) | ( ~n2889 & n2902 ) ;
  assign n2904 = ( n2899 & n2901 ) | ( n2899 & n2903 ) | ( n2901 & n2903 ) ;
  assign n2905 = ( n2865 & n2889 ) | ( n2865 & n2904 ) | ( n2889 & n2904 ) ;
  assign n2906 = n2813 | n2815 ;
  assign n2907 = ~n2816 & n2906 ;
  assign n2908 = n2891 | n2893 ;
  assign n2909 = ~n2894 & n2908 ;
  assign n2910 = n2907 & n2909 ;
  assign n2911 = ( ~n2816 & n2825 ) | ( ~n2816 & n2827 ) | ( n2825 & n2827 ) ;
  assign n2912 = ( n2816 & ~n2828 ) | ( n2816 & n2911 ) | ( ~n2828 & n2911 ) ;
  assign n2913 = ( ~n2894 & n2896 ) | ( ~n2894 & n2898 ) | ( n2896 & n2898 ) ;
  assign n2914 = ( n2894 & ~n2899 ) | ( n2894 & n2913 ) | ( ~n2899 & n2913 ) ;
  assign n2915 = ( n2910 & n2912 ) | ( n2910 & n2914 ) | ( n2912 & n2914 ) ;
  assign n2916 = ( ~n2828 & n2830 ) | ( ~n2828 & n2837 ) | ( n2830 & n2837 ) ;
  assign n2917 = ( n2828 & ~n2838 ) | ( n2828 & n2916 ) | ( ~n2838 & n2916 ) ;
  assign n2918 = ( ~n2899 & n2901 ) | ( ~n2899 & n2903 ) | ( n2901 & n2903 ) ;
  assign n2919 = ( n2899 & ~n2904 ) | ( n2899 & n2918 ) | ( ~n2904 & n2918 ) ;
  assign n2920 = ( n2915 & n2917 ) | ( n2915 & n2919 ) | ( n2917 & n2919 ) ;
  assign n2921 = ( ~n2795 & n2838 ) | ( ~n2795 & n2840 ) | ( n2838 & n2840 ) ;
  assign n2922 = ( n2795 & ~n2841 ) | ( n2795 & n2921 ) | ( ~n2841 & n2921 ) ;
  assign n2923 = ( n2865 & n2889 ) | ( n2865 & ~n2904 ) | ( n2889 & ~n2904 ) ;
  assign n2924 = ( n2904 & ~n2905 ) | ( n2904 & n2923 ) | ( ~n2905 & n2923 ) ;
  assign n2925 = ( n2920 & n2922 ) | ( n2920 & n2924 ) | ( n2922 & n2924 ) ;
  assign n2926 = ( n2841 & n2905 ) | ( n2841 & n2925 ) | ( n2905 & n2925 ) ;
  assign n2927 = ( x235 & x236 ) | ( x235 & x237 ) | ( x236 & x237 ) ;
  assign n2928 = ( x238 & x239 ) | ( x238 & x240 ) | ( x239 & x240 ) ;
  assign n2929 = ( ~x235 & x236 ) | ( ~x235 & x237 ) | ( x236 & x237 ) ;
  assign n2930 = ( x235 & ~n2927 ) | ( x235 & n2929 ) | ( ~n2927 & n2929 ) ;
  assign n2931 = ( ~x238 & x239 ) | ( ~x238 & x240 ) | ( x239 & x240 ) ;
  assign n2932 = ( x238 & ~n2928 ) | ( x238 & n2931 ) | ( ~n2928 & n2931 ) ;
  assign n2933 = n2930 & n2932 ;
  assign n2934 = ( n2927 & n2928 ) | ( n2927 & n2933 ) | ( n2928 & n2933 ) ;
  assign n2935 = ( x244 & x245 ) | ( x244 & x246 ) | ( x245 & x246 ) ;
  assign n2936 = ( x241 & x242 ) | ( x241 & x243 ) | ( x242 & x243 ) ;
  assign n2937 = n2935 & n2936 ;
  assign n2938 = n2930 | n2932 ;
  assign n2939 = ~n2933 & n2938 ;
  assign n2940 = ( ~x244 & x245 ) | ( ~x244 & x246 ) | ( x245 & x246 ) ;
  assign n2941 = ( x244 & ~n2935 ) | ( x244 & n2940 ) | ( ~n2935 & n2940 ) ;
  assign n2942 = ( ~x241 & x242 ) | ( ~x241 & x243 ) | ( x242 & x243 ) ;
  assign n2943 = ( x241 & ~n2936 ) | ( x241 & n2942 ) | ( ~n2936 & n2942 ) ;
  assign n2944 = ( n2939 & n2941 ) | ( n2939 & n2943 ) | ( n2941 & n2943 ) ;
  assign n2945 = ( ~n2927 & n2928 ) | ( ~n2927 & n2933 ) | ( n2928 & n2933 ) ;
  assign n2946 = ( n2927 & ~n2934 ) | ( n2927 & n2945 ) | ( ~n2934 & n2945 ) ;
  assign n2947 = n2935 | n2936 ;
  assign n2948 = ~n2937 & n2947 ;
  assign n2949 = ( n2944 & n2946 ) | ( n2944 & n2948 ) | ( n2946 & n2948 ) ;
  assign n2950 = ( n2934 & n2937 ) | ( n2934 & n2949 ) | ( n2937 & n2949 ) ;
  assign n2951 = ( x226 & x227 ) | ( x226 & x228 ) | ( x227 & x228 ) ;
  assign n2952 = ( x223 & x224 ) | ( x223 & x225 ) | ( x224 & x225 ) ;
  assign n2953 = ( ~x226 & x227 ) | ( ~x226 & x228 ) | ( x227 & x228 ) ;
  assign n2954 = ( x226 & ~n2951 ) | ( x226 & n2953 ) | ( ~n2951 & n2953 ) ;
  assign n2955 = ( ~x223 & x224 ) | ( ~x223 & x225 ) | ( x224 & x225 ) ;
  assign n2956 = ( x223 & ~n2952 ) | ( x223 & n2955 ) | ( ~n2952 & n2955 ) ;
  assign n2957 = n2954 & n2956 ;
  assign n2958 = ( n2951 & n2952 ) | ( n2951 & n2957 ) | ( n2952 & n2957 ) ;
  assign n2959 = ( x229 & x230 ) | ( x229 & x231 ) | ( x230 & x231 ) ;
  assign n2960 = ( x232 & x233 ) | ( x232 & x234 ) | ( x233 & x234 ) ;
  assign n2961 = n2959 & n2960 ;
  assign n2962 = n2954 | n2956 ;
  assign n2963 = ~n2957 & n2962 ;
  assign n2964 = ( ~x229 & x230 ) | ( ~x229 & x231 ) | ( x230 & x231 ) ;
  assign n2965 = ( x229 & ~n2959 ) | ( x229 & n2964 ) | ( ~n2959 & n2964 ) ;
  assign n2966 = ( ~x232 & x233 ) | ( ~x232 & x234 ) | ( x233 & x234 ) ;
  assign n2967 = ( x232 & ~n2960 ) | ( x232 & n2966 ) | ( ~n2960 & n2966 ) ;
  assign n2968 = ( n2963 & n2965 ) | ( n2963 & n2967 ) | ( n2965 & n2967 ) ;
  assign n2969 = ( ~n2951 & n2952 ) | ( ~n2951 & n2957 ) | ( n2952 & n2957 ) ;
  assign n2970 = ( n2951 & ~n2958 ) | ( n2951 & n2969 ) | ( ~n2958 & n2969 ) ;
  assign n2971 = n2959 | n2960 ;
  assign n2972 = ~n2961 & n2971 ;
  assign n2973 = ( n2968 & n2970 ) | ( n2968 & n2972 ) | ( n2970 & n2972 ) ;
  assign n2974 = ( n2958 & n2961 ) | ( n2958 & n2973 ) | ( n2961 & n2973 ) ;
  assign n2975 = ( ~n2939 & n2941 ) | ( ~n2939 & n2943 ) | ( n2941 & n2943 ) ;
  assign n2976 = ( n2939 & ~n2944 ) | ( n2939 & n2975 ) | ( ~n2944 & n2975 ) ;
  assign n2977 = ( ~n2963 & n2965 ) | ( ~n2963 & n2967 ) | ( n2965 & n2967 ) ;
  assign n2978 = ( n2963 & ~n2968 ) | ( n2963 & n2977 ) | ( ~n2968 & n2977 ) ;
  assign n2979 = n2976 & n2978 ;
  assign n2980 = ( ~n2944 & n2946 ) | ( ~n2944 & n2948 ) | ( n2946 & n2948 ) ;
  assign n2981 = ( n2944 & ~n2949 ) | ( n2944 & n2980 ) | ( ~n2949 & n2980 ) ;
  assign n2982 = ( ~n2968 & n2970 ) | ( ~n2968 & n2972 ) | ( n2970 & n2972 ) ;
  assign n2983 = ( n2968 & ~n2973 ) | ( n2968 & n2982 ) | ( ~n2973 & n2982 ) ;
  assign n2984 = ( n2979 & n2981 ) | ( n2979 & n2983 ) | ( n2981 & n2983 ) ;
  assign n2985 = ( n2934 & n2937 ) | ( n2934 & ~n2949 ) | ( n2937 & ~n2949 ) ;
  assign n2986 = ( n2949 & ~n2950 ) | ( n2949 & n2985 ) | ( ~n2950 & n2985 ) ;
  assign n2987 = ( n2958 & n2961 ) | ( n2958 & ~n2973 ) | ( n2961 & ~n2973 ) ;
  assign n2988 = ( n2973 & ~n2974 ) | ( n2973 & n2987 ) | ( ~n2974 & n2987 ) ;
  assign n2989 = ( n2984 & n2986 ) | ( n2984 & n2988 ) | ( n2986 & n2988 ) ;
  assign n2990 = ( n2950 & n2974 ) | ( n2950 & n2989 ) | ( n2974 & n2989 ) ;
  assign n2991 = ( x265 & x266 ) | ( x265 & x267 ) | ( x266 & x267 ) ;
  assign n2992 = ( x268 & x269 ) | ( x268 & x270 ) | ( x269 & x270 ) ;
  assign n2993 = ( ~x265 & x266 ) | ( ~x265 & x267 ) | ( x266 & x267 ) ;
  assign n2994 = ( x265 & ~n2991 ) | ( x265 & n2993 ) | ( ~n2991 & n2993 ) ;
  assign n2995 = ( ~x268 & x269 ) | ( ~x268 & x270 ) | ( x269 & x270 ) ;
  assign n2996 = ( x268 & ~n2992 ) | ( x268 & n2995 ) | ( ~n2992 & n2995 ) ;
  assign n2997 = n2994 & n2996 ;
  assign n2998 = ( n2991 & n2992 ) | ( n2991 & n2997 ) | ( n2992 & n2997 ) ;
  assign n2999 = ( x262 & x263 ) | ( x262 & x264 ) | ( x263 & x264 ) ;
  assign n3000 = ( x259 & x260 ) | ( x259 & x261 ) | ( x260 & x261 ) ;
  assign n3001 = n2999 & n3000 ;
  assign n3002 = n2994 | n2996 ;
  assign n3003 = ~n2997 & n3002 ;
  assign n3004 = ( ~x262 & x263 ) | ( ~x262 & x264 ) | ( x263 & x264 ) ;
  assign n3005 = ( x262 & ~n2999 ) | ( x262 & n3004 ) | ( ~n2999 & n3004 ) ;
  assign n3006 = ( ~x259 & x260 ) | ( ~x259 & x261 ) | ( x260 & x261 ) ;
  assign n3007 = ( x259 & ~n3000 ) | ( x259 & n3006 ) | ( ~n3000 & n3006 ) ;
  assign n3008 = ( n3003 & n3005 ) | ( n3003 & n3007 ) | ( n3005 & n3007 ) ;
  assign n3009 = ( ~n2991 & n2992 ) | ( ~n2991 & n2997 ) | ( n2992 & n2997 ) ;
  assign n3010 = ( n2991 & ~n2998 ) | ( n2991 & n3009 ) | ( ~n2998 & n3009 ) ;
  assign n3011 = n2999 | n3000 ;
  assign n3012 = ~n3001 & n3011 ;
  assign n3013 = ( n3008 & n3010 ) | ( n3008 & n3012 ) | ( n3010 & n3012 ) ;
  assign n3014 = ( n2998 & n3001 ) | ( n2998 & n3013 ) | ( n3001 & n3013 ) ;
  assign n3015 = ( x250 & x251 ) | ( x250 & x252 ) | ( x251 & x252 ) ;
  assign n3016 = ( x247 & x248 ) | ( x247 & x249 ) | ( x248 & x249 ) ;
  assign n3017 = ( ~x250 & x251 ) | ( ~x250 & x252 ) | ( x251 & x252 ) ;
  assign n3018 = ( x250 & ~n3015 ) | ( x250 & n3017 ) | ( ~n3015 & n3017 ) ;
  assign n3019 = ( ~x247 & x248 ) | ( ~x247 & x249 ) | ( x248 & x249 ) ;
  assign n3020 = ( x247 & ~n3016 ) | ( x247 & n3019 ) | ( ~n3016 & n3019 ) ;
  assign n3021 = n3018 & n3020 ;
  assign n3022 = ( n3015 & n3016 ) | ( n3015 & n3021 ) | ( n3016 & n3021 ) ;
  assign n3023 = ( x253 & x254 ) | ( x253 & x255 ) | ( x254 & x255 ) ;
  assign n3024 = ( x256 & x257 ) | ( x256 & x258 ) | ( x257 & x258 ) ;
  assign n3025 = ( ~x253 & x254 ) | ( ~x253 & x255 ) | ( x254 & x255 ) ;
  assign n3026 = ( x253 & ~n3023 ) | ( x253 & n3025 ) | ( ~n3023 & n3025 ) ;
  assign n3027 = ( ~x256 & x257 ) | ( ~x256 & x258 ) | ( x257 & x258 ) ;
  assign n3028 = ( x256 & ~n3024 ) | ( x256 & n3027 ) | ( ~n3024 & n3027 ) ;
  assign n3029 = n3026 & n3028 ;
  assign n3030 = ( n3023 & n3024 ) | ( n3023 & n3029 ) | ( n3024 & n3029 ) ;
  assign n3031 = ( ~n3015 & n3016 ) | ( ~n3015 & n3021 ) | ( n3016 & n3021 ) ;
  assign n3032 = ( n3015 & ~n3022 ) | ( n3015 & n3031 ) | ( ~n3022 & n3031 ) ;
  assign n3033 = ( n3023 & n3024 ) | ( n3023 & ~n3029 ) | ( n3024 & ~n3029 ) ;
  assign n3034 = n3023 | n3024 ;
  assign n3035 = n3018 | n3020 ;
  assign n3036 = ~n3021 & n3035 ;
  assign n3037 = ( n3026 & n3028 ) | ( n3026 & n3036 ) | ( n3028 & n3036 ) ;
  assign n3038 = ( n3033 & ~n3034 ) | ( n3033 & n3037 ) | ( ~n3034 & n3037 ) ;
  assign n3039 = ~n3030 & n3033 ;
  assign n3040 = ( n3032 & n3038 ) | ( n3032 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3041 = ( n3022 & n3030 ) | ( n3022 & n3040 ) | ( n3030 & n3040 ) ;
  assign n3042 = ( ~n3003 & n3005 ) | ( ~n3003 & n3007 ) | ( n3005 & n3007 ) ;
  assign n3043 = ( n3003 & ~n3008 ) | ( n3003 & n3042 ) | ( ~n3008 & n3042 ) ;
  assign n3044 = ( n3026 & n3028 ) | ( n3026 & ~n3036 ) | ( n3028 & ~n3036 ) ;
  assign n3045 = ( n3036 & ~n3037 ) | ( n3036 & n3044 ) | ( ~n3037 & n3044 ) ;
  assign n3046 = n3043 & n3045 ;
  assign n3047 = ( ~n3008 & n3010 ) | ( ~n3008 & n3012 ) | ( n3010 & n3012 ) ;
  assign n3048 = ( n3008 & ~n3013 ) | ( n3008 & n3047 ) | ( ~n3013 & n3047 ) ;
  assign n3049 = ( ~n3032 & n3038 ) | ( ~n3032 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3050 = ( n3032 & ~n3040 ) | ( n3032 & n3049 ) | ( ~n3040 & n3049 ) ;
  assign n3051 = ( n3046 & n3048 ) | ( n3046 & n3050 ) | ( n3048 & n3050 ) ;
  assign n3052 = ( n2998 & n3001 ) | ( n2998 & ~n3013 ) | ( n3001 & ~n3013 ) ;
  assign n3053 = ( n3013 & ~n3014 ) | ( n3013 & n3052 ) | ( ~n3014 & n3052 ) ;
  assign n3054 = ( ~n3022 & n3030 ) | ( ~n3022 & n3040 ) | ( n3030 & n3040 ) ;
  assign n3055 = ( n3022 & ~n3041 ) | ( n3022 & n3054 ) | ( ~n3041 & n3054 ) ;
  assign n3056 = ( n3051 & n3053 ) | ( n3051 & n3055 ) | ( n3053 & n3055 ) ;
  assign n3057 = ( n3014 & n3041 ) | ( n3014 & n3056 ) | ( n3041 & n3056 ) ;
  assign n3058 = n3043 | n3045 ;
  assign n3059 = ~n3046 & n3058 ;
  assign n3060 = n2976 | n2978 ;
  assign n3061 = ~n2979 & n3060 ;
  assign n3062 = n3059 & n3061 ;
  assign n3063 = ( ~n2979 & n2981 ) | ( ~n2979 & n2983 ) | ( n2981 & n2983 ) ;
  assign n3064 = ( n2979 & ~n2984 ) | ( n2979 & n3063 ) | ( ~n2984 & n3063 ) ;
  assign n3065 = ( n3046 & ~n3048 ) | ( n3046 & n3050 ) | ( ~n3048 & n3050 ) ;
  assign n3066 = ( n3048 & ~n3051 ) | ( n3048 & n3065 ) | ( ~n3051 & n3065 ) ;
  assign n3067 = ( n3062 & n3064 ) | ( n3062 & n3066 ) | ( n3064 & n3066 ) ;
  assign n3068 = ( ~n2984 & n2986 ) | ( ~n2984 & n2988 ) | ( n2986 & n2988 ) ;
  assign n3069 = ( n2984 & ~n2989 ) | ( n2984 & n3068 ) | ( ~n2989 & n3068 ) ;
  assign n3070 = ( ~n3051 & n3053 ) | ( ~n3051 & n3055 ) | ( n3053 & n3055 ) ;
  assign n3071 = ( n3051 & ~n3056 ) | ( n3051 & n3070 ) | ( ~n3056 & n3070 ) ;
  assign n3072 = ( n3067 & n3069 ) | ( n3067 & n3071 ) | ( n3069 & n3071 ) ;
  assign n3073 = ( n2950 & n2974 ) | ( n2950 & ~n2989 ) | ( n2974 & ~n2989 ) ;
  assign n3074 = ( n2989 & ~n2990 ) | ( n2989 & n3073 ) | ( ~n2990 & n3073 ) ;
  assign n3075 = ( n3014 & n3041 ) | ( n3014 & ~n3056 ) | ( n3041 & ~n3056 ) ;
  assign n3076 = ( n3056 & ~n3057 ) | ( n3056 & n3075 ) | ( ~n3057 & n3075 ) ;
  assign n3077 = ( n3072 & n3074 ) | ( n3072 & n3076 ) | ( n3074 & n3076 ) ;
  assign n3078 = ( n2990 & n3057 ) | ( n2990 & n3077 ) | ( n3057 & n3077 ) ;
  assign n3079 = n2907 | n2909 ;
  assign n3080 = ~n2910 & n3079 ;
  assign n3081 = n3059 | n3061 ;
  assign n3082 = ~n3062 & n3081 ;
  assign n3083 = n3080 & n3082 ;
  assign n3084 = ( ~n2910 & n2912 ) | ( ~n2910 & n2914 ) | ( n2912 & n2914 ) ;
  assign n3085 = ( n2910 & ~n2915 ) | ( n2910 & n3084 ) | ( ~n2915 & n3084 ) ;
  assign n3086 = ( n3062 & ~n3064 ) | ( n3062 & n3066 ) | ( ~n3064 & n3066 ) ;
  assign n3087 = ( n3064 & ~n3067 ) | ( n3064 & n3086 ) | ( ~n3067 & n3086 ) ;
  assign n3088 = ( n3083 & n3085 ) | ( n3083 & n3087 ) | ( n3085 & n3087 ) ;
  assign n3089 = ( n2915 & ~n2917 ) | ( n2915 & n2919 ) | ( ~n2917 & n2919 ) ;
  assign n3090 = ( n2917 & ~n2920 ) | ( n2917 & n3089 ) | ( ~n2920 & n3089 ) ;
  assign n3091 = ( ~n3067 & n3069 ) | ( ~n3067 & n3071 ) | ( n3069 & n3071 ) ;
  assign n3092 = ( n3067 & ~n3072 ) | ( n3067 & n3091 ) | ( ~n3072 & n3091 ) ;
  assign n3093 = ( n3088 & n3090 ) | ( n3088 & n3092 ) | ( n3090 & n3092 ) ;
  assign n3094 = ( ~n3072 & n3074 ) | ( ~n3072 & n3076 ) | ( n3074 & n3076 ) ;
  assign n3095 = ( n3072 & ~n3077 ) | ( n3072 & n3094 ) | ( ~n3077 & n3094 ) ;
  assign n3096 = ( n2920 & ~n2922 ) | ( n2920 & n2924 ) | ( ~n2922 & n2924 ) ;
  assign n3097 = ( n2922 & ~n2925 ) | ( n2922 & n3096 ) | ( ~n2925 & n3096 ) ;
  assign n3098 = ( n3093 & n3095 ) | ( n3093 & n3097 ) | ( n3095 & n3097 ) ;
  assign n3099 = ( n2841 & n2905 ) | ( n2841 & ~n2925 ) | ( n2905 & ~n2925 ) ;
  assign n3100 = ( n2925 & ~n2926 ) | ( n2925 & n3099 ) | ( ~n2926 & n3099 ) ;
  assign n3101 = ( n2990 & n3057 ) | ( n2990 & ~n3077 ) | ( n3057 & ~n3077 ) ;
  assign n3102 = ( n3077 & ~n3078 ) | ( n3077 & n3101 ) | ( ~n3078 & n3101 ) ;
  assign n3103 = ( n3098 & n3100 ) | ( n3098 & n3102 ) | ( n3100 & n3102 ) ;
  assign n3104 = ( n2926 & n3078 ) | ( n2926 & n3103 ) | ( n3078 & n3103 ) ;
  assign n3105 = n2747 | n2749 ;
  assign n3106 = ~n2750 & n3105 ;
  assign n3107 = n3080 | n3082 ;
  assign n3108 = ~n3083 & n3107 ;
  assign n3109 = n3106 & n3108 ;
  assign n3110 = ( n2750 & ~n2752 ) | ( n2750 & n2754 ) | ( ~n2752 & n2754 ) ;
  assign n3111 = ( n2752 & ~n2755 ) | ( n2752 & n3110 ) | ( ~n2755 & n3110 ) ;
  assign n3112 = ( n3083 & ~n3085 ) | ( n3083 & n3087 ) | ( ~n3085 & n3087 ) ;
  assign n3113 = ( n3085 & ~n3088 ) | ( n3085 & n3112 ) | ( ~n3088 & n3112 ) ;
  assign n3114 = ( n3109 & n3111 ) | ( n3109 & n3113 ) | ( n3111 & n3113 ) ;
  assign n3115 = ( ~n2755 & n2757 ) | ( ~n2755 & n2759 ) | ( n2757 & n2759 ) ;
  assign n3116 = ( n2755 & ~n2760 ) | ( n2755 & n3115 ) | ( ~n2760 & n3115 ) ;
  assign n3117 = ( n3088 & ~n3090 ) | ( n3088 & n3092 ) | ( ~n3090 & n3092 ) ;
  assign n3118 = ( n3090 & ~n3093 ) | ( n3090 & n3117 ) | ( ~n3093 & n3117 ) ;
  assign n3119 = ( n3114 & n3116 ) | ( n3114 & n3118 ) | ( n3116 & n3118 ) ;
  assign n3120 = ( ~n2760 & n2762 ) | ( ~n2760 & n2764 ) | ( n2762 & n2764 ) ;
  assign n3121 = ( n2760 & ~n2765 ) | ( n2760 & n3120 ) | ( ~n2765 & n3120 ) ;
  assign n3122 = ( ~n3093 & n3095 ) | ( ~n3093 & n3097 ) | ( n3095 & n3097 ) ;
  assign n3123 = ( n3093 & ~n3098 ) | ( n3093 & n3122 ) | ( ~n3098 & n3122 ) ;
  assign n3124 = ( n3119 & n3121 ) | ( n3119 & n3123 ) | ( n3121 & n3123 ) ;
  assign n3125 = ( ~n2765 & n2767 ) | ( ~n2765 & n2769 ) | ( n2767 & n2769 ) ;
  assign n3126 = ( n2765 & ~n2770 ) | ( n2765 & n3125 ) | ( ~n2770 & n3125 ) ;
  assign n3127 = ( ~n3098 & n3100 ) | ( ~n3098 & n3102 ) | ( n3100 & n3102 ) ;
  assign n3128 = ( n3098 & ~n3103 ) | ( n3098 & n3127 ) | ( ~n3103 & n3127 ) ;
  assign n3129 = ( n3124 & n3126 ) | ( n3124 & n3128 ) | ( n3126 & n3128 ) ;
  assign n3130 = ( n2596 & n2745 ) | ( n2596 & ~n2770 ) | ( n2745 & ~n2770 ) ;
  assign n3131 = ( n2770 & ~n2771 ) | ( n2770 & n3130 ) | ( ~n2771 & n3130 ) ;
  assign n3132 = ( n2926 & n3078 ) | ( n2926 & ~n3103 ) | ( n3078 & ~n3103 ) ;
  assign n3133 = ( n3103 & ~n3104 ) | ( n3103 & n3132 ) | ( ~n3104 & n3132 ) ;
  assign n3134 = ( n3129 & n3131 ) | ( n3129 & n3133 ) | ( n3131 & n3133 ) ;
  assign n3135 = ( n2771 & n3104 ) | ( n2771 & n3134 ) | ( n3104 & n3134 ) ;
  assign n3136 = ( x364 & x365 ) | ( x364 & x366 ) | ( x365 & x366 ) ;
  assign n3137 = ( x361 & x362 ) | ( x361 & x363 ) | ( x362 & x363 ) ;
  assign n3138 = ( ~x364 & x365 ) | ( ~x364 & x366 ) | ( x365 & x366 ) ;
  assign n3139 = ( x364 & ~n3136 ) | ( x364 & n3138 ) | ( ~n3136 & n3138 ) ;
  assign n3140 = ( ~x361 & x362 ) | ( ~x361 & x363 ) | ( x362 & x363 ) ;
  assign n3141 = ( x361 & ~n3137 ) | ( x361 & n3140 ) | ( ~n3137 & n3140 ) ;
  assign n3142 = n3139 & n3141 ;
  assign n3143 = ( n3136 & n3137 ) | ( n3136 & n3142 ) | ( n3137 & n3142 ) ;
  assign n3144 = ( x355 & x356 ) | ( x355 & x357 ) | ( x356 & x357 ) ;
  assign n3145 = ( x358 & x359 ) | ( x358 & x360 ) | ( x359 & x360 ) ;
  assign n3146 = n3144 & n3145 ;
  assign n3147 = n3139 | n3141 ;
  assign n3148 = ~n3142 & n3147 ;
  assign n3149 = ( ~x355 & x356 ) | ( ~x355 & x357 ) | ( x356 & x357 ) ;
  assign n3150 = ( x355 & ~n3144 ) | ( x355 & n3149 ) | ( ~n3144 & n3149 ) ;
  assign n3151 = ( ~x358 & x359 ) | ( ~x358 & x360 ) | ( x359 & x360 ) ;
  assign n3152 = ( x358 & ~n3145 ) | ( x358 & n3151 ) | ( ~n3145 & n3151 ) ;
  assign n3153 = ( n3148 & n3150 ) | ( n3148 & n3152 ) | ( n3150 & n3152 ) ;
  assign n3154 = ( ~n3136 & n3137 ) | ( ~n3136 & n3142 ) | ( n3137 & n3142 ) ;
  assign n3155 = ( n3136 & ~n3143 ) | ( n3136 & n3154 ) | ( ~n3143 & n3154 ) ;
  assign n3156 = n3144 | n3145 ;
  assign n3157 = ~n3146 & n3156 ;
  assign n3158 = ( n3153 & n3155 ) | ( n3153 & n3157 ) | ( n3155 & n3157 ) ;
  assign n3159 = ( n3143 & n3146 ) | ( n3143 & n3158 ) | ( n3146 & n3158 ) ;
  assign n3160 = ( ~x346 & x347 ) | ( ~x346 & x348 ) | ( x347 & x348 ) ;
  assign n3161 = ( x346 & x347 ) | ( x346 & x348 ) | ( x347 & x348 ) ;
  assign n3162 = ( x346 & n3160 ) | ( x346 & ~n3161 ) | ( n3160 & ~n3161 ) ;
  assign n3163 = ( ~x343 & x344 ) | ( ~x343 & x345 ) | ( x344 & x345 ) ;
  assign n3164 = ( x343 & x344 ) | ( x343 & x345 ) | ( x344 & x345 ) ;
  assign n3165 = ( x343 & n3163 ) | ( x343 & ~n3164 ) | ( n3163 & ~n3164 ) ;
  assign n3166 = n3162 | n3165 ;
  assign n3167 = n3162 & n3165 ;
  assign n3168 = n3166 & ~n3167 ;
  assign n3169 = ( ~x349 & x350 ) | ( ~x349 & x351 ) | ( x350 & x351 ) ;
  assign n3170 = ( x349 & x350 ) | ( x349 & x351 ) | ( x350 & x351 ) ;
  assign n3171 = ( x349 & n3169 ) | ( x349 & ~n3170 ) | ( n3169 & ~n3170 ) ;
  assign n3172 = ( ~x352 & x353 ) | ( ~x352 & x354 ) | ( x353 & x354 ) ;
  assign n3173 = ( x352 & x353 ) | ( x352 & x354 ) | ( x353 & x354 ) ;
  assign n3174 = ( x352 & n3172 ) | ( x352 & ~n3173 ) | ( n3172 & ~n3173 ) ;
  assign n3175 = ( ~n3168 & n3171 ) | ( ~n3168 & n3174 ) | ( n3171 & n3174 ) ;
  assign n3176 = ( n3168 & n3171 ) | ( n3168 & n3174 ) | ( n3171 & n3174 ) ;
  assign n3177 = ( n3168 & n3175 ) | ( n3168 & ~n3176 ) | ( n3175 & ~n3176 ) ;
  assign n3178 = ( ~n3148 & n3150 ) | ( ~n3148 & n3152 ) | ( n3150 & n3152 ) ;
  assign n3179 = ( n3148 & ~n3153 ) | ( n3148 & n3178 ) | ( ~n3153 & n3178 ) ;
  assign n3180 = n3177 & n3179 ;
  assign n3181 = ( ~n3161 & n3164 ) | ( ~n3161 & n3167 ) | ( n3164 & n3167 ) ;
  assign n3182 = ( n3161 & n3164 ) | ( n3161 & n3167 ) | ( n3164 & n3167 ) ;
  assign n3183 = ( n3161 & n3181 ) | ( n3161 & ~n3182 ) | ( n3181 & ~n3182 ) ;
  assign n3184 = n3176 & n3183 ;
  assign n3185 = n3176 | n3183 ;
  assign n3186 = ~n3184 & n3185 ;
  assign n3187 = ( n3170 & n3173 ) | ( n3170 & n3186 ) | ( n3173 & n3186 ) ;
  assign n3188 = ( ~n3170 & n3173 ) | ( ~n3170 & n3186 ) | ( n3173 & n3186 ) ;
  assign n3189 = ( n3170 & ~n3187 ) | ( n3170 & n3188 ) | ( ~n3187 & n3188 ) ;
  assign n3190 = ( ~n3153 & n3155 ) | ( ~n3153 & n3157 ) | ( n3155 & n3157 ) ;
  assign n3191 = ( n3153 & ~n3158 ) | ( n3153 & n3190 ) | ( ~n3158 & n3190 ) ;
  assign n3192 = ( n3180 & n3189 ) | ( n3180 & n3191 ) | ( n3189 & n3191 ) ;
  assign n3193 = ( n3173 & n3185 ) | ( n3173 & ~n3188 ) | ( n3185 & ~n3188 ) ;
  assign n3194 = n3170 & n3173 ;
  assign n3195 = n3184 & n3194 ;
  assign n3196 = ( n3182 & n3193 ) | ( n3182 & ~n3195 ) | ( n3193 & ~n3195 ) ;
  assign n3197 = n3182 & n3195 ;
  assign n3198 = n3182 & n3193 ;
  assign n3199 = ( n3196 & n3197 ) | ( n3196 & ~n3198 ) | ( n3197 & ~n3198 ) ;
  assign n3200 = ( n3143 & n3146 ) | ( n3143 & ~n3158 ) | ( n3146 & ~n3158 ) ;
  assign n3201 = ( n3158 & ~n3159 ) | ( n3158 & n3200 ) | ( ~n3159 & n3200 ) ;
  assign n3202 = ( n3192 & n3199 ) | ( n3192 & n3201 ) | ( n3199 & n3201 ) ;
  assign n3203 = ( n3182 & n3184 ) | ( n3182 & ~n3199 ) | ( n3184 & ~n3199 ) ;
  assign n3204 = ( n3159 & n3202 ) | ( n3159 & n3203 ) | ( n3202 & n3203 ) ;
  assign n3205 = ( x319 & x320 ) | ( x319 & x321 ) | ( x320 & x321 ) ;
  assign n3206 = ( x322 & x323 ) | ( x322 & x324 ) | ( x323 & x324 ) ;
  assign n3207 = ( ~x319 & x320 ) | ( ~x319 & x321 ) | ( x320 & x321 ) ;
  assign n3208 = ( x319 & ~n3205 ) | ( x319 & n3207 ) | ( ~n3205 & n3207 ) ;
  assign n3209 = ( ~x322 & x323 ) | ( ~x322 & x324 ) | ( x323 & x324 ) ;
  assign n3210 = ( x322 & ~n3206 ) | ( x322 & n3209 ) | ( ~n3206 & n3209 ) ;
  assign n3211 = n3208 & n3210 ;
  assign n3212 = ( n3205 & n3206 ) | ( n3205 & n3211 ) | ( n3206 & n3211 ) ;
  assign n3213 = n3208 | n3210 ;
  assign n3214 = ~n3211 & n3213 ;
  assign n3215 = ( ~x328 & x329 ) | ( ~x328 & x330 ) | ( x329 & x330 ) ;
  assign n3216 = ( x328 & x329 ) | ( x328 & x330 ) | ( x329 & x330 ) ;
  assign n3217 = ( x328 & n3215 ) | ( x328 & ~n3216 ) | ( n3215 & ~n3216 ) ;
  assign n3218 = ( ~x325 & x326 ) | ( ~x325 & x327 ) | ( x326 & x327 ) ;
  assign n3219 = ( x325 & x326 ) | ( x325 & x327 ) | ( x326 & x327 ) ;
  assign n3220 = ( x325 & n3218 ) | ( x325 & ~n3219 ) | ( n3218 & ~n3219 ) ;
  assign n3221 = ( n3214 & n3217 ) | ( n3214 & n3220 ) | ( n3217 & n3220 ) ;
  assign n3222 = ( ~n3205 & n3206 ) | ( ~n3205 & n3211 ) | ( n3206 & n3211 ) ;
  assign n3223 = ( n3205 & ~n3212 ) | ( n3205 & n3222 ) | ( ~n3212 & n3222 ) ;
  assign n3224 = n3216 & n3219 ;
  assign n3225 = n3216 | n3219 ;
  assign n3226 = ~n3224 & n3225 ;
  assign n3227 = ( n3221 & n3223 ) | ( n3221 & n3226 ) | ( n3223 & n3226 ) ;
  assign n3228 = ( ~n3214 & n3217 ) | ( ~n3214 & n3220 ) | ( n3217 & n3220 ) ;
  assign n3229 = ( n3221 & ~n3223 ) | ( n3221 & n3226 ) | ( ~n3223 & n3226 ) ;
  assign n3230 = n3228 & n3229 ;
  assign n3231 = n3227 & ~n3230 ;
  assign n3232 = n3217 & n3220 ;
  assign n3233 = ( n3216 & n3219 ) | ( n3216 & n3232 ) | ( n3219 & n3232 ) ;
  assign n3234 = ( n3212 & n3231 ) | ( n3212 & n3233 ) | ( n3231 & n3233 ) ;
  assign n3235 = ( x334 & x335 ) | ( x334 & x336 ) | ( x335 & x336 ) ;
  assign n3236 = ( x331 & x332 ) | ( x331 & x333 ) | ( x332 & x333 ) ;
  assign n3237 = ( ~x334 & x335 ) | ( ~x334 & x336 ) | ( x335 & x336 ) ;
  assign n3238 = ( x334 & ~n3235 ) | ( x334 & n3237 ) | ( ~n3235 & n3237 ) ;
  assign n3239 = ( ~x331 & x332 ) | ( ~x331 & x333 ) | ( x332 & x333 ) ;
  assign n3240 = ( x331 & ~n3236 ) | ( x331 & n3239 ) | ( ~n3236 & n3239 ) ;
  assign n3241 = n3238 & n3240 ;
  assign n3242 = ( n3235 & n3236 ) | ( n3235 & n3241 ) | ( n3236 & n3241 ) ;
  assign n3243 = ( x337 & x338 ) | ( x337 & x339 ) | ( x338 & x339 ) ;
  assign n3244 = ( x340 & x341 ) | ( x340 & x342 ) | ( x341 & x342 ) ;
  assign n3245 = n3243 & n3244 ;
  assign n3246 = n3238 | n3240 ;
  assign n3247 = ~n3241 & n3246 ;
  assign n3248 = ( ~x337 & x338 ) | ( ~x337 & x339 ) | ( x338 & x339 ) ;
  assign n3249 = ( x337 & ~n3243 ) | ( x337 & n3248 ) | ( ~n3243 & n3248 ) ;
  assign n3250 = ( ~x340 & x341 ) | ( ~x340 & x342 ) | ( x341 & x342 ) ;
  assign n3251 = ( x340 & ~n3244 ) | ( x340 & n3250 ) | ( ~n3244 & n3250 ) ;
  assign n3252 = ( n3247 & n3249 ) | ( n3247 & n3251 ) | ( n3249 & n3251 ) ;
  assign n3253 = ( ~n3235 & n3236 ) | ( ~n3235 & n3241 ) | ( n3236 & n3241 ) ;
  assign n3254 = ( n3235 & ~n3242 ) | ( n3235 & n3253 ) | ( ~n3242 & n3253 ) ;
  assign n3255 = n3243 | n3244 ;
  assign n3256 = ~n3245 & n3255 ;
  assign n3257 = ( n3252 & n3254 ) | ( n3252 & n3256 ) | ( n3254 & n3256 ) ;
  assign n3258 = ( n3242 & n3245 ) | ( n3242 & n3257 ) | ( n3245 & n3257 ) ;
  assign n3259 = ( ~n3247 & n3249 ) | ( ~n3247 & n3251 ) | ( n3249 & n3251 ) ;
  assign n3260 = ( n3247 & ~n3252 ) | ( n3247 & n3259 ) | ( ~n3252 & n3259 ) ;
  assign n3261 = ( n3214 & ~n3221 ) | ( n3214 & n3228 ) | ( ~n3221 & n3228 ) ;
  assign n3262 = n3260 & n3261 ;
  assign n3263 = ( ~n3252 & n3254 ) | ( ~n3252 & n3256 ) | ( n3254 & n3256 ) ;
  assign n3264 = ( n3252 & ~n3257 ) | ( n3252 & n3263 ) | ( ~n3257 & n3263 ) ;
  assign n3265 = ( n3223 & ~n3227 ) | ( n3223 & n3229 ) | ( ~n3227 & n3229 ) ;
  assign n3266 = ( n3262 & n3264 ) | ( n3262 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3267 = ( ~n3212 & n3231 ) | ( ~n3212 & n3233 ) | ( n3231 & n3233 ) ;
  assign n3268 = ( n3212 & ~n3234 ) | ( n3212 & n3267 ) | ( ~n3234 & n3267 ) ;
  assign n3269 = ( n3242 & n3245 ) | ( n3242 & ~n3257 ) | ( n3245 & ~n3257 ) ;
  assign n3270 = ( n3257 & ~n3258 ) | ( n3257 & n3269 ) | ( ~n3258 & n3269 ) ;
  assign n3271 = ( n3266 & n3268 ) | ( n3266 & n3270 ) | ( n3268 & n3270 ) ;
  assign n3272 = ( n3234 & n3258 ) | ( n3234 & n3271 ) | ( n3258 & n3271 ) ;
  assign n3273 = n3260 | n3261 ;
  assign n3274 = ~n3262 & n3273 ;
  assign n3275 = n3177 | n3179 ;
  assign n3276 = ~n3180 & n3275 ;
  assign n3277 = n3274 & n3276 ;
  assign n3278 = ( ~n3180 & n3189 ) | ( ~n3180 & n3191 ) | ( n3189 & n3191 ) ;
  assign n3279 = ( n3180 & ~n3192 ) | ( n3180 & n3278 ) | ( ~n3192 & n3278 ) ;
  assign n3280 = ( ~n3262 & n3264 ) | ( ~n3262 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3281 = ( n3262 & ~n3266 ) | ( n3262 & n3280 ) | ( ~n3266 & n3280 ) ;
  assign n3282 = ( n3277 & n3279 ) | ( n3277 & n3281 ) | ( n3279 & n3281 ) ;
  assign n3283 = ( ~n3192 & n3199 ) | ( ~n3192 & n3201 ) | ( n3199 & n3201 ) ;
  assign n3284 = ( n3192 & ~n3202 ) | ( n3192 & n3283 ) | ( ~n3202 & n3283 ) ;
  assign n3285 = ( n3266 & ~n3268 ) | ( n3266 & n3270 ) | ( ~n3268 & n3270 ) ;
  assign n3286 = ( n3268 & ~n3271 ) | ( n3268 & n3285 ) | ( ~n3271 & n3285 ) ;
  assign n3287 = ( n3282 & n3284 ) | ( n3282 & n3286 ) | ( n3284 & n3286 ) ;
  assign n3288 = ( n3159 & ~n3202 ) | ( n3159 & n3203 ) | ( ~n3202 & n3203 ) ;
  assign n3289 = ( n3202 & ~n3204 ) | ( n3202 & n3288 ) | ( ~n3204 & n3288 ) ;
  assign n3290 = ( n3234 & n3258 ) | ( n3234 & ~n3271 ) | ( n3258 & ~n3271 ) ;
  assign n3291 = ( n3271 & ~n3272 ) | ( n3271 & n3290 ) | ( ~n3272 & n3290 ) ;
  assign n3292 = ( n3287 & n3289 ) | ( n3287 & n3291 ) | ( n3289 & n3291 ) ;
  assign n3293 = ( n3204 & n3272 ) | ( n3204 & n3292 ) | ( n3272 & n3292 ) ;
  assign n3294 = ( x298 & x299 ) | ( x298 & x300 ) | ( x299 & x300 ) ;
  assign n3295 = ( x295 & x296 ) | ( x295 & x297 ) | ( x296 & x297 ) ;
  assign n3296 = ( ~x298 & x299 ) | ( ~x298 & x300 ) | ( x299 & x300 ) ;
  assign n3297 = ( x298 & ~n3294 ) | ( x298 & n3296 ) | ( ~n3294 & n3296 ) ;
  assign n3298 = ( ~x295 & x296 ) | ( ~x295 & x297 ) | ( x296 & x297 ) ;
  assign n3299 = ( x295 & ~n3295 ) | ( x295 & n3298 ) | ( ~n3295 & n3298 ) ;
  assign n3300 = n3297 & n3299 ;
  assign n3301 = ( n3294 & n3295 ) | ( n3294 & n3300 ) | ( n3295 & n3300 ) ;
  assign n3302 = ( x304 & x305 ) | ( x304 & x306 ) | ( x305 & x306 ) ;
  assign n3303 = ( x301 & x302 ) | ( x301 & x303 ) | ( x302 & x303 ) ;
  assign n3304 = n3302 & n3303 ;
  assign n3305 = n3297 | n3299 ;
  assign n3306 = ~n3300 & n3305 ;
  assign n3307 = ( ~x304 & x305 ) | ( ~x304 & x306 ) | ( x305 & x306 ) ;
  assign n3308 = ( x304 & ~n3302 ) | ( x304 & n3307 ) | ( ~n3302 & n3307 ) ;
  assign n3309 = ( ~x301 & x302 ) | ( ~x301 & x303 ) | ( x302 & x303 ) ;
  assign n3310 = ( x301 & ~n3303 ) | ( x301 & n3309 ) | ( ~n3303 & n3309 ) ;
  assign n3311 = ( n3306 & n3308 ) | ( n3306 & n3310 ) | ( n3308 & n3310 ) ;
  assign n3312 = ( ~n3294 & n3295 ) | ( ~n3294 & n3300 ) | ( n3295 & n3300 ) ;
  assign n3313 = ( n3294 & ~n3301 ) | ( n3294 & n3312 ) | ( ~n3301 & n3312 ) ;
  assign n3314 = n3302 | n3303 ;
  assign n3315 = ~n3304 & n3314 ;
  assign n3316 = ( n3311 & n3313 ) | ( n3311 & n3315 ) | ( n3313 & n3315 ) ;
  assign n3317 = ( n3301 & n3304 ) | ( n3301 & n3316 ) | ( n3304 & n3316 ) ;
  assign n3318 = ( x307 & x308 ) | ( x307 & x309 ) | ( x308 & x309 ) ;
  assign n3319 = ( x310 & x311 ) | ( x310 & x312 ) | ( x311 & x312 ) ;
  assign n3320 = ( ~x307 & x308 ) | ( ~x307 & x309 ) | ( x308 & x309 ) ;
  assign n3321 = ( x307 & ~n3318 ) | ( x307 & n3320 ) | ( ~n3318 & n3320 ) ;
  assign n3322 = ( ~x310 & x311 ) | ( ~x310 & x312 ) | ( x311 & x312 ) ;
  assign n3323 = ( x310 & ~n3319 ) | ( x310 & n3322 ) | ( ~n3319 & n3322 ) ;
  assign n3324 = n3321 & n3323 ;
  assign n3325 = ( n3318 & n3319 ) | ( n3318 & n3324 ) | ( n3319 & n3324 ) ;
  assign n3326 = ( x313 & x314 ) | ( x313 & x315 ) | ( x314 & x315 ) ;
  assign n3327 = ( x316 & x317 ) | ( x316 & x318 ) | ( x317 & x318 ) ;
  assign n3328 = n3326 & n3327 ;
  assign n3329 = n3321 | n3323 ;
  assign n3330 = ~n3324 & n3329 ;
  assign n3331 = ( ~x313 & x314 ) | ( ~x313 & x315 ) | ( x314 & x315 ) ;
  assign n3332 = ( x313 & ~n3326 ) | ( x313 & n3331 ) | ( ~n3326 & n3331 ) ;
  assign n3333 = ( ~x316 & x317 ) | ( ~x316 & x318 ) | ( x317 & x318 ) ;
  assign n3334 = ( x316 & ~n3327 ) | ( x316 & n3333 ) | ( ~n3327 & n3333 ) ;
  assign n3335 = ( n3330 & n3332 ) | ( n3330 & n3334 ) | ( n3332 & n3334 ) ;
  assign n3336 = ( ~n3318 & n3319 ) | ( ~n3318 & n3324 ) | ( n3319 & n3324 ) ;
  assign n3337 = ( n3318 & ~n3325 ) | ( n3318 & n3336 ) | ( ~n3325 & n3336 ) ;
  assign n3338 = n3326 | n3327 ;
  assign n3339 = ~n3328 & n3338 ;
  assign n3340 = ( n3335 & n3337 ) | ( n3335 & n3339 ) | ( n3337 & n3339 ) ;
  assign n3341 = ( n3325 & n3328 ) | ( n3325 & n3340 ) | ( n3328 & n3340 ) ;
  assign n3342 = ( ~n3330 & n3332 ) | ( ~n3330 & n3334 ) | ( n3332 & n3334 ) ;
  assign n3343 = ( n3330 & ~n3335 ) | ( n3330 & n3342 ) | ( ~n3335 & n3342 ) ;
  assign n3344 = ( ~n3306 & n3308 ) | ( ~n3306 & n3310 ) | ( n3308 & n3310 ) ;
  assign n3345 = ( n3306 & ~n3311 ) | ( n3306 & n3344 ) | ( ~n3311 & n3344 ) ;
  assign n3346 = n3343 & n3345 ;
  assign n3347 = ( ~n3335 & n3337 ) | ( ~n3335 & n3339 ) | ( n3337 & n3339 ) ;
  assign n3348 = ( n3335 & ~n3340 ) | ( n3335 & n3347 ) | ( ~n3340 & n3347 ) ;
  assign n3349 = ( ~n3311 & n3313 ) | ( ~n3311 & n3315 ) | ( n3313 & n3315 ) ;
  assign n3350 = ( n3311 & ~n3316 ) | ( n3311 & n3349 ) | ( ~n3316 & n3349 ) ;
  assign n3351 = ( n3346 & n3348 ) | ( n3346 & n3350 ) | ( n3348 & n3350 ) ;
  assign n3352 = ( n3301 & n3304 ) | ( n3301 & ~n3316 ) | ( n3304 & ~n3316 ) ;
  assign n3353 = ( n3316 & ~n3317 ) | ( n3316 & n3352 ) | ( ~n3317 & n3352 ) ;
  assign n3354 = ( n3325 & n3328 ) | ( n3325 & ~n3340 ) | ( n3328 & ~n3340 ) ;
  assign n3355 = ( n3340 & ~n3341 ) | ( n3340 & n3354 ) | ( ~n3341 & n3354 ) ;
  assign n3356 = ( n3351 & n3353 ) | ( n3351 & n3355 ) | ( n3353 & n3355 ) ;
  assign n3357 = ( n3317 & n3341 ) | ( n3317 & n3356 ) | ( n3341 & n3356 ) ;
  assign n3358 = ( x286 & x287 ) | ( x286 & x288 ) | ( x287 & x288 ) ;
  assign n3359 = ( x283 & x284 ) | ( x283 & x285 ) | ( x284 & x285 ) ;
  assign n3360 = ( ~x286 & x287 ) | ( ~x286 & x288 ) | ( x287 & x288 ) ;
  assign n3361 = ( x286 & ~n3358 ) | ( x286 & n3360 ) | ( ~n3358 & n3360 ) ;
  assign n3362 = ( ~x283 & x284 ) | ( ~x283 & x285 ) | ( x284 & x285 ) ;
  assign n3363 = ( x283 & ~n3359 ) | ( x283 & n3362 ) | ( ~n3359 & n3362 ) ;
  assign n3364 = n3361 & n3363 ;
  assign n3365 = ( n3358 & n3359 ) | ( n3358 & n3364 ) | ( n3359 & n3364 ) ;
  assign n3366 = ( x292 & x293 ) | ( x292 & x294 ) | ( x293 & x294 ) ;
  assign n3367 = ( x289 & x290 ) | ( x289 & x291 ) | ( x290 & x291 ) ;
  assign n3368 = n3366 & n3367 ;
  assign n3369 = n3361 | n3363 ;
  assign n3370 = ~n3364 & n3369 ;
  assign n3371 = ( ~x292 & x293 ) | ( ~x292 & x294 ) | ( x293 & x294 ) ;
  assign n3372 = ( x292 & ~n3366 ) | ( x292 & n3371 ) | ( ~n3366 & n3371 ) ;
  assign n3373 = ( ~x289 & x290 ) | ( ~x289 & x291 ) | ( x290 & x291 ) ;
  assign n3374 = ( x289 & ~n3367 ) | ( x289 & n3373 ) | ( ~n3367 & n3373 ) ;
  assign n3375 = ( n3370 & n3372 ) | ( n3370 & n3374 ) | ( n3372 & n3374 ) ;
  assign n3376 = ( ~n3358 & n3359 ) | ( ~n3358 & n3364 ) | ( n3359 & n3364 ) ;
  assign n3377 = ( n3358 & ~n3365 ) | ( n3358 & n3376 ) | ( ~n3365 & n3376 ) ;
  assign n3378 = n3366 | n3367 ;
  assign n3379 = ~n3368 & n3378 ;
  assign n3380 = ( n3375 & n3377 ) | ( n3375 & n3379 ) | ( n3377 & n3379 ) ;
  assign n3381 = ( n3365 & n3368 ) | ( n3365 & n3380 ) | ( n3368 & n3380 ) ;
  assign n3382 = ( x271 & x272 ) | ( x271 & x273 ) | ( x272 & x273 ) ;
  assign n3383 = ( x274 & x275 ) | ( x274 & x276 ) | ( x275 & x276 ) ;
  assign n3384 = ( ~x271 & x272 ) | ( ~x271 & x273 ) | ( x272 & x273 ) ;
  assign n3385 = ( x271 & ~n3382 ) | ( x271 & n3384 ) | ( ~n3382 & n3384 ) ;
  assign n3386 = ( ~x274 & x275 ) | ( ~x274 & x276 ) | ( x275 & x276 ) ;
  assign n3387 = ( x274 & ~n3383 ) | ( x274 & n3386 ) | ( ~n3383 & n3386 ) ;
  assign n3388 = n3385 & n3387 ;
  assign n3389 = ( n3382 & n3383 ) | ( n3382 & n3388 ) | ( n3383 & n3388 ) ;
  assign n3390 = ( x280 & x281 ) | ( x280 & x282 ) | ( x281 & x282 ) ;
  assign n3391 = ( x277 & x278 ) | ( x277 & x279 ) | ( x278 & x279 ) ;
  assign n3392 = n3390 & n3391 ;
  assign n3393 = n3385 | n3387 ;
  assign n3394 = ~n3388 & n3393 ;
  assign n3395 = ( ~x280 & x281 ) | ( ~x280 & x282 ) | ( x281 & x282 ) ;
  assign n3396 = ( x280 & ~n3390 ) | ( x280 & n3395 ) | ( ~n3390 & n3395 ) ;
  assign n3397 = ( ~x277 & x278 ) | ( ~x277 & x279 ) | ( x278 & x279 ) ;
  assign n3398 = ( x277 & ~n3391 ) | ( x277 & n3397 ) | ( ~n3391 & n3397 ) ;
  assign n3399 = ( n3394 & n3396 ) | ( n3394 & n3398 ) | ( n3396 & n3398 ) ;
  assign n3400 = ( ~n3382 & n3383 ) | ( ~n3382 & n3388 ) | ( n3383 & n3388 ) ;
  assign n3401 = ( n3382 & ~n3389 ) | ( n3382 & n3400 ) | ( ~n3389 & n3400 ) ;
  assign n3402 = n3390 | n3391 ;
  assign n3403 = ~n3392 & n3402 ;
  assign n3404 = ( n3399 & n3401 ) | ( n3399 & n3403 ) | ( n3401 & n3403 ) ;
  assign n3405 = ( n3389 & n3392 ) | ( n3389 & n3404 ) | ( n3392 & n3404 ) ;
  assign n3406 = ( ~n3394 & n3396 ) | ( ~n3394 & n3398 ) | ( n3396 & n3398 ) ;
  assign n3407 = ( n3394 & ~n3399 ) | ( n3394 & n3406 ) | ( ~n3399 & n3406 ) ;
  assign n3408 = ( ~n3370 & n3372 ) | ( ~n3370 & n3374 ) | ( n3372 & n3374 ) ;
  assign n3409 = ( n3370 & ~n3375 ) | ( n3370 & n3408 ) | ( ~n3375 & n3408 ) ;
  assign n3410 = n3407 & n3409 ;
  assign n3411 = ( ~n3399 & n3401 ) | ( ~n3399 & n3403 ) | ( n3401 & n3403 ) ;
  assign n3412 = ( n3399 & ~n3404 ) | ( n3399 & n3411 ) | ( ~n3404 & n3411 ) ;
  assign n3413 = ( ~n3375 & n3377 ) | ( ~n3375 & n3379 ) | ( n3377 & n3379 ) ;
  assign n3414 = ( n3375 & ~n3380 ) | ( n3375 & n3413 ) | ( ~n3380 & n3413 ) ;
  assign n3415 = ( n3410 & n3412 ) | ( n3410 & n3414 ) | ( n3412 & n3414 ) ;
  assign n3416 = ( n3365 & n3368 ) | ( n3365 & ~n3380 ) | ( n3368 & ~n3380 ) ;
  assign n3417 = ( n3380 & ~n3381 ) | ( n3380 & n3416 ) | ( ~n3381 & n3416 ) ;
  assign n3418 = ( n3389 & n3392 ) | ( n3389 & ~n3404 ) | ( n3392 & ~n3404 ) ;
  assign n3419 = ( n3404 & ~n3405 ) | ( n3404 & n3418 ) | ( ~n3405 & n3418 ) ;
  assign n3420 = ( n3415 & n3417 ) | ( n3415 & n3419 ) | ( n3417 & n3419 ) ;
  assign n3421 = ( n3381 & n3405 ) | ( n3381 & n3420 ) | ( n3405 & n3420 ) ;
  assign n3422 = n3407 | n3409 ;
  assign n3423 = ~n3410 & n3422 ;
  assign n3424 = n3343 | n3345 ;
  assign n3425 = ~n3346 & n3424 ;
  assign n3426 = n3423 & n3425 ;
  assign n3427 = ( ~n3410 & n3412 ) | ( ~n3410 & n3414 ) | ( n3412 & n3414 ) ;
  assign n3428 = ( n3410 & ~n3415 ) | ( n3410 & n3427 ) | ( ~n3415 & n3427 ) ;
  assign n3429 = ( n3346 & ~n3348 ) | ( n3346 & n3350 ) | ( ~n3348 & n3350 ) ;
  assign n3430 = ( n3348 & ~n3351 ) | ( n3348 & n3429 ) | ( ~n3351 & n3429 ) ;
  assign n3431 = ( n3426 & n3428 ) | ( n3426 & n3430 ) | ( n3428 & n3430 ) ;
  assign n3432 = ( ~n3415 & n3417 ) | ( ~n3415 & n3419 ) | ( n3417 & n3419 ) ;
  assign n3433 = ( n3415 & ~n3420 ) | ( n3415 & n3432 ) | ( ~n3420 & n3432 ) ;
  assign n3434 = ( ~n3351 & n3353 ) | ( ~n3351 & n3355 ) | ( n3353 & n3355 ) ;
  assign n3435 = ( n3351 & ~n3356 ) | ( n3351 & n3434 ) | ( ~n3356 & n3434 ) ;
  assign n3436 = ( n3431 & n3433 ) | ( n3431 & n3435 ) | ( n3433 & n3435 ) ;
  assign n3437 = ( n3317 & n3341 ) | ( n3317 & ~n3356 ) | ( n3341 & ~n3356 ) ;
  assign n3438 = ( n3356 & ~n3357 ) | ( n3356 & n3437 ) | ( ~n3357 & n3437 ) ;
  assign n3439 = ( n3381 & n3405 ) | ( n3381 & ~n3420 ) | ( n3405 & ~n3420 ) ;
  assign n3440 = ( n3420 & ~n3421 ) | ( n3420 & n3439 ) | ( ~n3421 & n3439 ) ;
  assign n3441 = ( n3436 & n3438 ) | ( n3436 & n3440 ) | ( n3438 & n3440 ) ;
  assign n3442 = ( n3357 & n3421 ) | ( n3357 & n3441 ) | ( n3421 & n3441 ) ;
  assign n3443 = n3423 | n3425 ;
  assign n3444 = ~n3426 & n3443 ;
  assign n3445 = n3274 | n3276 ;
  assign n3446 = ~n3277 & n3445 ;
  assign n3447 = n3444 & n3446 ;
  assign n3448 = ( ~n3426 & n3428 ) | ( ~n3426 & n3430 ) | ( n3428 & n3430 ) ;
  assign n3449 = ( n3426 & ~n3431 ) | ( n3426 & n3448 ) | ( ~n3431 & n3448 ) ;
  assign n3450 = ( n3277 & ~n3279 ) | ( n3277 & n3281 ) | ( ~n3279 & n3281 ) ;
  assign n3451 = ( n3279 & ~n3282 ) | ( n3279 & n3450 ) | ( ~n3282 & n3450 ) ;
  assign n3452 = ( n3447 & n3449 ) | ( n3447 & n3451 ) | ( n3449 & n3451 ) ;
  assign n3453 = ( ~n3282 & n3284 ) | ( ~n3282 & n3286 ) | ( n3284 & n3286 ) ;
  assign n3454 = ( n3282 & ~n3287 ) | ( n3282 & n3453 ) | ( ~n3287 & n3453 ) ;
  assign n3455 = ( ~n3431 & n3433 ) | ( ~n3431 & n3435 ) | ( n3433 & n3435 ) ;
  assign n3456 = ( n3431 & ~n3436 ) | ( n3431 & n3455 ) | ( ~n3436 & n3455 ) ;
  assign n3457 = ( n3452 & n3454 ) | ( n3452 & n3456 ) | ( n3454 & n3456 ) ;
  assign n3458 = ( ~n3436 & n3438 ) | ( ~n3436 & n3440 ) | ( n3438 & n3440 ) ;
  assign n3459 = ( n3436 & ~n3441 ) | ( n3436 & n3458 ) | ( ~n3441 & n3458 ) ;
  assign n3460 = ( ~n3287 & n3289 ) | ( ~n3287 & n3291 ) | ( n3289 & n3291 ) ;
  assign n3461 = ( n3287 & ~n3292 ) | ( n3287 & n3460 ) | ( ~n3292 & n3460 ) ;
  assign n3462 = ( n3457 & n3459 ) | ( n3457 & n3461 ) | ( n3459 & n3461 ) ;
  assign n3463 = ( n3204 & n3272 ) | ( n3204 & ~n3292 ) | ( n3272 & ~n3292 ) ;
  assign n3464 = ( n3292 & ~n3293 ) | ( n3292 & n3463 ) | ( ~n3293 & n3463 ) ;
  assign n3465 = ( n3357 & n3421 ) | ( n3357 & ~n3441 ) | ( n3421 & ~n3441 ) ;
  assign n3466 = ( n3441 & ~n3442 ) | ( n3441 & n3465 ) | ( ~n3442 & n3465 ) ;
  assign n3467 = ( n3462 & n3464 ) | ( n3462 & n3466 ) | ( n3464 & n3466 ) ;
  assign n3468 = ( n3293 & n3442 ) | ( n3293 & n3467 ) | ( n3442 & n3467 ) ;
  assign n3469 = ( x403 & x404 ) | ( x403 & x405 ) | ( x404 & x405 ) ;
  assign n3470 = ( x406 & x407 ) | ( x406 & x408 ) | ( x407 & x408 ) ;
  assign n3471 = ( ~x403 & x404 ) | ( ~x403 & x405 ) | ( x404 & x405 ) ;
  assign n3472 = ( x403 & ~n3469 ) | ( x403 & n3471 ) | ( ~n3469 & n3471 ) ;
  assign n3473 = ( ~x406 & x407 ) | ( ~x406 & x408 ) | ( x407 & x408 ) ;
  assign n3474 = ( x406 & ~n3470 ) | ( x406 & n3473 ) | ( ~n3470 & n3473 ) ;
  assign n3475 = n3472 & n3474 ;
  assign n3476 = ( n3469 & n3470 ) | ( n3469 & n3475 ) | ( n3470 & n3475 ) ;
  assign n3477 = ( x409 & x410 ) | ( x409 & x411 ) | ( x410 & x411 ) ;
  assign n3478 = ( x412 & x413 ) | ( x412 & x414 ) | ( x413 & x414 ) ;
  assign n3479 = n3477 & n3478 ;
  assign n3480 = n3472 | n3474 ;
  assign n3481 = ~n3475 & n3480 ;
  assign n3482 = ( ~x409 & x410 ) | ( ~x409 & x411 ) | ( x410 & x411 ) ;
  assign n3483 = ( x409 & ~n3477 ) | ( x409 & n3482 ) | ( ~n3477 & n3482 ) ;
  assign n3484 = ( ~x412 & x413 ) | ( ~x412 & x414 ) | ( x413 & x414 ) ;
  assign n3485 = ( x412 & ~n3478 ) | ( x412 & n3484 ) | ( ~n3478 & n3484 ) ;
  assign n3486 = ( n3481 & n3483 ) | ( n3481 & n3485 ) | ( n3483 & n3485 ) ;
  assign n3487 = ( ~n3469 & n3470 ) | ( ~n3469 & n3475 ) | ( n3470 & n3475 ) ;
  assign n3488 = ( n3469 & ~n3476 ) | ( n3469 & n3487 ) | ( ~n3476 & n3487 ) ;
  assign n3489 = n3477 | n3478 ;
  assign n3490 = ~n3479 & n3489 ;
  assign n3491 = ( n3486 & n3488 ) | ( n3486 & n3490 ) | ( n3488 & n3490 ) ;
  assign n3492 = ( n3476 & n3479 ) | ( n3476 & n3491 ) | ( n3479 & n3491 ) ;
  assign n3493 = ( x391 & x392 ) | ( x391 & x393 ) | ( x392 & x393 ) ;
  assign n3494 = ( x394 & x395 ) | ( x394 & x396 ) | ( x395 & x396 ) ;
  assign n3495 = ( ~x391 & x392 ) | ( ~x391 & x393 ) | ( x392 & x393 ) ;
  assign n3496 = ( x391 & ~n3493 ) | ( x391 & n3495 ) | ( ~n3493 & n3495 ) ;
  assign n3497 = ( ~x394 & x395 ) | ( ~x394 & x396 ) | ( x395 & x396 ) ;
  assign n3498 = ( x394 & ~n3494 ) | ( x394 & n3497 ) | ( ~n3494 & n3497 ) ;
  assign n3499 = n3496 & n3498 ;
  assign n3500 = ( n3493 & n3494 ) | ( n3493 & n3499 ) | ( n3494 & n3499 ) ;
  assign n3501 = ( x397 & x398 ) | ( x397 & x399 ) | ( x398 & x399 ) ;
  assign n3502 = ( x400 & x401 ) | ( x400 & x402 ) | ( x401 & x402 ) ;
  assign n3503 = n3501 & n3502 ;
  assign n3504 = n3496 | n3498 ;
  assign n3505 = ~n3499 & n3504 ;
  assign n3506 = ( ~x397 & x398 ) | ( ~x397 & x399 ) | ( x398 & x399 ) ;
  assign n3507 = ( x397 & ~n3501 ) | ( x397 & n3506 ) | ( ~n3501 & n3506 ) ;
  assign n3508 = ( ~x400 & x401 ) | ( ~x400 & x402 ) | ( x401 & x402 ) ;
  assign n3509 = ( x400 & ~n3502 ) | ( x400 & n3508 ) | ( ~n3502 & n3508 ) ;
  assign n3510 = ( n3505 & n3507 ) | ( n3505 & n3509 ) | ( n3507 & n3509 ) ;
  assign n3511 = ( ~n3493 & n3494 ) | ( ~n3493 & n3499 ) | ( n3494 & n3499 ) ;
  assign n3512 = ( n3493 & ~n3500 ) | ( n3493 & n3511 ) | ( ~n3500 & n3511 ) ;
  assign n3513 = n3501 | n3502 ;
  assign n3514 = ~n3503 & n3513 ;
  assign n3515 = ( n3510 & n3512 ) | ( n3510 & n3514 ) | ( n3512 & n3514 ) ;
  assign n3516 = ( n3500 & n3503 ) | ( n3500 & n3515 ) | ( n3503 & n3515 ) ;
  assign n3517 = ( ~n3505 & n3507 ) | ( ~n3505 & n3509 ) | ( n3507 & n3509 ) ;
  assign n3518 = ( n3505 & ~n3510 ) | ( n3505 & n3517 ) | ( ~n3510 & n3517 ) ;
  assign n3519 = ( ~n3481 & n3483 ) | ( ~n3481 & n3485 ) | ( n3483 & n3485 ) ;
  assign n3520 = ( n3481 & ~n3486 ) | ( n3481 & n3519 ) | ( ~n3486 & n3519 ) ;
  assign n3521 = n3518 & n3520 ;
  assign n3522 = ( ~n3486 & n3488 ) | ( ~n3486 & n3490 ) | ( n3488 & n3490 ) ;
  assign n3523 = ( n3486 & ~n3491 ) | ( n3486 & n3522 ) | ( ~n3491 & n3522 ) ;
  assign n3524 = ( ~n3510 & n3512 ) | ( ~n3510 & n3514 ) | ( n3512 & n3514 ) ;
  assign n3525 = ( n3510 & ~n3515 ) | ( n3510 & n3524 ) | ( ~n3515 & n3524 ) ;
  assign n3526 = ( n3521 & n3523 ) | ( n3521 & n3525 ) | ( n3523 & n3525 ) ;
  assign n3527 = ( n3476 & n3479 ) | ( n3476 & ~n3491 ) | ( n3479 & ~n3491 ) ;
  assign n3528 = ( n3491 & ~n3492 ) | ( n3491 & n3527 ) | ( ~n3492 & n3527 ) ;
  assign n3529 = ( n3500 & n3503 ) | ( n3500 & ~n3515 ) | ( n3503 & ~n3515 ) ;
  assign n3530 = ( n3515 & ~n3516 ) | ( n3515 & n3529 ) | ( ~n3516 & n3529 ) ;
  assign n3531 = ( n3526 & n3528 ) | ( n3526 & n3530 ) | ( n3528 & n3530 ) ;
  assign n3532 = ( n3492 & n3516 ) | ( n3492 & n3531 ) | ( n3516 & n3531 ) ;
  assign n3533 = ( x382 & x383 ) | ( x382 & x384 ) | ( x383 & x384 ) ;
  assign n3534 = ( x379 & x380 ) | ( x379 & x381 ) | ( x380 & x381 ) ;
  assign n3535 = ( ~x382 & x383 ) | ( ~x382 & x384 ) | ( x383 & x384 ) ;
  assign n3536 = ( x382 & ~n3533 ) | ( x382 & n3535 ) | ( ~n3533 & n3535 ) ;
  assign n3537 = ( ~x379 & x380 ) | ( ~x379 & x381 ) | ( x380 & x381 ) ;
  assign n3538 = ( x379 & ~n3534 ) | ( x379 & n3537 ) | ( ~n3534 & n3537 ) ;
  assign n3539 = n3536 & n3538 ;
  assign n3540 = ( n3533 & n3534 ) | ( n3533 & n3539 ) | ( n3534 & n3539 ) ;
  assign n3541 = ( x385 & x386 ) | ( x385 & x387 ) | ( x386 & x387 ) ;
  assign n3542 = ( x388 & x389 ) | ( x388 & x390 ) | ( x389 & x390 ) ;
  assign n3543 = n3541 & n3542 ;
  assign n3544 = n3536 | n3538 ;
  assign n3545 = ~n3539 & n3544 ;
  assign n3546 = ( ~x385 & x386 ) | ( ~x385 & x387 ) | ( x386 & x387 ) ;
  assign n3547 = ( x385 & ~n3541 ) | ( x385 & n3546 ) | ( ~n3541 & n3546 ) ;
  assign n3548 = ( ~x388 & x389 ) | ( ~x388 & x390 ) | ( x389 & x390 ) ;
  assign n3549 = ( x388 & ~n3542 ) | ( x388 & n3548 ) | ( ~n3542 & n3548 ) ;
  assign n3550 = ( n3545 & n3547 ) | ( n3545 & n3549 ) | ( n3547 & n3549 ) ;
  assign n3551 = ( ~n3533 & n3534 ) | ( ~n3533 & n3539 ) | ( n3534 & n3539 ) ;
  assign n3552 = ( n3533 & ~n3540 ) | ( n3533 & n3551 ) | ( ~n3540 & n3551 ) ;
  assign n3553 = n3541 | n3542 ;
  assign n3554 = ~n3543 & n3553 ;
  assign n3555 = ( n3550 & n3552 ) | ( n3550 & n3554 ) | ( n3552 & n3554 ) ;
  assign n3556 = ( n3540 & n3543 ) | ( n3540 & n3555 ) | ( n3543 & n3555 ) ;
  assign n3557 = ( x370 & x371 ) | ( x370 & x372 ) | ( x371 & x372 ) ;
  assign n3558 = ( x367 & x368 ) | ( x367 & x369 ) | ( x368 & x369 ) ;
  assign n3559 = ( ~x370 & x371 ) | ( ~x370 & x372 ) | ( x371 & x372 ) ;
  assign n3560 = ( x370 & ~n3557 ) | ( x370 & n3559 ) | ( ~n3557 & n3559 ) ;
  assign n3561 = ( ~x367 & x368 ) | ( ~x367 & x369 ) | ( x368 & x369 ) ;
  assign n3562 = ( x367 & ~n3558 ) | ( x367 & n3561 ) | ( ~n3558 & n3561 ) ;
  assign n3563 = n3560 & n3562 ;
  assign n3564 = ( n3557 & n3558 ) | ( n3557 & n3563 ) | ( n3558 & n3563 ) ;
  assign n3565 = ( x373 & x374 ) | ( x373 & x375 ) | ( x374 & x375 ) ;
  assign n3566 = ( x376 & x377 ) | ( x376 & x378 ) | ( x377 & x378 ) ;
  assign n3567 = n3565 & n3566 ;
  assign n3568 = n3560 | n3562 ;
  assign n3569 = ~n3563 & n3568 ;
  assign n3570 = ( ~x373 & x374 ) | ( ~x373 & x375 ) | ( x374 & x375 ) ;
  assign n3571 = ( x373 & ~n3565 ) | ( x373 & n3570 ) | ( ~n3565 & n3570 ) ;
  assign n3572 = ( ~x376 & x377 ) | ( ~x376 & x378 ) | ( x377 & x378 ) ;
  assign n3573 = ( x376 & ~n3566 ) | ( x376 & n3572 ) | ( ~n3566 & n3572 ) ;
  assign n3574 = ( n3569 & n3571 ) | ( n3569 & n3573 ) | ( n3571 & n3573 ) ;
  assign n3575 = ( ~n3557 & n3558 ) | ( ~n3557 & n3563 ) | ( n3558 & n3563 ) ;
  assign n3576 = ( n3557 & ~n3564 ) | ( n3557 & n3575 ) | ( ~n3564 & n3575 ) ;
  assign n3577 = n3565 | n3566 ;
  assign n3578 = ~n3567 & n3577 ;
  assign n3579 = ( n3574 & n3576 ) | ( n3574 & n3578 ) | ( n3576 & n3578 ) ;
  assign n3580 = ( n3564 & n3567 ) | ( n3564 & n3579 ) | ( n3567 & n3579 ) ;
  assign n3581 = ( ~n3569 & n3571 ) | ( ~n3569 & n3573 ) | ( n3571 & n3573 ) ;
  assign n3582 = ( n3569 & ~n3574 ) | ( n3569 & n3581 ) | ( ~n3574 & n3581 ) ;
  assign n3583 = ( ~n3545 & n3547 ) | ( ~n3545 & n3549 ) | ( n3547 & n3549 ) ;
  assign n3584 = ( n3545 & ~n3550 ) | ( n3545 & n3583 ) | ( ~n3550 & n3583 ) ;
  assign n3585 = n3582 & n3584 ;
  assign n3586 = ( ~n3550 & n3552 ) | ( ~n3550 & n3554 ) | ( n3552 & n3554 ) ;
  assign n3587 = ( n3550 & ~n3555 ) | ( n3550 & n3586 ) | ( ~n3555 & n3586 ) ;
  assign n3588 = ( ~n3574 & n3576 ) | ( ~n3574 & n3578 ) | ( n3576 & n3578 ) ;
  assign n3589 = ( n3574 & ~n3579 ) | ( n3574 & n3588 ) | ( ~n3579 & n3588 ) ;
  assign n3590 = ( n3585 & n3587 ) | ( n3585 & n3589 ) | ( n3587 & n3589 ) ;
  assign n3591 = ( n3540 & n3543 ) | ( n3540 & ~n3555 ) | ( n3543 & ~n3555 ) ;
  assign n3592 = ( n3555 & ~n3556 ) | ( n3555 & n3591 ) | ( ~n3556 & n3591 ) ;
  assign n3593 = ( n3564 & n3567 ) | ( n3564 & ~n3579 ) | ( n3567 & ~n3579 ) ;
  assign n3594 = ( n3579 & ~n3580 ) | ( n3579 & n3593 ) | ( ~n3580 & n3593 ) ;
  assign n3595 = ( n3590 & n3592 ) | ( n3590 & n3594 ) | ( n3592 & n3594 ) ;
  assign n3596 = ( n3556 & n3580 ) | ( n3556 & n3595 ) | ( n3580 & n3595 ) ;
  assign n3597 = n3518 | n3520 ;
  assign n3598 = ~n3521 & n3597 ;
  assign n3599 = n3582 | n3584 ;
  assign n3600 = ~n3585 & n3599 ;
  assign n3601 = n3598 & n3600 ;
  assign n3602 = ( ~n3521 & n3523 ) | ( ~n3521 & n3525 ) | ( n3523 & n3525 ) ;
  assign n3603 = ( n3521 & ~n3526 ) | ( n3521 & n3602 ) | ( ~n3526 & n3602 ) ;
  assign n3604 = ( ~n3585 & n3587 ) | ( ~n3585 & n3589 ) | ( n3587 & n3589 ) ;
  assign n3605 = ( n3585 & ~n3590 ) | ( n3585 & n3604 ) | ( ~n3590 & n3604 ) ;
  assign n3606 = ( n3601 & n3603 ) | ( n3601 & n3605 ) | ( n3603 & n3605 ) ;
  assign n3607 = ( ~n3590 & n3592 ) | ( ~n3590 & n3594 ) | ( n3592 & n3594 ) ;
  assign n3608 = ( n3590 & ~n3595 ) | ( n3590 & n3607 ) | ( ~n3595 & n3607 ) ;
  assign n3609 = ( ~n3526 & n3528 ) | ( ~n3526 & n3530 ) | ( n3528 & n3530 ) ;
  assign n3610 = ( n3526 & ~n3531 ) | ( n3526 & n3609 ) | ( ~n3531 & n3609 ) ;
  assign n3611 = ( n3606 & n3608 ) | ( n3606 & n3610 ) | ( n3608 & n3610 ) ;
  assign n3612 = ( n3492 & n3516 ) | ( n3492 & ~n3531 ) | ( n3516 & ~n3531 ) ;
  assign n3613 = ( n3531 & ~n3532 ) | ( n3531 & n3612 ) | ( ~n3532 & n3612 ) ;
  assign n3614 = ( n3556 & n3580 ) | ( n3556 & ~n3595 ) | ( n3580 & ~n3595 ) ;
  assign n3615 = ( n3595 & ~n3596 ) | ( n3595 & n3614 ) | ( ~n3596 & n3614 ) ;
  assign n3616 = ( n3611 & n3613 ) | ( n3611 & n3615 ) | ( n3613 & n3615 ) ;
  assign n3617 = ( n3532 & n3596 ) | ( n3532 & n3616 ) | ( n3596 & n3616 ) ;
  assign n3618 = ( x457 & x458 ) | ( x457 & x459 ) | ( x458 & x459 ) ;
  assign n3619 = ( x460 & x461 ) | ( x460 & x462 ) | ( x461 & x462 ) ;
  assign n3620 = ( ~x457 & x458 ) | ( ~x457 & x459 ) | ( x458 & x459 ) ;
  assign n3621 = ( x457 & ~n3618 ) | ( x457 & n3620 ) | ( ~n3618 & n3620 ) ;
  assign n3622 = ( ~x460 & x461 ) | ( ~x460 & x462 ) | ( x461 & x462 ) ;
  assign n3623 = ( x460 & ~n3619 ) | ( x460 & n3622 ) | ( ~n3619 & n3622 ) ;
  assign n3624 = n3621 & n3623 ;
  assign n3625 = ( n3618 & n3619 ) | ( n3618 & n3624 ) | ( n3619 & n3624 ) ;
  assign n3626 = ( x454 & x455 ) | ( x454 & x456 ) | ( x455 & x456 ) ;
  assign n3627 = ( x451 & x452 ) | ( x451 & x453 ) | ( x452 & x453 ) ;
  assign n3628 = n3626 & n3627 ;
  assign n3629 = n3621 | n3623 ;
  assign n3630 = ~n3624 & n3629 ;
  assign n3631 = ( ~x454 & x455 ) | ( ~x454 & x456 ) | ( x455 & x456 ) ;
  assign n3632 = ( x454 & ~n3626 ) | ( x454 & n3631 ) | ( ~n3626 & n3631 ) ;
  assign n3633 = ( ~x451 & x452 ) | ( ~x451 & x453 ) | ( x452 & x453 ) ;
  assign n3634 = ( x451 & ~n3627 ) | ( x451 & n3633 ) | ( ~n3627 & n3633 ) ;
  assign n3635 = ( n3630 & n3632 ) | ( n3630 & n3634 ) | ( n3632 & n3634 ) ;
  assign n3636 = ( ~n3618 & n3619 ) | ( ~n3618 & n3624 ) | ( n3619 & n3624 ) ;
  assign n3637 = ( n3618 & ~n3625 ) | ( n3618 & n3636 ) | ( ~n3625 & n3636 ) ;
  assign n3638 = n3626 | n3627 ;
  assign n3639 = ~n3628 & n3638 ;
  assign n3640 = ( n3635 & n3637 ) | ( n3635 & n3639 ) | ( n3637 & n3639 ) ;
  assign n3641 = ( n3625 & n3628 ) | ( n3625 & n3640 ) | ( n3628 & n3640 ) ;
  assign n3642 = ( x439 & x440 ) | ( x439 & x441 ) | ( x440 & x441 ) ;
  assign n3643 = ( x442 & x443 ) | ( x442 & x444 ) | ( x443 & x444 ) ;
  assign n3644 = ( ~x439 & x440 ) | ( ~x439 & x441 ) | ( x440 & x441 ) ;
  assign n3645 = ( x439 & ~n3642 ) | ( x439 & n3644 ) | ( ~n3642 & n3644 ) ;
  assign n3646 = ( ~x442 & x443 ) | ( ~x442 & x444 ) | ( x443 & x444 ) ;
  assign n3647 = ( x442 & ~n3643 ) | ( x442 & n3646 ) | ( ~n3643 & n3646 ) ;
  assign n3648 = n3645 & n3647 ;
  assign n3649 = ( n3642 & n3643 ) | ( n3642 & n3648 ) | ( n3643 & n3648 ) ;
  assign n3650 = ( x448 & x449 ) | ( x448 & x450 ) | ( x449 & x450 ) ;
  assign n3651 = ( x445 & x446 ) | ( x445 & x447 ) | ( x446 & x447 ) ;
  assign n3652 = n3650 & n3651 ;
  assign n3653 = n3645 | n3647 ;
  assign n3654 = ~n3648 & n3653 ;
  assign n3655 = ( ~x448 & x449 ) | ( ~x448 & x450 ) | ( x449 & x450 ) ;
  assign n3656 = ( x448 & ~n3650 ) | ( x448 & n3655 ) | ( ~n3650 & n3655 ) ;
  assign n3657 = ( ~x445 & x446 ) | ( ~x445 & x447 ) | ( x446 & x447 ) ;
  assign n3658 = ( x445 & ~n3651 ) | ( x445 & n3657 ) | ( ~n3651 & n3657 ) ;
  assign n3659 = ( n3654 & n3656 ) | ( n3654 & n3658 ) | ( n3656 & n3658 ) ;
  assign n3660 = ( ~n3642 & n3643 ) | ( ~n3642 & n3648 ) | ( n3643 & n3648 ) ;
  assign n3661 = ( n3642 & ~n3649 ) | ( n3642 & n3660 ) | ( ~n3649 & n3660 ) ;
  assign n3662 = n3650 | n3651 ;
  assign n3663 = ~n3652 & n3662 ;
  assign n3664 = ( n3659 & n3661 ) | ( n3659 & n3663 ) | ( n3661 & n3663 ) ;
  assign n3665 = ( n3649 & n3652 ) | ( n3649 & n3664 ) | ( n3652 & n3664 ) ;
  assign n3666 = ( ~n3630 & n3632 ) | ( ~n3630 & n3634 ) | ( n3632 & n3634 ) ;
  assign n3667 = ( n3630 & ~n3635 ) | ( n3630 & n3666 ) | ( ~n3635 & n3666 ) ;
  assign n3668 = ( ~n3654 & n3656 ) | ( ~n3654 & n3658 ) | ( n3656 & n3658 ) ;
  assign n3669 = ( n3654 & ~n3659 ) | ( n3654 & n3668 ) | ( ~n3659 & n3668 ) ;
  assign n3670 = n3667 & n3669 ;
  assign n3671 = ( ~n3659 & n3661 ) | ( ~n3659 & n3663 ) | ( n3661 & n3663 ) ;
  assign n3672 = ( n3659 & ~n3664 ) | ( n3659 & n3671 ) | ( ~n3664 & n3671 ) ;
  assign n3673 = ( ~n3635 & n3637 ) | ( ~n3635 & n3639 ) | ( n3637 & n3639 ) ;
  assign n3674 = ( n3635 & ~n3640 ) | ( n3635 & n3673 ) | ( ~n3640 & n3673 ) ;
  assign n3675 = ( n3670 & n3672 ) | ( n3670 & n3674 ) | ( n3672 & n3674 ) ;
  assign n3676 = ( n3625 & n3628 ) | ( n3625 & ~n3640 ) | ( n3628 & ~n3640 ) ;
  assign n3677 = ( n3640 & ~n3641 ) | ( n3640 & n3676 ) | ( ~n3641 & n3676 ) ;
  assign n3678 = ( n3649 & n3652 ) | ( n3649 & ~n3664 ) | ( n3652 & ~n3664 ) ;
  assign n3679 = ( n3664 & ~n3665 ) | ( n3664 & n3678 ) | ( ~n3665 & n3678 ) ;
  assign n3680 = ( n3675 & n3677 ) | ( n3675 & n3679 ) | ( n3677 & n3679 ) ;
  assign n3681 = ( n3641 & n3665 ) | ( n3641 & n3680 ) | ( n3665 & n3680 ) ;
  assign n3682 = ( x418 & x419 ) | ( x418 & x420 ) | ( x419 & x420 ) ;
  assign n3683 = ( x415 & x416 ) | ( x415 & x417 ) | ( x416 & x417 ) ;
  assign n3684 = ( ~x418 & x419 ) | ( ~x418 & x420 ) | ( x419 & x420 ) ;
  assign n3685 = ( x418 & ~n3682 ) | ( x418 & n3684 ) | ( ~n3682 & n3684 ) ;
  assign n3686 = ( ~x415 & x416 ) | ( ~x415 & x417 ) | ( x416 & x417 ) ;
  assign n3687 = ( x415 & ~n3683 ) | ( x415 & n3686 ) | ( ~n3683 & n3686 ) ;
  assign n3688 = n3685 & n3687 ;
  assign n3689 = ( n3682 & n3683 ) | ( n3682 & n3688 ) | ( n3683 & n3688 ) ;
  assign n3690 = ( x421 & x422 ) | ( x421 & x423 ) | ( x422 & x423 ) ;
  assign n3691 = ( x424 & x425 ) | ( x424 & x426 ) | ( x425 & x426 ) ;
  assign n3692 = ( ~x421 & x422 ) | ( ~x421 & x423 ) | ( x422 & x423 ) ;
  assign n3693 = ( x421 & ~n3690 ) | ( x421 & n3692 ) | ( ~n3690 & n3692 ) ;
  assign n3694 = ( ~x424 & x425 ) | ( ~x424 & x426 ) | ( x425 & x426 ) ;
  assign n3695 = ( x424 & ~n3691 ) | ( x424 & n3694 ) | ( ~n3691 & n3694 ) ;
  assign n3696 = n3693 & n3695 ;
  assign n3697 = ( n3690 & n3691 ) | ( n3690 & n3696 ) | ( n3691 & n3696 ) ;
  assign n3698 = ( ~n3682 & n3683 ) | ( ~n3682 & n3688 ) | ( n3683 & n3688 ) ;
  assign n3699 = ( n3682 & ~n3689 ) | ( n3682 & n3698 ) | ( ~n3689 & n3698 ) ;
  assign n3700 = ( n3690 & n3691 ) | ( n3690 & ~n3696 ) | ( n3691 & ~n3696 ) ;
  assign n3701 = n3690 | n3691 ;
  assign n3702 = n3685 | n3687 ;
  assign n3703 = ~n3688 & n3702 ;
  assign n3704 = ( n3693 & n3695 ) | ( n3693 & n3703 ) | ( n3695 & n3703 ) ;
  assign n3705 = ( n3700 & ~n3701 ) | ( n3700 & n3704 ) | ( ~n3701 & n3704 ) ;
  assign n3706 = ~n3697 & n3700 ;
  assign n3707 = ( n3699 & n3705 ) | ( n3699 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3708 = ( n3689 & n3697 ) | ( n3689 & n3707 ) | ( n3697 & n3707 ) ;
  assign n3709 = ( x427 & x428 ) | ( x427 & x429 ) | ( x428 & x429 ) ;
  assign n3710 = ( x430 & x431 ) | ( x430 & x432 ) | ( x431 & x432 ) ;
  assign n3711 = ( ~x427 & x428 ) | ( ~x427 & x429 ) | ( x428 & x429 ) ;
  assign n3712 = ( x427 & ~n3709 ) | ( x427 & n3711 ) | ( ~n3709 & n3711 ) ;
  assign n3713 = ( ~x430 & x431 ) | ( ~x430 & x432 ) | ( x431 & x432 ) ;
  assign n3714 = ( x430 & ~n3710 ) | ( x430 & n3713 ) | ( ~n3710 & n3713 ) ;
  assign n3715 = n3712 & n3714 ;
  assign n3716 = ( n3709 & n3710 ) | ( n3709 & n3715 ) | ( n3710 & n3715 ) ;
  assign n3717 = ( x433 & x434 ) | ( x433 & x435 ) | ( x434 & x435 ) ;
  assign n3718 = ( x436 & x437 ) | ( x436 & x438 ) | ( x437 & x438 ) ;
  assign n3719 = n3717 & n3718 ;
  assign n3720 = n3712 | n3714 ;
  assign n3721 = ~n3715 & n3720 ;
  assign n3722 = ( ~x433 & x434 ) | ( ~x433 & x435 ) | ( x434 & x435 ) ;
  assign n3723 = ( x433 & ~n3717 ) | ( x433 & n3722 ) | ( ~n3717 & n3722 ) ;
  assign n3724 = ( ~x436 & x437 ) | ( ~x436 & x438 ) | ( x437 & x438 ) ;
  assign n3725 = ( x436 & ~n3718 ) | ( x436 & n3724 ) | ( ~n3718 & n3724 ) ;
  assign n3726 = ( n3721 & n3723 ) | ( n3721 & n3725 ) | ( n3723 & n3725 ) ;
  assign n3727 = ( ~n3709 & n3710 ) | ( ~n3709 & n3715 ) | ( n3710 & n3715 ) ;
  assign n3728 = ( n3709 & ~n3716 ) | ( n3709 & n3727 ) | ( ~n3716 & n3727 ) ;
  assign n3729 = n3717 | n3718 ;
  assign n3730 = ~n3719 & n3729 ;
  assign n3731 = ( n3726 & n3728 ) | ( n3726 & n3730 ) | ( n3728 & n3730 ) ;
  assign n3732 = ( n3716 & n3719 ) | ( n3716 & n3731 ) | ( n3719 & n3731 ) ;
  assign n3733 = ( ~n3721 & n3723 ) | ( ~n3721 & n3725 ) | ( n3723 & n3725 ) ;
  assign n3734 = ( n3721 & ~n3726 ) | ( n3721 & n3733 ) | ( ~n3726 & n3733 ) ;
  assign n3735 = ( n3693 & n3695 ) | ( n3693 & ~n3703 ) | ( n3695 & ~n3703 ) ;
  assign n3736 = ( n3703 & ~n3704 ) | ( n3703 & n3735 ) | ( ~n3704 & n3735 ) ;
  assign n3737 = n3734 & n3736 ;
  assign n3738 = ( ~n3726 & n3728 ) | ( ~n3726 & n3730 ) | ( n3728 & n3730 ) ;
  assign n3739 = ( n3726 & ~n3731 ) | ( n3726 & n3738 ) | ( ~n3731 & n3738 ) ;
  assign n3740 = ( ~n3699 & n3705 ) | ( ~n3699 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3741 = ( n3699 & ~n3707 ) | ( n3699 & n3740 ) | ( ~n3707 & n3740 ) ;
  assign n3742 = ( n3737 & n3739 ) | ( n3737 & n3741 ) | ( n3739 & n3741 ) ;
  assign n3743 = ( ~n3689 & n3697 ) | ( ~n3689 & n3707 ) | ( n3697 & n3707 ) ;
  assign n3744 = ( n3689 & ~n3708 ) | ( n3689 & n3743 ) | ( ~n3708 & n3743 ) ;
  assign n3745 = ( n3716 & n3719 ) | ( n3716 & ~n3731 ) | ( n3719 & ~n3731 ) ;
  assign n3746 = ( n3731 & ~n3732 ) | ( n3731 & n3745 ) | ( ~n3732 & n3745 ) ;
  assign n3747 = ( n3742 & n3744 ) | ( n3742 & n3746 ) | ( n3744 & n3746 ) ;
  assign n3748 = ( n3708 & n3732 ) | ( n3708 & n3747 ) | ( n3732 & n3747 ) ;
  assign n3749 = n3734 | n3736 ;
  assign n3750 = ~n3737 & n3749 ;
  assign n3751 = n3667 | n3669 ;
  assign n3752 = ~n3670 & n3751 ;
  assign n3753 = n3750 & n3752 ;
  assign n3754 = ( n3670 & ~n3672 ) | ( n3670 & n3674 ) | ( ~n3672 & n3674 ) ;
  assign n3755 = ( n3672 & ~n3675 ) | ( n3672 & n3754 ) | ( ~n3675 & n3754 ) ;
  assign n3756 = ( n3737 & ~n3739 ) | ( n3737 & n3741 ) | ( ~n3739 & n3741 ) ;
  assign n3757 = ( n3739 & ~n3742 ) | ( n3739 & n3756 ) | ( ~n3742 & n3756 ) ;
  assign n3758 = ( n3753 & n3755 ) | ( n3753 & n3757 ) | ( n3755 & n3757 ) ;
  assign n3759 = ( ~n3742 & n3744 ) | ( ~n3742 & n3746 ) | ( n3744 & n3746 ) ;
  assign n3760 = ( n3742 & ~n3747 ) | ( n3742 & n3759 ) | ( ~n3747 & n3759 ) ;
  assign n3761 = ( ~n3675 & n3677 ) | ( ~n3675 & n3679 ) | ( n3677 & n3679 ) ;
  assign n3762 = ( n3675 & ~n3680 ) | ( n3675 & n3761 ) | ( ~n3680 & n3761 ) ;
  assign n3763 = ( n3758 & n3760 ) | ( n3758 & n3762 ) | ( n3760 & n3762 ) ;
  assign n3764 = ( n3641 & n3665 ) | ( n3641 & ~n3680 ) | ( n3665 & ~n3680 ) ;
  assign n3765 = ( n3680 & ~n3681 ) | ( n3680 & n3764 ) | ( ~n3681 & n3764 ) ;
  assign n3766 = ( ~n3708 & n3732 ) | ( ~n3708 & n3747 ) | ( n3732 & n3747 ) ;
  assign n3767 = ( n3708 & ~n3748 ) | ( n3708 & n3766 ) | ( ~n3748 & n3766 ) ;
  assign n3768 = ( n3763 & n3765 ) | ( n3763 & n3767 ) | ( n3765 & n3767 ) ;
  assign n3769 = ( n3681 & n3748 ) | ( n3681 & n3768 ) | ( n3748 & n3768 ) ;
  assign n3770 = n3598 | n3600 ;
  assign n3771 = ~n3601 & n3770 ;
  assign n3772 = n3750 | n3752 ;
  assign n3773 = ~n3753 & n3772 ;
  assign n3774 = n3771 & n3773 ;
  assign n3775 = ( n3601 & ~n3603 ) | ( n3601 & n3605 ) | ( ~n3603 & n3605 ) ;
  assign n3776 = ( n3603 & ~n3606 ) | ( n3603 & n3775 ) | ( ~n3606 & n3775 ) ;
  assign n3777 = ( ~n3753 & n3755 ) | ( ~n3753 & n3757 ) | ( n3755 & n3757 ) ;
  assign n3778 = ( n3753 & ~n3758 ) | ( n3753 & n3777 ) | ( ~n3758 & n3777 ) ;
  assign n3779 = ( n3774 & n3776 ) | ( n3774 & n3778 ) | ( n3776 & n3778 ) ;
  assign n3780 = ( ~n3758 & n3760 ) | ( ~n3758 & n3762 ) | ( n3760 & n3762 ) ;
  assign n3781 = ( n3758 & ~n3763 ) | ( n3758 & n3780 ) | ( ~n3763 & n3780 ) ;
  assign n3782 = ( ~n3606 & n3608 ) | ( ~n3606 & n3610 ) | ( n3608 & n3610 ) ;
  assign n3783 = ( n3606 & ~n3611 ) | ( n3606 & n3782 ) | ( ~n3611 & n3782 ) ;
  assign n3784 = ( n3779 & n3781 ) | ( n3779 & n3783 ) | ( n3781 & n3783 ) ;
  assign n3785 = ( n3611 & ~n3613 ) | ( n3611 & n3615 ) | ( ~n3613 & n3615 ) ;
  assign n3786 = ( n3613 & ~n3616 ) | ( n3613 & n3785 ) | ( ~n3616 & n3785 ) ;
  assign n3787 = ( ~n3763 & n3765 ) | ( ~n3763 & n3767 ) | ( n3765 & n3767 ) ;
  assign n3788 = ( n3763 & ~n3768 ) | ( n3763 & n3787 ) | ( ~n3768 & n3787 ) ;
  assign n3789 = ( n3784 & n3786 ) | ( n3784 & n3788 ) | ( n3786 & n3788 ) ;
  assign n3790 = ( ~n3532 & n3596 ) | ( ~n3532 & n3616 ) | ( n3596 & n3616 ) ;
  assign n3791 = ( n3532 & ~n3617 ) | ( n3532 & n3790 ) | ( ~n3617 & n3790 ) ;
  assign n3792 = ( n3681 & n3748 ) | ( n3681 & ~n3768 ) | ( n3748 & ~n3768 ) ;
  assign n3793 = ( n3768 & ~n3769 ) | ( n3768 & n3792 ) | ( ~n3769 & n3792 ) ;
  assign n3794 = ( n3789 & n3791 ) | ( n3789 & n3793 ) | ( n3791 & n3793 ) ;
  assign n3795 = ( n3617 & n3769 ) | ( n3617 & n3794 ) | ( n3769 & n3794 ) ;
  assign n3796 = n3771 | n3773 ;
  assign n3797 = ~n3774 & n3796 ;
  assign n3798 = n3444 | n3446 ;
  assign n3799 = ~n3447 & n3798 ;
  assign n3800 = n3797 & n3799 ;
  assign n3801 = ( n3774 & ~n3776 ) | ( n3774 & n3778 ) | ( ~n3776 & n3778 ) ;
  assign n3802 = ( n3776 & ~n3779 ) | ( n3776 & n3801 ) | ( ~n3779 & n3801 ) ;
  assign n3803 = ( ~n3447 & n3449 ) | ( ~n3447 & n3451 ) | ( n3449 & n3451 ) ;
  assign n3804 = ( n3447 & ~n3452 ) | ( n3447 & n3803 ) | ( ~n3452 & n3803 ) ;
  assign n3805 = ( n3800 & n3802 ) | ( n3800 & n3804 ) | ( n3802 & n3804 ) ;
  assign n3806 = ( n3452 & ~n3454 ) | ( n3452 & n3456 ) | ( ~n3454 & n3456 ) ;
  assign n3807 = ( n3454 & ~n3457 ) | ( n3454 & n3806 ) | ( ~n3457 & n3806 ) ;
  assign n3808 = ( ~n3779 & n3781 ) | ( ~n3779 & n3783 ) | ( n3781 & n3783 ) ;
  assign n3809 = ( n3779 & ~n3784 ) | ( n3779 & n3808 ) | ( ~n3784 & n3808 ) ;
  assign n3810 = ( n3805 & n3807 ) | ( n3805 & n3809 ) | ( n3807 & n3809 ) ;
  assign n3811 = ( ~n3457 & n3459 ) | ( ~n3457 & n3461 ) | ( n3459 & n3461 ) ;
  assign n3812 = ( n3457 & ~n3462 ) | ( n3457 & n3811 ) | ( ~n3462 & n3811 ) ;
  assign n3813 = ( n3784 & ~n3786 ) | ( n3784 & n3788 ) | ( ~n3786 & n3788 ) ;
  assign n3814 = ( n3786 & ~n3789 ) | ( n3786 & n3813 ) | ( ~n3789 & n3813 ) ;
  assign n3815 = ( n3810 & n3812 ) | ( n3810 & n3814 ) | ( n3812 & n3814 ) ;
  assign n3816 = ( ~n3789 & n3791 ) | ( ~n3789 & n3793 ) | ( n3791 & n3793 ) ;
  assign n3817 = ( n3789 & ~n3794 ) | ( n3789 & n3816 ) | ( ~n3794 & n3816 ) ;
  assign n3818 = ( ~n3462 & n3464 ) | ( ~n3462 & n3466 ) | ( n3464 & n3466 ) ;
  assign n3819 = ( n3462 & ~n3467 ) | ( n3462 & n3818 ) | ( ~n3467 & n3818 ) ;
  assign n3820 = ( n3815 & n3817 ) | ( n3815 & n3819 ) | ( n3817 & n3819 ) ;
  assign n3821 = ( ~n3293 & n3442 ) | ( ~n3293 & n3467 ) | ( n3442 & n3467 ) ;
  assign n3822 = ( n3293 & ~n3468 ) | ( n3293 & n3821 ) | ( ~n3468 & n3821 ) ;
  assign n3823 = ( n3617 & n3769 ) | ( n3617 & ~n3794 ) | ( n3769 & ~n3794 ) ;
  assign n3824 = ( n3794 & ~n3795 ) | ( n3794 & n3823 ) | ( ~n3795 & n3823 ) ;
  assign n3825 = ( n3820 & n3822 ) | ( n3820 & n3824 ) | ( n3822 & n3824 ) ;
  assign n3826 = ( n3468 & n3795 ) | ( n3468 & n3825 ) | ( n3795 & n3825 ) ;
  assign n3827 = ( n3109 & ~n3111 ) | ( n3109 & n3113 ) | ( ~n3111 & n3113 ) ;
  assign n3828 = ( n3111 & ~n3114 ) | ( n3111 & n3827 ) | ( ~n3114 & n3827 ) ;
  assign n3829 = n3106 | n3108 ;
  assign n3830 = ~n3109 & n3829 ;
  assign n3831 = n3797 | n3799 ;
  assign n3832 = ~n3800 & n3831 ;
  assign n3833 = n3830 & n3832 ;
  assign n3834 = ( n3800 & ~n3802 ) | ( n3800 & n3804 ) | ( ~n3802 & n3804 ) ;
  assign n3835 = ( n3802 & ~n3805 ) | ( n3802 & n3834 ) | ( ~n3805 & n3834 ) ;
  assign n3836 = n3833 | n3835 ;
  assign n3837 = ( n3802 & n3804 ) | ( n3802 & n3833 ) | ( n3804 & n3833 ) ;
  assign n3838 = ( n3802 & n3804 ) | ( n3802 & ~n3833 ) | ( n3804 & ~n3833 ) ;
  assign n3839 = n3837 & ~n3838 ;
  assign n3840 = ( n3828 & n3836 ) | ( n3828 & n3839 ) | ( n3836 & n3839 ) ;
  assign n3841 = ( n3114 & ~n3116 ) | ( n3114 & n3118 ) | ( ~n3116 & n3118 ) ;
  assign n3842 = ( n3116 & ~n3119 ) | ( n3116 & n3841 ) | ( ~n3119 & n3841 ) ;
  assign n3843 = ( ~n3805 & n3807 ) | ( ~n3805 & n3809 ) | ( n3807 & n3809 ) ;
  assign n3844 = ( n3805 & ~n3810 ) | ( n3805 & n3843 ) | ( ~n3810 & n3843 ) ;
  assign n3845 = ( n3840 & n3842 ) | ( n3840 & n3844 ) | ( n3842 & n3844 ) ;
  assign n3846 = ( n3119 & ~n3121 ) | ( n3119 & n3123 ) | ( ~n3121 & n3123 ) ;
  assign n3847 = ( n3121 & ~n3124 ) | ( n3121 & n3846 ) | ( ~n3124 & n3846 ) ;
  assign n3848 = ( ~n3810 & n3812 ) | ( ~n3810 & n3814 ) | ( n3812 & n3814 ) ;
  assign n3849 = ( n3810 & ~n3815 ) | ( n3810 & n3848 ) | ( ~n3815 & n3848 ) ;
  assign n3850 = ( n3845 & n3847 ) | ( n3845 & n3849 ) | ( n3847 & n3849 ) ;
  assign n3851 = ( ~n3124 & n3126 ) | ( ~n3124 & n3128 ) | ( n3126 & n3128 ) ;
  assign n3852 = ( n3124 & ~n3129 ) | ( n3124 & n3851 ) | ( ~n3129 & n3851 ) ;
  assign n3853 = ( ~n3815 & n3817 ) | ( ~n3815 & n3819 ) | ( n3817 & n3819 ) ;
  assign n3854 = ( n3815 & ~n3820 ) | ( n3815 & n3853 ) | ( ~n3820 & n3853 ) ;
  assign n3855 = ( n3850 & n3852 ) | ( n3850 & n3854 ) | ( n3852 & n3854 ) ;
  assign n3856 = ( ~n3820 & n3822 ) | ( ~n3820 & n3824 ) | ( n3822 & n3824 ) ;
  assign n3857 = ( n3820 & ~n3825 ) | ( n3820 & n3856 ) | ( ~n3825 & n3856 ) ;
  assign n3858 = ( n3129 & ~n3131 ) | ( n3129 & n3133 ) | ( ~n3131 & n3133 ) ;
  assign n3859 = ( n3131 & ~n3134 ) | ( n3131 & n3858 ) | ( ~n3134 & n3858 ) ;
  assign n3860 = ( n3855 & n3857 ) | ( n3855 & n3859 ) | ( n3857 & n3859 ) ;
  assign n3861 = ( n2771 & n3104 ) | ( n2771 & ~n3134 ) | ( n3104 & ~n3134 ) ;
  assign n3862 = ( n3134 & ~n3135 ) | ( n3134 & n3861 ) | ( ~n3135 & n3861 ) ;
  assign n3863 = ( n3468 & n3795 ) | ( n3468 & ~n3825 ) | ( n3795 & ~n3825 ) ;
  assign n3864 = ( n3825 & ~n3826 ) | ( n3825 & n3863 ) | ( ~n3826 & n3863 ) ;
  assign n3865 = ( n3860 & n3862 ) | ( n3860 & n3864 ) | ( n3862 & n3864 ) ;
  assign n3866 = ( n3135 & n3826 ) | ( n3135 & n3865 ) | ( n3826 & n3865 ) ;
  assign n3867 = ( ~n3135 & n3826 ) | ( ~n3135 & n3865 ) | ( n3826 & n3865 ) ;
  assign n3868 = ( n3135 & ~n3866 ) | ( n3135 & n3867 ) | ( ~n3866 & n3867 ) ;
  assign n3869 = ( ~x862 & x863 ) | ( ~x862 & x864 ) | ( x863 & x864 ) ;
  assign n3870 = ( x862 & x863 ) | ( x862 & x864 ) | ( x863 & x864 ) ;
  assign n3871 = ( x862 & n3869 ) | ( x862 & ~n3870 ) | ( n3869 & ~n3870 ) ;
  assign n3872 = ( ~x859 & x860 ) | ( ~x859 & x861 ) | ( x860 & x861 ) ;
  assign n3873 = ( x859 & x860 ) | ( x859 & x861 ) | ( x860 & x861 ) ;
  assign n3874 = ( x859 & n3872 ) | ( x859 & ~n3873 ) | ( n3872 & ~n3873 ) ;
  assign n3875 = n3871 | n3874 ;
  assign n3876 = n3871 & n3874 ;
  assign n3877 = n3875 & ~n3876 ;
  assign n3878 = ( ~x868 & x869 ) | ( ~x868 & x870 ) | ( x869 & x870 ) ;
  assign n3879 = ( x868 & x869 ) | ( x868 & x870 ) | ( x869 & x870 ) ;
  assign n3880 = ( x868 & n3878 ) | ( x868 & ~n3879 ) | ( n3878 & ~n3879 ) ;
  assign n3881 = ( ~x865 & x866 ) | ( ~x865 & x867 ) | ( x866 & x867 ) ;
  assign n3882 = ( x865 & x866 ) | ( x865 & x867 ) | ( x866 & x867 ) ;
  assign n3883 = ( x865 & n3881 ) | ( x865 & ~n3882 ) | ( n3881 & ~n3882 ) ;
  assign n3884 = ( ~n3877 & n3880 ) | ( ~n3877 & n3883 ) | ( n3880 & n3883 ) ;
  assign n3885 = ( n3877 & n3880 ) | ( n3877 & n3883 ) | ( n3880 & n3883 ) ;
  assign n3886 = ( n3877 & n3884 ) | ( n3877 & ~n3885 ) | ( n3884 & ~n3885 ) ;
  assign n3887 = ( ~x850 & x851 ) | ( ~x850 & x852 ) | ( x851 & x852 ) ;
  assign n3888 = ( x850 & x851 ) | ( x850 & x852 ) | ( x851 & x852 ) ;
  assign n3889 = ( x850 & n3887 ) | ( x850 & ~n3888 ) | ( n3887 & ~n3888 ) ;
  assign n3890 = ( ~x847 & x848 ) | ( ~x847 & x849 ) | ( x848 & x849 ) ;
  assign n3891 = ( x847 & x848 ) | ( x847 & x849 ) | ( x848 & x849 ) ;
  assign n3892 = ( x847 & n3890 ) | ( x847 & ~n3891 ) | ( n3890 & ~n3891 ) ;
  assign n3893 = n3889 | n3892 ;
  assign n3894 = n3889 & n3892 ;
  assign n3895 = n3893 & ~n3894 ;
  assign n3896 = ( ~x856 & x857 ) | ( ~x856 & x858 ) | ( x857 & x858 ) ;
  assign n3897 = ( x856 & x857 ) | ( x856 & x858 ) | ( x857 & x858 ) ;
  assign n3898 = ( x856 & n3896 ) | ( x856 & ~n3897 ) | ( n3896 & ~n3897 ) ;
  assign n3899 = ( ~x853 & x854 ) | ( ~x853 & x855 ) | ( x854 & x855 ) ;
  assign n3900 = ( x853 & x854 ) | ( x853 & x855 ) | ( x854 & x855 ) ;
  assign n3901 = ( x853 & n3899 ) | ( x853 & ~n3900 ) | ( n3899 & ~n3900 ) ;
  assign n3902 = n3898 & n3901 ;
  assign n3903 = n3898 | n3901 ;
  assign n3904 = ~n3902 & n3903 ;
  assign n3905 = n3895 | n3904 ;
  assign n3906 = n3895 & n3904 ;
  assign n3907 = n3905 & ~n3906 ;
  assign n3908 = ( ~x886 & x887 ) | ( ~x886 & x888 ) | ( x887 & x888 ) ;
  assign n3909 = ( x886 & x887 ) | ( x886 & x888 ) | ( x887 & x888 ) ;
  assign n3910 = ( x886 & n3908 ) | ( x886 & ~n3909 ) | ( n3908 & ~n3909 ) ;
  assign n3911 = ( ~x883 & x884 ) | ( ~x883 & x885 ) | ( x884 & x885 ) ;
  assign n3912 = ( x883 & x884 ) | ( x883 & x885 ) | ( x884 & x885 ) ;
  assign n3913 = ( x883 & n3911 ) | ( x883 & ~n3912 ) | ( n3911 & ~n3912 ) ;
  assign n3914 = n3910 & n3913 ;
  assign n3915 = n3910 | n3913 ;
  assign n3916 = ~n3914 & n3915 ;
  assign n3917 = ( ~x892 & x893 ) | ( ~x892 & x894 ) | ( x893 & x894 ) ;
  assign n3918 = ( x892 & x893 ) | ( x892 & x894 ) | ( x893 & x894 ) ;
  assign n3919 = ( x892 & n3917 ) | ( x892 & ~n3918 ) | ( n3917 & ~n3918 ) ;
  assign n3920 = ( ~x889 & x890 ) | ( ~x889 & x891 ) | ( x890 & x891 ) ;
  assign n3921 = ( x889 & x890 ) | ( x889 & x891 ) | ( x890 & x891 ) ;
  assign n3922 = ( x889 & n3920 ) | ( x889 & ~n3921 ) | ( n3920 & ~n3921 ) ;
  assign n3923 = ( n3916 & n3919 ) | ( n3916 & n3922 ) | ( n3919 & n3922 ) ;
  assign n3924 = ( ~n3916 & n3919 ) | ( ~n3916 & n3922 ) | ( n3919 & n3922 ) ;
  assign n3925 = ( n3916 & ~n3923 ) | ( n3916 & n3924 ) | ( ~n3923 & n3924 ) ;
  assign n3926 = ( ~x874 & x875 ) | ( ~x874 & x876 ) | ( x875 & x876 ) ;
  assign n3927 = ( x874 & x875 ) | ( x874 & x876 ) | ( x875 & x876 ) ;
  assign n3928 = ( x874 & n3926 ) | ( x874 & ~n3927 ) | ( n3926 & ~n3927 ) ;
  assign n3929 = ( ~x871 & x872 ) | ( ~x871 & x873 ) | ( x872 & x873 ) ;
  assign n3930 = ( x871 & x872 ) | ( x871 & x873 ) | ( x872 & x873 ) ;
  assign n3931 = ( x871 & n3929 ) | ( x871 & ~n3930 ) | ( n3929 & ~n3930 ) ;
  assign n3932 = n3928 & n3931 ;
  assign n3933 = n3928 | n3931 ;
  assign n3934 = ~n3932 & n3933 ;
  assign n3935 = ( ~x880 & x881 ) | ( ~x880 & x882 ) | ( x881 & x882 ) ;
  assign n3936 = ( x880 & x881 ) | ( x880 & x882 ) | ( x881 & x882 ) ;
  assign n3937 = ( x880 & n3935 ) | ( x880 & ~n3936 ) | ( n3935 & ~n3936 ) ;
  assign n3938 = ( ~x877 & x878 ) | ( ~x877 & x879 ) | ( x878 & x879 ) ;
  assign n3939 = ( x877 & x878 ) | ( x877 & x879 ) | ( x878 & x879 ) ;
  assign n3940 = ( x877 & n3938 ) | ( x877 & ~n3939 ) | ( n3938 & ~n3939 ) ;
  assign n3941 = ( n3934 & n3937 ) | ( n3934 & n3940 ) | ( n3937 & n3940 ) ;
  assign n3942 = ( ~n3934 & n3937 ) | ( ~n3934 & n3940 ) | ( n3937 & n3940 ) ;
  assign n3943 = ( n3934 & ~n3941 ) | ( n3934 & n3942 ) | ( ~n3941 & n3942 ) ;
  assign n3944 = n3925 & n3943 ;
  assign n3945 = n3925 | n3943 ;
  assign n3946 = ~n3944 & n3945 ;
  assign n3947 = ( n3886 & n3907 ) | ( n3886 & n3946 ) | ( n3907 & n3946 ) ;
  assign n3948 = ( ~n3886 & n3907 ) | ( ~n3886 & n3946 ) | ( n3907 & n3946 ) ;
  assign n3949 = ( n3886 & ~n3947 ) | ( n3886 & n3948 ) | ( ~n3947 & n3948 ) ;
  assign n3950 = ( ~x922 & x923 ) | ( ~x922 & x924 ) | ( x923 & x924 ) ;
  assign n3951 = ( x922 & x923 ) | ( x922 & x924 ) | ( x923 & x924 ) ;
  assign n3952 = ( x922 & n3950 ) | ( x922 & ~n3951 ) | ( n3950 & ~n3951 ) ;
  assign n3953 = ( ~x919 & x920 ) | ( ~x919 & x921 ) | ( x920 & x921 ) ;
  assign n3954 = ( x919 & x920 ) | ( x919 & x921 ) | ( x920 & x921 ) ;
  assign n3955 = ( x919 & n3953 ) | ( x919 & ~n3954 ) | ( n3953 & ~n3954 ) ;
  assign n3956 = n3952 & n3955 ;
  assign n3957 = n3952 | n3955 ;
  assign n3958 = ~n3956 & n3957 ;
  assign n3959 = ( ~x925 & x926 ) | ( ~x925 & x927 ) | ( x926 & x927 ) ;
  assign n3960 = ( x925 & x926 ) | ( x925 & x927 ) | ( x926 & x927 ) ;
  assign n3961 = ( x925 & n3959 ) | ( x925 & ~n3960 ) | ( n3959 & ~n3960 ) ;
  assign n3962 = ( ~x928 & x929 ) | ( ~x928 & x930 ) | ( x929 & x930 ) ;
  assign n3963 = ( x928 & x929 ) | ( x928 & x930 ) | ( x929 & x930 ) ;
  assign n3964 = ( x928 & n3962 ) | ( x928 & ~n3963 ) | ( n3962 & ~n3963 ) ;
  assign n3965 = ( n3958 & n3961 ) | ( n3958 & n3964 ) | ( n3961 & n3964 ) ;
  assign n3966 = ( ~n3958 & n3961 ) | ( ~n3958 & n3964 ) | ( n3961 & n3964 ) ;
  assign n3967 = ( n3958 & ~n3965 ) | ( n3958 & n3966 ) | ( ~n3965 & n3966 ) ;
  assign n3968 = ( ~x931 & x932 ) | ( ~x931 & x933 ) | ( x932 & x933 ) ;
  assign n3969 = ( x931 & x932 ) | ( x931 & x933 ) | ( x932 & x933 ) ;
  assign n3970 = ( x931 & n3968 ) | ( x931 & ~n3969 ) | ( n3968 & ~n3969 ) ;
  assign n3971 = ( ~x934 & x935 ) | ( ~x934 & x936 ) | ( x935 & x936 ) ;
  assign n3972 = ( x934 & x935 ) | ( x934 & x936 ) | ( x935 & x936 ) ;
  assign n3973 = ( x934 & n3971 ) | ( x934 & ~n3972 ) | ( n3971 & ~n3972 ) ;
  assign n3974 = n3970 & n3973 ;
  assign n3975 = n3970 | n3973 ;
  assign n3976 = ~n3974 & n3975 ;
  assign n3977 = ( ~x940 & x941 ) | ( ~x940 & x942 ) | ( x941 & x942 ) ;
  assign n3978 = ( x940 & x941 ) | ( x940 & x942 ) | ( x941 & x942 ) ;
  assign n3979 = ( x940 & n3977 ) | ( x940 & ~n3978 ) | ( n3977 & ~n3978 ) ;
  assign n3980 = ( ~x937 & x938 ) | ( ~x937 & x939 ) | ( x938 & x939 ) ;
  assign n3981 = ( x937 & x938 ) | ( x937 & x939 ) | ( x938 & x939 ) ;
  assign n3982 = ( x937 & n3980 ) | ( x937 & ~n3981 ) | ( n3980 & ~n3981 ) ;
  assign n3983 = ( n3976 & n3979 ) | ( n3976 & n3982 ) | ( n3979 & n3982 ) ;
  assign n3984 = ( ~n3976 & n3979 ) | ( ~n3976 & n3982 ) | ( n3979 & n3982 ) ;
  assign n3985 = ( n3976 & ~n3983 ) | ( n3976 & n3984 ) | ( ~n3983 & n3984 ) ;
  assign n3986 = n3967 & n3985 ;
  assign n3987 = n3967 | n3985 ;
  assign n3988 = ~n3986 & n3987 ;
  assign n3989 = ( ~x895 & x896 ) | ( ~x895 & x897 ) | ( x896 & x897 ) ;
  assign n3990 = ( x895 & x896 ) | ( x895 & x897 ) | ( x896 & x897 ) ;
  assign n3991 = ( x895 & n3989 ) | ( x895 & ~n3990 ) | ( n3989 & ~n3990 ) ;
  assign n3992 = ( ~x898 & x899 ) | ( ~x898 & x900 ) | ( x899 & x900 ) ;
  assign n3993 = ( x898 & x899 ) | ( x898 & x900 ) | ( x899 & x900 ) ;
  assign n3994 = ( x898 & n3992 ) | ( x898 & ~n3993 ) | ( n3992 & ~n3993 ) ;
  assign n3995 = n3991 & n3994 ;
  assign n3996 = n3991 | n3994 ;
  assign n3997 = ~n3995 & n3996 ;
  assign n3998 = ( ~x904 & x905 ) | ( ~x904 & x906 ) | ( x905 & x906 ) ;
  assign n3999 = ( x904 & x905 ) | ( x904 & x906 ) | ( x905 & x906 ) ;
  assign n4000 = ( x904 & n3998 ) | ( x904 & ~n3999 ) | ( n3998 & ~n3999 ) ;
  assign n4001 = ( ~x901 & x902 ) | ( ~x901 & x903 ) | ( x902 & x903 ) ;
  assign n4002 = ( x901 & x902 ) | ( x901 & x903 ) | ( x902 & x903 ) ;
  assign n4003 = ( x901 & n4001 ) | ( x901 & ~n4002 ) | ( n4001 & ~n4002 ) ;
  assign n4004 = ( n3997 & n4000 ) | ( n3997 & n4003 ) | ( n4000 & n4003 ) ;
  assign n4005 = ( ~n3997 & n4000 ) | ( ~n3997 & n4003 ) | ( n4000 & n4003 ) ;
  assign n4006 = ( n3997 & ~n4004 ) | ( n3997 & n4005 ) | ( ~n4004 & n4005 ) ;
  assign n4007 = ( ~x910 & x911 ) | ( ~x910 & x912 ) | ( x911 & x912 ) ;
  assign n4008 = ( x910 & x911 ) | ( x910 & x912 ) | ( x911 & x912 ) ;
  assign n4009 = ( x910 & n4007 ) | ( x910 & ~n4008 ) | ( n4007 & ~n4008 ) ;
  assign n4010 = ( ~x907 & x908 ) | ( ~x907 & x909 ) | ( x908 & x909 ) ;
  assign n4011 = ( x907 & x908 ) | ( x907 & x909 ) | ( x908 & x909 ) ;
  assign n4012 = ( x907 & n4010 ) | ( x907 & ~n4011 ) | ( n4010 & ~n4011 ) ;
  assign n4013 = n4009 & n4012 ;
  assign n4014 = n4009 | n4012 ;
  assign n4015 = ~n4013 & n4014 ;
  assign n4016 = ( ~x913 & x914 ) | ( ~x913 & x915 ) | ( x914 & x915 ) ;
  assign n4017 = ( x913 & x914 ) | ( x913 & x915 ) | ( x914 & x915 ) ;
  assign n4018 = ( x913 & n4016 ) | ( x913 & ~n4017 ) | ( n4016 & ~n4017 ) ;
  assign n4019 = ( ~x916 & x917 ) | ( ~x916 & x918 ) | ( x917 & x918 ) ;
  assign n4020 = ( x916 & x917 ) | ( x916 & x918 ) | ( x917 & x918 ) ;
  assign n4021 = ( x916 & n4019 ) | ( x916 & ~n4020 ) | ( n4019 & ~n4020 ) ;
  assign n4022 = ( n4015 & n4018 ) | ( n4015 & n4021 ) | ( n4018 & n4021 ) ;
  assign n4023 = ( ~n4015 & n4018 ) | ( ~n4015 & n4021 ) | ( n4018 & n4021 ) ;
  assign n4024 = ( n4015 & ~n4022 ) | ( n4015 & n4023 ) | ( ~n4022 & n4023 ) ;
  assign n4025 = n4006 & n4024 ;
  assign n4026 = n4006 | n4024 ;
  assign n4027 = ~n4025 & n4026 ;
  assign n4028 = n3988 & n4027 ;
  assign n4029 = n3988 | n4027 ;
  assign n4030 = ~n4028 & n4029 ;
  assign n4031 = n3949 & n4030 ;
  assign n4032 = n3949 | n4030 ;
  assign n4033 = ~n4031 & n4032 ;
  assign n4034 = ( ~x0 & x1 ) | ( ~x0 & x2 ) | ( x1 & x2 ) ;
  assign n4035 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n4036 = ( x0 & n4034 ) | ( x0 & ~n4035 ) | ( n4034 & ~n4035 ) ;
  assign n4037 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n4038 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n4039 = ( x3 & n4037 ) | ( x3 & ~n4038 ) | ( n4037 & ~n4038 ) ;
  assign n4040 = ( x6 & n4036 ) | ( x6 & n4039 ) | ( n4036 & n4039 ) ;
  assign n4041 = ( ~x6 & n4036 ) | ( ~x6 & n4039 ) | ( n4036 & n4039 ) ;
  assign n4042 = ( x6 & ~n4040 ) | ( x6 & n4041 ) | ( ~n4040 & n4041 ) ;
  assign n4043 = x997 & x998 ;
  assign n4044 = x997 | x998 ;
  assign n4045 = ~n4043 & n4044 ;
  assign n4046 = ( x999 & ~n4042 ) | ( x999 & n4045 ) | ( ~n4042 & n4045 ) ;
  assign n4047 = ( x999 & n4042 ) | ( x999 & n4045 ) | ( n4042 & n4045 ) ;
  assign n4048 = ( n4042 & n4046 ) | ( n4042 & ~n4047 ) | ( n4046 & ~n4047 ) ;
  assign n4049 = ( ~x994 & x995 ) | ( ~x994 & x996 ) | ( x995 & x996 ) ;
  assign n4050 = ( x994 & x995 ) | ( x994 & x996 ) | ( x995 & x996 ) ;
  assign n4051 = ( x994 & n4049 ) | ( x994 & ~n4050 ) | ( n4049 & ~n4050 ) ;
  assign n4052 = ( ~x991 & x992 ) | ( ~x991 & x993 ) | ( x992 & x993 ) ;
  assign n4053 = ( x991 & x992 ) | ( x991 & x993 ) | ( x992 & x993 ) ;
  assign n4054 = ( x991 & n4052 ) | ( x991 & ~n4053 ) | ( n4052 & ~n4053 ) ;
  assign n4055 = ( n4048 & n4051 ) | ( n4048 & n4054 ) | ( n4051 & n4054 ) ;
  assign n4056 = ( ~n4048 & n4051 ) | ( ~n4048 & n4054 ) | ( n4051 & n4054 ) ;
  assign n4057 = ( n4048 & ~n4055 ) | ( n4048 & n4056 ) | ( ~n4055 & n4056 ) ;
  assign n4058 = ( ~x7 & x8 ) | ( ~x7 & x9 ) | ( x8 & x9 ) ;
  assign n4059 = ( x7 & x8 ) | ( x7 & x9 ) | ( x8 & x9 ) ;
  assign n4060 = ( x7 & n4058 ) | ( x7 & ~n4059 ) | ( n4058 & ~n4059 ) ;
  assign n4061 = ( ~x10 & x11 ) | ( ~x10 & x12 ) | ( x11 & x12 ) ;
  assign n4062 = ( x10 & x11 ) | ( x10 & x12 ) | ( x11 & x12 ) ;
  assign n4063 = ( x10 & n4061 ) | ( x10 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = n4060 | n4063 ;
  assign n4065 = n4060 & n4063 ;
  assign n4066 = n4064 & ~n4065 ;
  assign n4067 = ( ~x16 & x17 ) | ( ~x16 & x18 ) | ( x17 & x18 ) ;
  assign n4068 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n4069 = ( x16 & n4067 ) | ( x16 & ~n4068 ) | ( n4067 & ~n4068 ) ;
  assign n4070 = ( ~x13 & x14 ) | ( ~x13 & x15 ) | ( x14 & x15 ) ;
  assign n4071 = ( x13 & x14 ) | ( x13 & x15 ) | ( x14 & x15 ) ;
  assign n4072 = ( x13 & n4070 ) | ( x13 & ~n4071 ) | ( n4070 & ~n4071 ) ;
  assign n4073 = ( n4066 & n4069 ) | ( n4066 & n4072 ) | ( n4069 & n4072 ) ;
  assign n4074 = ( ~n4066 & n4069 ) | ( ~n4066 & n4072 ) | ( n4069 & n4072 ) ;
  assign n4075 = ( n4066 & ~n4073 ) | ( n4066 & n4074 ) | ( ~n4073 & n4074 ) ;
  assign n4076 = ( ~x19 & x20 ) | ( ~x19 & x21 ) | ( x20 & x21 ) ;
  assign n4077 = ( x19 & x20 ) | ( x19 & x21 ) | ( x20 & x21 ) ;
  assign n4078 = ( x19 & n4076 ) | ( x19 & ~n4077 ) | ( n4076 & ~n4077 ) ;
  assign n4079 = ( ~x22 & x23 ) | ( ~x22 & x24 ) | ( x23 & x24 ) ;
  assign n4080 = ( x22 & x23 ) | ( x22 & x24 ) | ( x23 & x24 ) ;
  assign n4081 = ( x22 & n4079 ) | ( x22 & ~n4080 ) | ( n4079 & ~n4080 ) ;
  assign n4082 = n4078 | n4081 ;
  assign n4083 = n4078 & n4081 ;
  assign n4084 = n4082 & ~n4083 ;
  assign n4085 = ( ~x28 & x29 ) | ( ~x28 & x30 ) | ( x29 & x30 ) ;
  assign n4086 = ( x28 & x29 ) | ( x28 & x30 ) | ( x29 & x30 ) ;
  assign n4087 = ( x28 & n4085 ) | ( x28 & ~n4086 ) | ( n4085 & ~n4086 ) ;
  assign n4088 = ( ~x25 & x26 ) | ( ~x25 & x27 ) | ( x26 & x27 ) ;
  assign n4089 = ( x25 & x26 ) | ( x25 & x27 ) | ( x26 & x27 ) ;
  assign n4090 = ( x25 & n4088 ) | ( x25 & ~n4089 ) | ( n4088 & ~n4089 ) ;
  assign n4091 = ( n4084 & n4087 ) | ( n4084 & n4090 ) | ( n4087 & n4090 ) ;
  assign n4092 = ( ~n4084 & n4087 ) | ( ~n4084 & n4090 ) | ( n4087 & n4090 ) ;
  assign n4093 = ( n4084 & ~n4091 ) | ( n4084 & n4092 ) | ( ~n4091 & n4092 ) ;
  assign n4094 = ( n4057 & n4075 ) | ( n4057 & n4093 ) | ( n4075 & n4093 ) ;
  assign n4095 = ( ~n4057 & n4075 ) | ( ~n4057 & n4093 ) | ( n4075 & n4093 ) ;
  assign n4096 = ( n4057 & ~n4094 ) | ( n4057 & n4095 ) | ( ~n4094 & n4095 ) ;
  assign n4097 = ( ~x58 & x59 ) | ( ~x58 & x60 ) | ( x59 & x60 ) ;
  assign n4098 = ( x58 & x59 ) | ( x58 & x60 ) | ( x59 & x60 ) ;
  assign n4099 = ( x58 & n4097 ) | ( x58 & ~n4098 ) | ( n4097 & ~n4098 ) ;
  assign n4100 = ( ~x55 & x56 ) | ( ~x55 & x57 ) | ( x56 & x57 ) ;
  assign n4101 = ( x55 & x56 ) | ( x55 & x57 ) | ( x56 & x57 ) ;
  assign n4102 = ( x55 & n4100 ) | ( x55 & ~n4101 ) | ( n4100 & ~n4101 ) ;
  assign n4103 = n4099 & n4102 ;
  assign n4104 = n4099 | n4102 ;
  assign n4105 = ~n4103 & n4104 ;
  assign n4106 = ( ~x61 & x62 ) | ( ~x61 & x63 ) | ( x62 & x63 ) ;
  assign n4107 = ( x61 & x62 ) | ( x61 & x63 ) | ( x62 & x63 ) ;
  assign n4108 = ( x61 & n4106 ) | ( x61 & ~n4107 ) | ( n4106 & ~n4107 ) ;
  assign n4109 = ( ~x64 & x65 ) | ( ~x64 & x66 ) | ( x65 & x66 ) ;
  assign n4110 = ( x64 & x65 ) | ( x64 & x66 ) | ( x65 & x66 ) ;
  assign n4111 = ( x64 & n4109 ) | ( x64 & ~n4110 ) | ( n4109 & ~n4110 ) ;
  assign n4112 = ( n4105 & n4108 ) | ( n4105 & n4111 ) | ( n4108 & n4111 ) ;
  assign n4113 = ( ~n4105 & n4108 ) | ( ~n4105 & n4111 ) | ( n4108 & n4111 ) ;
  assign n4114 = ( n4105 & ~n4112 ) | ( n4105 & n4113 ) | ( ~n4112 & n4113 ) ;
  assign n4115 = ( ~x73 & x74 ) | ( ~x73 & x75 ) | ( x74 & x75 ) ;
  assign n4116 = ( x73 & x74 ) | ( x73 & x75 ) | ( x74 & x75 ) ;
  assign n4117 = ( x73 & n4115 ) | ( x73 & ~n4116 ) | ( n4115 & ~n4116 ) ;
  assign n4118 = ( ~x76 & x77 ) | ( ~x76 & x78 ) | ( x77 & x78 ) ;
  assign n4119 = ( x76 & x77 ) | ( x76 & x78 ) | ( x77 & x78 ) ;
  assign n4120 = ( x76 & n4118 ) | ( x76 & ~n4119 ) | ( n4118 & ~n4119 ) ;
  assign n4121 = n4117 & n4120 ;
  assign n4122 = n4117 | n4120 ;
  assign n4123 = ~n4121 & n4122 ;
  assign n4124 = ( ~x70 & x71 ) | ( ~x70 & x72 ) | ( x71 & x72 ) ;
  assign n4125 = ( x70 & x71 ) | ( x70 & x72 ) | ( x71 & x72 ) ;
  assign n4126 = ( x70 & n4124 ) | ( x70 & ~n4125 ) | ( n4124 & ~n4125 ) ;
  assign n4127 = ( ~x67 & x68 ) | ( ~x67 & x69 ) | ( x68 & x69 ) ;
  assign n4128 = ( x67 & x68 ) | ( x67 & x69 ) | ( x68 & x69 ) ;
  assign n4129 = ( x67 & n4127 ) | ( x67 & ~n4128 ) | ( n4127 & ~n4128 ) ;
  assign n4130 = ( n4123 & n4126 ) | ( n4123 & n4129 ) | ( n4126 & n4129 ) ;
  assign n4131 = ( ~n4123 & n4126 ) | ( ~n4123 & n4129 ) | ( n4126 & n4129 ) ;
  assign n4132 = ( n4123 & ~n4130 ) | ( n4123 & n4131 ) | ( ~n4130 & n4131 ) ;
  assign n4133 = n4114 & n4132 ;
  assign n4134 = n4114 | n4132 ;
  assign n4135 = ~n4133 & n4134 ;
  assign n4136 = ( ~x31 & x32 ) | ( ~x31 & x33 ) | ( x32 & x33 ) ;
  assign n4137 = ( x31 & x32 ) | ( x31 & x33 ) | ( x32 & x33 ) ;
  assign n4138 = ( x31 & n4136 ) | ( x31 & ~n4137 ) | ( n4136 & ~n4137 ) ;
  assign n4139 = ( ~x34 & x35 ) | ( ~x34 & x36 ) | ( x35 & x36 ) ;
  assign n4140 = ( x34 & x35 ) | ( x34 & x36 ) | ( x35 & x36 ) ;
  assign n4141 = ( x34 & n4139 ) | ( x34 & ~n4140 ) | ( n4139 & ~n4140 ) ;
  assign n4142 = n4138 & n4141 ;
  assign n4143 = n4138 | n4141 ;
  assign n4144 = ~n4142 & n4143 ;
  assign n4145 = ( ~x37 & x38 ) | ( ~x37 & x39 ) | ( x38 & x39 ) ;
  assign n4146 = ( x37 & x38 ) | ( x37 & x39 ) | ( x38 & x39 ) ;
  assign n4147 = ( x37 & n4145 ) | ( x37 & ~n4146 ) | ( n4145 & ~n4146 ) ;
  assign n4148 = ( ~x40 & x41 ) | ( ~x40 & x42 ) | ( x41 & x42 ) ;
  assign n4149 = ( x40 & x41 ) | ( x40 & x42 ) | ( x41 & x42 ) ;
  assign n4150 = ( x40 & n4148 ) | ( x40 & ~n4149 ) | ( n4148 & ~n4149 ) ;
  assign n4151 = ( n4144 & n4147 ) | ( n4144 & n4150 ) | ( n4147 & n4150 ) ;
  assign n4152 = ( ~n4144 & n4147 ) | ( ~n4144 & n4150 ) | ( n4147 & n4150 ) ;
  assign n4153 = ( n4144 & ~n4151 ) | ( n4144 & n4152 ) | ( ~n4151 & n4152 ) ;
  assign n4154 = ( ~x46 & x47 ) | ( ~x46 & x48 ) | ( x47 & x48 ) ;
  assign n4155 = ( x46 & x47 ) | ( x46 & x48 ) | ( x47 & x48 ) ;
  assign n4156 = ( x46 & n4154 ) | ( x46 & ~n4155 ) | ( n4154 & ~n4155 ) ;
  assign n4157 = ( ~x43 & x44 ) | ( ~x43 & x45 ) | ( x44 & x45 ) ;
  assign n4158 = ( x43 & x44 ) | ( x43 & x45 ) | ( x44 & x45 ) ;
  assign n4159 = ( x43 & n4157 ) | ( x43 & ~n4158 ) | ( n4157 & ~n4158 ) ;
  assign n4160 = n4156 & n4159 ;
  assign n4161 = n4156 | n4159 ;
  assign n4162 = ~n4160 & n4161 ;
  assign n4163 = ( ~x52 & x53 ) | ( ~x52 & x54 ) | ( x53 & x54 ) ;
  assign n4164 = ( x52 & x53 ) | ( x52 & x54 ) | ( x53 & x54 ) ;
  assign n4165 = ( x52 & n4163 ) | ( x52 & ~n4164 ) | ( n4163 & ~n4164 ) ;
  assign n4166 = ( ~x49 & x50 ) | ( ~x49 & x51 ) | ( x50 & x51 ) ;
  assign n4167 = ( x49 & x50 ) | ( x49 & x51 ) | ( x50 & x51 ) ;
  assign n4168 = ( x49 & n4166 ) | ( x49 & ~n4167 ) | ( n4166 & ~n4167 ) ;
  assign n4169 = ( n4162 & n4165 ) | ( n4162 & n4168 ) | ( n4165 & n4168 ) ;
  assign n4170 = ( ~n4162 & n4165 ) | ( ~n4162 & n4168 ) | ( n4165 & n4168 ) ;
  assign n4171 = ( n4162 & ~n4169 ) | ( n4162 & n4170 ) | ( ~n4169 & n4170 ) ;
  assign n4172 = n4153 & n4171 ;
  assign n4173 = n4153 | n4171 ;
  assign n4174 = ~n4172 & n4173 ;
  assign n4175 = n4135 & n4174 ;
  assign n4176 = n4135 | n4174 ;
  assign n4177 = ~n4175 & n4176 ;
  assign n4178 = ( ~x955 & x956 ) | ( ~x955 & x957 ) | ( x956 & x957 ) ;
  assign n4179 = ( x955 & x956 ) | ( x955 & x957 ) | ( x956 & x957 ) ;
  assign n4180 = ( x955 & n4178 ) | ( x955 & ~n4179 ) | ( n4178 & ~n4179 ) ;
  assign n4181 = ( ~x958 & x959 ) | ( ~x958 & x960 ) | ( x959 & x960 ) ;
  assign n4182 = ( x958 & x959 ) | ( x958 & x960 ) | ( x959 & x960 ) ;
  assign n4183 = ( x958 & n4181 ) | ( x958 & ~n4182 ) | ( n4181 & ~n4182 ) ;
  assign n4184 = n4180 | n4183 ;
  assign n4185 = n4180 & n4183 ;
  assign n4186 = n4184 & ~n4185 ;
  assign n4187 = ( ~x964 & x965 ) | ( ~x964 & x966 ) | ( x965 & x966 ) ;
  assign n4188 = ( x964 & x965 ) | ( x964 & x966 ) | ( x965 & x966 ) ;
  assign n4189 = ( x964 & n4187 ) | ( x964 & ~n4188 ) | ( n4187 & ~n4188 ) ;
  assign n4190 = ( ~x961 & x962 ) | ( ~x961 & x963 ) | ( x962 & x963 ) ;
  assign n4191 = ( x961 & x962 ) | ( x961 & x963 ) | ( x962 & x963 ) ;
  assign n4192 = ( x961 & n4190 ) | ( x961 & ~n4191 ) | ( n4190 & ~n4191 ) ;
  assign n4193 = ( n4186 & n4189 ) | ( n4186 & n4192 ) | ( n4189 & n4192 ) ;
  assign n4194 = ( ~n4186 & n4189 ) | ( ~n4186 & n4192 ) | ( n4189 & n4192 ) ;
  assign n4195 = ( n4186 & ~n4193 ) | ( n4186 & n4194 ) | ( ~n4193 & n4194 ) ;
  assign n4196 = ( x949 & x950 ) | ( x949 & x951 ) | ( x950 & x951 ) ;
  assign n4197 = ( ~x949 & x950 ) | ( ~x949 & x951 ) | ( x950 & x951 ) ;
  assign n4198 = ( x949 & ~n4196 ) | ( x949 & n4197 ) | ( ~n4196 & n4197 ) ;
  assign n4199 = ( x952 & x953 ) | ( x952 & x954 ) | ( x953 & x954 ) ;
  assign n4200 = ( ~x952 & x953 ) | ( ~x952 & x954 ) | ( x953 & x954 ) ;
  assign n4201 = ( x952 & ~n4199 ) | ( x952 & n4200 ) | ( ~n4199 & n4200 ) ;
  assign n4202 = n4198 & n4201 ;
  assign n4203 = n4198 | n4201 ;
  assign n4204 = ~n4202 & n4203 ;
  assign n4205 = ( x943 & x944 ) | ( x943 & x945 ) | ( x944 & x945 ) ;
  assign n4206 = ( ~x943 & x944 ) | ( ~x943 & x945 ) | ( x944 & x945 ) ;
  assign n4207 = ( x943 & ~n4205 ) | ( x943 & n4206 ) | ( ~n4205 & n4206 ) ;
  assign n4208 = ( x946 & x947 ) | ( x946 & x948 ) | ( x947 & x948 ) ;
  assign n4209 = ( ~x946 & x947 ) | ( ~x946 & x948 ) | ( x947 & x948 ) ;
  assign n4210 = ( x946 & ~n4208 ) | ( x946 & n4209 ) | ( ~n4208 & n4209 ) ;
  assign n4211 = n4207 & n4210 ;
  assign n4212 = n4207 | n4210 ;
  assign n4213 = ~n4211 & n4212 ;
  assign n4214 = n4204 & n4213 ;
  assign n4215 = n4204 | n4213 ;
  assign n4216 = ~n4214 & n4215 ;
  assign n4217 = n4195 & n4216 ;
  assign n4218 = n4195 | n4216 ;
  assign n4219 = ~n4217 & n4218 ;
  assign n4220 = ( ~x970 & x971 ) | ( ~x970 & x972 ) | ( x971 & x972 ) ;
  assign n4221 = ( x970 & x971 ) | ( x970 & x972 ) | ( x971 & x972 ) ;
  assign n4222 = ( x970 & n4220 ) | ( x970 & ~n4221 ) | ( n4220 & ~n4221 ) ;
  assign n4223 = x967 & x968 ;
  assign n4224 = x967 | x968 ;
  assign n4225 = ~n4223 & n4224 ;
  assign n4226 = ( ~x969 & n4222 ) | ( ~x969 & n4225 ) | ( n4222 & n4225 ) ;
  assign n4227 = ( x969 & n4222 ) | ( x969 & n4225 ) | ( n4222 & n4225 ) ;
  assign n4228 = ( x969 & n4226 ) | ( x969 & ~n4227 ) | ( n4226 & ~n4227 ) ;
  assign n4229 = ( ~x976 & x977 ) | ( ~x976 & x978 ) | ( x977 & x978 ) ;
  assign n4230 = ( x976 & x977 ) | ( x976 & x978 ) | ( x977 & x978 ) ;
  assign n4231 = ( x976 & n4229 ) | ( x976 & ~n4230 ) | ( n4229 & ~n4230 ) ;
  assign n4232 = ( ~x973 & x974 ) | ( ~x973 & x975 ) | ( x974 & x975 ) ;
  assign n4233 = ( x973 & x974 ) | ( x973 & x975 ) | ( x974 & x975 ) ;
  assign n4234 = ( x973 & n4232 ) | ( x973 & ~n4233 ) | ( n4232 & ~n4233 ) ;
  assign n4235 = ( n4228 & n4231 ) | ( n4228 & n4234 ) | ( n4231 & n4234 ) ;
  assign n4236 = ( ~n4228 & n4231 ) | ( ~n4228 & n4234 ) | ( n4231 & n4234 ) ;
  assign n4237 = ( n4228 & ~n4235 ) | ( n4228 & n4236 ) | ( ~n4235 & n4236 ) ;
  assign n4238 = ( ~x982 & x983 ) | ( ~x982 & x984 ) | ( x983 & x984 ) ;
  assign n4239 = ( x982 & x983 ) | ( x982 & x984 ) | ( x983 & x984 ) ;
  assign n4240 = ( x982 & n4238 ) | ( x982 & ~n4239 ) | ( n4238 & ~n4239 ) ;
  assign n4241 = ( ~x979 & x980 ) | ( ~x979 & x981 ) | ( x980 & x981 ) ;
  assign n4242 = ( x979 & x980 ) | ( x979 & x981 ) | ( x980 & x981 ) ;
  assign n4243 = ( x979 & n4241 ) | ( x979 & ~n4242 ) | ( n4241 & ~n4242 ) ;
  assign n4244 = n4240 & n4243 ;
  assign n4245 = n4240 | n4243 ;
  assign n4246 = ~n4244 & n4245 ;
  assign n4247 = ( ~x988 & x989 ) | ( ~x988 & x990 ) | ( x989 & x990 ) ;
  assign n4248 = ( x988 & x989 ) | ( x988 & x990 ) | ( x989 & x990 ) ;
  assign n4249 = ( x988 & n4247 ) | ( x988 & ~n4248 ) | ( n4247 & ~n4248 ) ;
  assign n4250 = ( ~x985 & x986 ) | ( ~x985 & x987 ) | ( x986 & x987 ) ;
  assign n4251 = ( x985 & x986 ) | ( x985 & x987 ) | ( x986 & x987 ) ;
  assign n4252 = ( x985 & n4250 ) | ( x985 & ~n4251 ) | ( n4250 & ~n4251 ) ;
  assign n4253 = ( n4246 & n4249 ) | ( n4246 & n4252 ) | ( n4249 & n4252 ) ;
  assign n4254 = ( ~n4246 & n4249 ) | ( ~n4246 & n4252 ) | ( n4249 & n4252 ) ;
  assign n4255 = ( n4246 & ~n4253 ) | ( n4246 & n4254 ) | ( ~n4253 & n4254 ) ;
  assign n4256 = n4237 & n4255 ;
  assign n4257 = n4237 | n4255 ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4259 = n4219 & n4258 ;
  assign n4260 = n4219 | n4258 ;
  assign n4261 = ~n4259 & n4260 ;
  assign n4262 = ( n4096 & n4177 ) | ( n4096 & n4261 ) | ( n4177 & n4261 ) ;
  assign n4263 = ( ~n4096 & n4177 ) | ( ~n4096 & n4261 ) | ( n4177 & n4261 ) ;
  assign n4264 = ( n4096 & ~n4262 ) | ( n4096 & n4263 ) | ( ~n4262 & n4263 ) ;
  assign n4265 = n4033 & n4264 ;
  assign n4266 = n4033 | n4264 ;
  assign n4267 = ~n4265 & n4266 ;
  assign n4268 = ( n3830 & n3832 ) | ( n3830 & n4267 ) | ( n3832 & n4267 ) ;
  assign n4269 = ~n3833 & n4268 ;
  assign n4270 = ( n3828 & n3833 ) | ( n3828 & n3835 ) | ( n3833 & n3835 ) ;
  assign n4271 = ( ~n3828 & n3833 ) | ( ~n3828 & n3835 ) | ( n3833 & n3835 ) ;
  assign n4272 = ( n3828 & ~n4270 ) | ( n3828 & n4271 ) | ( ~n4270 & n4271 ) ;
  assign n4273 = ( ~n4179 & n4182 ) | ( ~n4179 & n4185 ) | ( n4182 & n4185 ) ;
  assign n4274 = ( n4179 & n4182 ) | ( n4179 & n4185 ) | ( n4182 & n4185 ) ;
  assign n4275 = ( n4179 & n4273 ) | ( n4179 & ~n4274 ) | ( n4273 & ~n4274 ) ;
  assign n4276 = n4193 & n4275 ;
  assign n4277 = n4193 | n4275 ;
  assign n4278 = ~n4276 & n4277 ;
  assign n4279 = ( n4188 & n4191 ) | ( n4188 & n4278 ) | ( n4191 & n4278 ) ;
  assign n4280 = ( n4188 & n4191 ) | ( n4188 & ~n4278 ) | ( n4191 & ~n4278 ) ;
  assign n4281 = ( n4278 & ~n4279 ) | ( n4278 & n4280 ) | ( ~n4279 & n4280 ) ;
  assign n4282 = ( ~n4205 & n4208 ) | ( ~n4205 & n4211 ) | ( n4208 & n4211 ) ;
  assign n4283 = ( n4205 & n4208 ) | ( n4205 & n4211 ) | ( n4208 & n4211 ) ;
  assign n4284 = ( n4205 & n4282 ) | ( n4205 & ~n4283 ) | ( n4282 & ~n4283 ) ;
  assign n4285 = ( n4198 & n4201 ) | ( n4198 & n4213 ) | ( n4201 & n4213 ) ;
  assign n4286 = n4196 & n4199 ;
  assign n4287 = n4196 | n4199 ;
  assign n4288 = ~n4286 & n4287 ;
  assign n4289 = ( n4284 & n4285 ) | ( n4284 & n4288 ) | ( n4285 & n4288 ) ;
  assign n4290 = ( ~n4284 & n4285 ) | ( ~n4284 & n4288 ) | ( n4285 & n4288 ) ;
  assign n4291 = ( n4284 & ~n4289 ) | ( n4284 & n4290 ) | ( ~n4289 & n4290 ) ;
  assign n4292 = ( n4217 & n4281 ) | ( n4217 & n4291 ) | ( n4281 & n4291 ) ;
  assign n4293 = ( n4217 & ~n4281 ) | ( n4217 & n4291 ) | ( ~n4281 & n4291 ) ;
  assign n4294 = ( n4281 & ~n4292 ) | ( n4281 & n4293 ) | ( ~n4292 & n4293 ) ;
  assign n4295 = ( ~n4239 & n4242 ) | ( ~n4239 & n4244 ) | ( n4242 & n4244 ) ;
  assign n4296 = ( n4239 & n4242 ) | ( n4239 & n4244 ) | ( n4242 & n4244 ) ;
  assign n4297 = ( n4239 & n4295 ) | ( n4239 & ~n4296 ) | ( n4295 & ~n4296 ) ;
  assign n4298 = n4248 & n4251 ;
  assign n4299 = n4248 | n4251 ;
  assign n4300 = ~n4298 & n4299 ;
  assign n4301 = ( ~n4253 & n4297 ) | ( ~n4253 & n4300 ) | ( n4297 & n4300 ) ;
  assign n4302 = ( n4253 & n4297 ) | ( n4253 & n4300 ) | ( n4297 & n4300 ) ;
  assign n4303 = ( n4253 & n4301 ) | ( n4253 & ~n4302 ) | ( n4301 & ~n4302 ) ;
  assign n4304 = ( n4221 & n4223 ) | ( n4221 & ~n4227 ) | ( n4223 & ~n4227 ) ;
  assign n4305 = ( n4221 & n4223 ) | ( n4221 & n4227 ) | ( n4223 & n4227 ) ;
  assign n4306 = ( n4227 & n4304 ) | ( n4227 & ~n4305 ) | ( n4304 & ~n4305 ) ;
  assign n4307 = n4230 & n4233 ;
  assign n4308 = n4230 | n4233 ;
  assign n4309 = ~n4307 & n4308 ;
  assign n4310 = ( ~n4235 & n4306 ) | ( ~n4235 & n4309 ) | ( n4306 & n4309 ) ;
  assign n4311 = ( n4235 & n4306 ) | ( n4235 & n4309 ) | ( n4306 & n4309 ) ;
  assign n4312 = ( n4235 & n4310 ) | ( n4235 & ~n4311 ) | ( n4310 & ~n4311 ) ;
  assign n4313 = ( n4256 & n4303 ) | ( n4256 & n4312 ) | ( n4303 & n4312 ) ;
  assign n4314 = ( n4256 & ~n4303 ) | ( n4256 & n4312 ) | ( ~n4303 & n4312 ) ;
  assign n4315 = ( n4303 & ~n4313 ) | ( n4303 & n4314 ) | ( ~n4313 & n4314 ) ;
  assign n4316 = ( n4259 & n4294 ) | ( n4259 & n4315 ) | ( n4294 & n4315 ) ;
  assign n4317 = ( n4259 & ~n4294 ) | ( n4259 & n4315 ) | ( ~n4294 & n4315 ) ;
  assign n4318 = ( n4294 & ~n4316 ) | ( n4294 & n4317 ) | ( ~n4316 & n4317 ) ;
  assign n4319 = ( n4035 & n4038 ) | ( n4035 & ~n4040 ) | ( n4038 & ~n4040 ) ;
  assign n4320 = ( n4035 & n4038 ) | ( n4035 & n4040 ) | ( n4038 & n4040 ) ;
  assign n4321 = ( n4040 & n4319 ) | ( n4040 & ~n4320 ) | ( n4319 & ~n4320 ) ;
  assign n4322 = x999 | n4043 ;
  assign n4323 = ( n4042 & n4044 ) | ( n4042 & n4322 ) | ( n4044 & n4322 ) ;
  assign n4324 = n4321 & n4323 ;
  assign n4325 = x999 & n4043 ;
  assign n4326 = n4042 & n4325 ;
  assign n4327 = n4321 & n4326 ;
  assign n4328 = ( n4321 & n4323 ) | ( n4321 & ~n4326 ) | ( n4323 & ~n4326 ) ;
  assign n4329 = ( ~n4324 & n4327 ) | ( ~n4324 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4330 = n4050 & n4053 ;
  assign n4331 = n4050 | n4053 ;
  assign n4332 = ~n4330 & n4331 ;
  assign n4333 = ( n4055 & n4329 ) | ( n4055 & n4332 ) | ( n4329 & n4332 ) ;
  assign n4334 = ( n4055 & ~n4329 ) | ( n4055 & n4332 ) | ( ~n4329 & n4332 ) ;
  assign n4335 = ( n4329 & ~n4333 ) | ( n4329 & n4334 ) | ( ~n4333 & n4334 ) ;
  assign n4336 = ( ~n4059 & n4062 ) | ( ~n4059 & n4065 ) | ( n4062 & n4065 ) ;
  assign n4337 = ( n4059 & n4062 ) | ( n4059 & n4065 ) | ( n4062 & n4065 ) ;
  assign n4338 = ( n4059 & n4336 ) | ( n4059 & ~n4337 ) | ( n4336 & ~n4337 ) ;
  assign n4339 = n4068 & n4071 ;
  assign n4340 = n4068 | n4071 ;
  assign n4341 = ~n4339 & n4340 ;
  assign n4342 = ( n4073 & n4338 ) | ( n4073 & n4341 ) | ( n4338 & n4341 ) ;
  assign n4343 = ( ~n4073 & n4338 ) | ( ~n4073 & n4341 ) | ( n4338 & n4341 ) ;
  assign n4344 = ( n4073 & ~n4342 ) | ( n4073 & n4343 ) | ( ~n4342 & n4343 ) ;
  assign n4345 = ( ~n4077 & n4080 ) | ( ~n4077 & n4083 ) | ( n4080 & n4083 ) ;
  assign n4346 = ( n4077 & n4080 ) | ( n4077 & n4083 ) | ( n4080 & n4083 ) ;
  assign n4347 = ( n4077 & n4345 ) | ( n4077 & ~n4346 ) | ( n4345 & ~n4346 ) ;
  assign n4348 = n4086 & n4089 ;
  assign n4349 = n4086 | n4089 ;
  assign n4350 = ~n4348 & n4349 ;
  assign n4351 = ( n4091 & n4347 ) | ( n4091 & n4350 ) | ( n4347 & n4350 ) ;
  assign n4352 = ( ~n4091 & n4347 ) | ( ~n4091 & n4350 ) | ( n4347 & n4350 ) ;
  assign n4353 = ( n4091 & ~n4351 ) | ( n4091 & n4352 ) | ( ~n4351 & n4352 ) ;
  assign n4354 = n4344 | n4353 ;
  assign n4355 = n4344 & n4353 ;
  assign n4356 = n4354 & ~n4355 ;
  assign n4357 = ( n4094 & n4335 ) | ( n4094 & n4356 ) | ( n4335 & n4356 ) ;
  assign n4358 = ( ~n4094 & n4335 ) | ( ~n4094 & n4356 ) | ( n4335 & n4356 ) ;
  assign n4359 = ( n4094 & ~n4357 ) | ( n4094 & n4358 ) | ( ~n4357 & n4358 ) ;
  assign n4360 = n4096 & n4177 ;
  assign n4361 = ( ~n4116 & n4119 ) | ( ~n4116 & n4121 ) | ( n4119 & n4121 ) ;
  assign n4362 = ( n4116 & n4119 ) | ( n4116 & n4121 ) | ( n4119 & n4121 ) ;
  assign n4363 = ( n4116 & n4361 ) | ( n4116 & ~n4362 ) | ( n4361 & ~n4362 ) ;
  assign n4364 = n4125 & n4128 ;
  assign n4365 = n4125 | n4128 ;
  assign n4366 = ~n4364 & n4365 ;
  assign n4367 = ( ~n4130 & n4363 ) | ( ~n4130 & n4366 ) | ( n4363 & n4366 ) ;
  assign n4368 = ( n4130 & n4363 ) | ( n4130 & n4366 ) | ( n4363 & n4366 ) ;
  assign n4369 = ( n4130 & n4367 ) | ( n4130 & ~n4368 ) | ( n4367 & ~n4368 ) ;
  assign n4370 = ( ~n4098 & n4101 ) | ( ~n4098 & n4103 ) | ( n4101 & n4103 ) ;
  assign n4371 = ( n4098 & n4101 ) | ( n4098 & n4103 ) | ( n4101 & n4103 ) ;
  assign n4372 = ( n4098 & n4370 ) | ( n4098 & ~n4371 ) | ( n4370 & ~n4371 ) ;
  assign n4373 = n4107 & n4110 ;
  assign n4374 = n4107 | n4110 ;
  assign n4375 = ~n4373 & n4374 ;
  assign n4376 = ( ~n4112 & n4372 ) | ( ~n4112 & n4375 ) | ( n4372 & n4375 ) ;
  assign n4377 = ( n4112 & n4372 ) | ( n4112 & n4375 ) | ( n4372 & n4375 ) ;
  assign n4378 = ( n4112 & n4376 ) | ( n4112 & ~n4377 ) | ( n4376 & ~n4377 ) ;
  assign n4379 = ( n4133 & n4369 ) | ( n4133 & n4378 ) | ( n4369 & n4378 ) ;
  assign n4380 = ( n4133 & ~n4369 ) | ( n4133 & n4378 ) | ( ~n4369 & n4378 ) ;
  assign n4381 = ( n4369 & ~n4379 ) | ( n4369 & n4380 ) | ( ~n4379 & n4380 ) ;
  assign n4382 = ( ~n4155 & n4158 ) | ( ~n4155 & n4160 ) | ( n4158 & n4160 ) ;
  assign n4383 = ( n4155 & n4158 ) | ( n4155 & n4160 ) | ( n4158 & n4160 ) ;
  assign n4384 = ( n4155 & n4382 ) | ( n4155 & ~n4383 ) | ( n4382 & ~n4383 ) ;
  assign n4385 = n4164 & n4167 ;
  assign n4386 = n4164 | n4167 ;
  assign n4387 = ~n4385 & n4386 ;
  assign n4388 = ( n4169 & n4384 ) | ( n4169 & n4387 ) | ( n4384 & n4387 ) ;
  assign n4389 = ( ~n4169 & n4384 ) | ( ~n4169 & n4387 ) | ( n4384 & n4387 ) ;
  assign n4390 = ( n4169 & ~n4388 ) | ( n4169 & n4389 ) | ( ~n4388 & n4389 ) ;
  assign n4391 = ( ~n4137 & n4140 ) | ( ~n4137 & n4142 ) | ( n4140 & n4142 ) ;
  assign n4392 = ( n4137 & n4140 ) | ( n4137 & n4142 ) | ( n4140 & n4142 ) ;
  assign n4393 = ( n4137 & n4391 ) | ( n4137 & ~n4392 ) | ( n4391 & ~n4392 ) ;
  assign n4394 = n4146 & n4149 ;
  assign n4395 = n4146 | n4149 ;
  assign n4396 = ~n4394 & n4395 ;
  assign n4397 = ( ~n4151 & n4393 ) | ( ~n4151 & n4396 ) | ( n4393 & n4396 ) ;
  assign n4398 = ( n4151 & n4393 ) | ( n4151 & n4396 ) | ( n4393 & n4396 ) ;
  assign n4399 = ( n4151 & n4397 ) | ( n4151 & ~n4398 ) | ( n4397 & ~n4398 ) ;
  assign n4400 = ( n4172 & n4390 ) | ( n4172 & n4399 ) | ( n4390 & n4399 ) ;
  assign n4401 = ( n4172 & ~n4390 ) | ( n4172 & n4399 ) | ( ~n4390 & n4399 ) ;
  assign n4402 = ( n4390 & ~n4400 ) | ( n4390 & n4401 ) | ( ~n4400 & n4401 ) ;
  assign n4403 = ( n4175 & n4381 ) | ( n4175 & n4402 ) | ( n4381 & n4402 ) ;
  assign n4404 = ( ~n4175 & n4381 ) | ( ~n4175 & n4402 ) | ( n4381 & n4402 ) ;
  assign n4405 = ( n4175 & ~n4403 ) | ( n4175 & n4404 ) | ( ~n4403 & n4404 ) ;
  assign n4406 = ( n4359 & n4360 ) | ( n4359 & n4405 ) | ( n4360 & n4405 ) ;
  assign n4407 = ( ~n4359 & n4360 ) | ( ~n4359 & n4405 ) | ( n4360 & n4405 ) ;
  assign n4408 = ( n4359 & ~n4406 ) | ( n4359 & n4407 ) | ( ~n4406 & n4407 ) ;
  assign n4409 = n4262 & ~n4360 ;
  assign n4410 = ( n4318 & n4408 ) | ( n4318 & n4409 ) | ( n4408 & n4409 ) ;
  assign n4411 = ( ~n4318 & n4408 ) | ( ~n4318 & n4409 ) | ( n4408 & n4409 ) ;
  assign n4412 = ( n4318 & ~n4410 ) | ( n4318 & n4411 ) | ( ~n4410 & n4411 ) ;
  assign n4413 = n3897 | n3900 ;
  assign n4414 = n3897 & n3900 ;
  assign n4415 = n4413 & ~n4414 ;
  assign n4416 = ( n3895 & n3898 ) | ( n3895 & n3901 ) | ( n3898 & n3901 ) ;
  assign n4417 = ( ~n3888 & n3891 ) | ( ~n3888 & n3894 ) | ( n3891 & n3894 ) ;
  assign n4418 = ( n3888 & n3891 ) | ( n3888 & n3894 ) | ( n3891 & n3894 ) ;
  assign n4419 = ( n3888 & n4417 ) | ( n3888 & ~n4418 ) | ( n4417 & ~n4418 ) ;
  assign n4420 = ( n4415 & n4416 ) | ( n4415 & n4419 ) | ( n4416 & n4419 ) ;
  assign n4421 = ( ~n4415 & n4416 ) | ( ~n4415 & n4419 ) | ( n4416 & n4419 ) ;
  assign n4422 = ( n4415 & ~n4420 ) | ( n4415 & n4421 ) | ( ~n4420 & n4421 ) ;
  assign n4423 = ( ~n3870 & n3873 ) | ( ~n3870 & n3876 ) | ( n3873 & n3876 ) ;
  assign n4424 = ( n3870 & n3873 ) | ( n3870 & n3876 ) | ( n3873 & n3876 ) ;
  assign n4425 = ( n3870 & n4423 ) | ( n3870 & ~n4424 ) | ( n4423 & ~n4424 ) ;
  assign n4426 = ( ~n3879 & n3882 ) | ( ~n3879 & n4425 ) | ( n3882 & n4425 ) ;
  assign n4427 = ( n3879 & n3882 ) | ( n3879 & n4425 ) | ( n3882 & n4425 ) ;
  assign n4428 = ( n3879 & n4426 ) | ( n3879 & ~n4427 ) | ( n4426 & ~n4427 ) ;
  assign n4429 = ( ~n3885 & n4422 ) | ( ~n3885 & n4428 ) | ( n4422 & n4428 ) ;
  assign n4430 = ( n3885 & n4422 ) | ( n3885 & n4428 ) | ( n4422 & n4428 ) ;
  assign n4431 = ( n3885 & n4429 ) | ( n3885 & ~n4430 ) | ( n4429 & ~n4430 ) ;
  assign n4432 = ( ~n3909 & n3912 ) | ( ~n3909 & n3914 ) | ( n3912 & n3914 ) ;
  assign n4433 = ( n3909 & n3912 ) | ( n3909 & n3914 ) | ( n3912 & n3914 ) ;
  assign n4434 = ( n3909 & n4432 ) | ( n3909 & ~n4433 ) | ( n4432 & ~n4433 ) ;
  assign n4435 = n3918 & n3921 ;
  assign n4436 = n3918 | n3921 ;
  assign n4437 = ~n4435 & n4436 ;
  assign n4438 = ( ~n3923 & n4434 ) | ( ~n3923 & n4437 ) | ( n4434 & n4437 ) ;
  assign n4439 = ( n3923 & n4434 ) | ( n3923 & n4437 ) | ( n4434 & n4437 ) ;
  assign n4440 = ( n3923 & n4438 ) | ( n3923 & ~n4439 ) | ( n4438 & ~n4439 ) ;
  assign n4441 = ( ~n3927 & n3930 ) | ( ~n3927 & n3932 ) | ( n3930 & n3932 ) ;
  assign n4442 = ( n3927 & n3930 ) | ( n3927 & n3932 ) | ( n3930 & n3932 ) ;
  assign n4443 = ( n3927 & n4441 ) | ( n3927 & ~n4442 ) | ( n4441 & ~n4442 ) ;
  assign n4444 = n3936 & n3939 ;
  assign n4445 = n3936 | n3939 ;
  assign n4446 = ~n4444 & n4445 ;
  assign n4447 = ( n3941 & n4443 ) | ( n3941 & n4446 ) | ( n4443 & n4446 ) ;
  assign n4448 = ( ~n3941 & n4443 ) | ( ~n3941 & n4446 ) | ( n4443 & n4446 ) ;
  assign n4449 = ( n3941 & ~n4447 ) | ( n3941 & n4448 ) | ( ~n4447 & n4448 ) ;
  assign n4450 = ( n3944 & n4440 ) | ( n3944 & n4449 ) | ( n4440 & n4449 ) ;
  assign n4451 = ( n3944 & ~n4440 ) | ( n3944 & n4449 ) | ( ~n4440 & n4449 ) ;
  assign n4452 = ( n4440 & ~n4450 ) | ( n4440 & n4451 ) | ( ~n4450 & n4451 ) ;
  assign n4453 = ( ~n3947 & n4431 ) | ( ~n3947 & n4452 ) | ( n4431 & n4452 ) ;
  assign n4454 = ( n3947 & n4431 ) | ( n3947 & n4452 ) | ( n4431 & n4452 ) ;
  assign n4455 = ( n3947 & n4453 ) | ( n3947 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = ( ~n3951 & n3954 ) | ( ~n3951 & n3956 ) | ( n3954 & n3956 ) ;
  assign n4457 = ( n3951 & n3954 ) | ( n3951 & n3956 ) | ( n3954 & n3956 ) ;
  assign n4458 = ( n3951 & n4456 ) | ( n3951 & ~n4457 ) | ( n4456 & ~n4457 ) ;
  assign n4459 = n3960 & n3963 ;
  assign n4460 = n3960 | n3963 ;
  assign n4461 = ~n4459 & n4460 ;
  assign n4462 = ( ~n3965 & n4458 ) | ( ~n3965 & n4461 ) | ( n4458 & n4461 ) ;
  assign n4463 = ( n3965 & n4458 ) | ( n3965 & n4461 ) | ( n4458 & n4461 ) ;
  assign n4464 = ( n3965 & n4462 ) | ( n3965 & ~n4463 ) | ( n4462 & ~n4463 ) ;
  assign n4465 = ( ~n3969 & n3972 ) | ( ~n3969 & n3974 ) | ( n3972 & n3974 ) ;
  assign n4466 = ( n3969 & n3972 ) | ( n3969 & n3974 ) | ( n3972 & n3974 ) ;
  assign n4467 = ( n3969 & n4465 ) | ( n3969 & ~n4466 ) | ( n4465 & ~n4466 ) ;
  assign n4468 = n3978 & n3981 ;
  assign n4469 = n3978 | n3981 ;
  assign n4470 = ~n4468 & n4469 ;
  assign n4471 = ( n3983 & n4467 ) | ( n3983 & n4470 ) | ( n4467 & n4470 ) ;
  assign n4472 = ( ~n3983 & n4467 ) | ( ~n3983 & n4470 ) | ( n4467 & n4470 ) ;
  assign n4473 = ( n3983 & ~n4471 ) | ( n3983 & n4472 ) | ( ~n4471 & n4472 ) ;
  assign n4474 = ( n3986 & n4464 ) | ( n3986 & n4473 ) | ( n4464 & n4473 ) ;
  assign n4475 = ( ~n3986 & n4464 ) | ( ~n3986 & n4473 ) | ( n4464 & n4473 ) ;
  assign n4476 = ( n3986 & ~n4474 ) | ( n3986 & n4475 ) | ( ~n4474 & n4475 ) ;
  assign n4477 = ( ~n3990 & n3993 ) | ( ~n3990 & n3995 ) | ( n3993 & n3995 ) ;
  assign n4478 = ( n3990 & n3993 ) | ( n3990 & n3995 ) | ( n3993 & n3995 ) ;
  assign n4479 = ( n3990 & n4477 ) | ( n3990 & ~n4478 ) | ( n4477 & ~n4478 ) ;
  assign n4480 = n3999 & n4002 ;
  assign n4481 = n3999 | n4002 ;
  assign n4482 = ~n4480 & n4481 ;
  assign n4483 = ( ~n4004 & n4479 ) | ( ~n4004 & n4482 ) | ( n4479 & n4482 ) ;
  assign n4484 = ( n4004 & n4479 ) | ( n4004 & n4482 ) | ( n4479 & n4482 ) ;
  assign n4485 = ( n4004 & n4483 ) | ( n4004 & ~n4484 ) | ( n4483 & ~n4484 ) ;
  assign n4486 = ( ~n4008 & n4011 ) | ( ~n4008 & n4013 ) | ( n4011 & n4013 ) ;
  assign n4487 = ( n4008 & n4011 ) | ( n4008 & n4013 ) | ( n4011 & n4013 ) ;
  assign n4488 = ( n4008 & n4486 ) | ( n4008 & ~n4487 ) | ( n4486 & ~n4487 ) ;
  assign n4489 = n4017 & n4020 ;
  assign n4490 = n4017 | n4020 ;
  assign n4491 = ~n4489 & n4490 ;
  assign n4492 = ( n4022 & n4488 ) | ( n4022 & n4491 ) | ( n4488 & n4491 ) ;
  assign n4493 = ( ~n4022 & n4488 ) | ( ~n4022 & n4491 ) | ( n4488 & n4491 ) ;
  assign n4494 = ( n4022 & ~n4492 ) | ( n4022 & n4493 ) | ( ~n4492 & n4493 ) ;
  assign n4495 = ( n4025 & n4485 ) | ( n4025 & n4494 ) | ( n4485 & n4494 ) ;
  assign n4496 = ( n4025 & ~n4485 ) | ( n4025 & n4494 ) | ( ~n4485 & n4494 ) ;
  assign n4497 = ( n4485 & ~n4495 ) | ( n4485 & n4496 ) | ( ~n4495 & n4496 ) ;
  assign n4498 = ( n4028 & n4476 ) | ( n4028 & n4497 ) | ( n4476 & n4497 ) ;
  assign n4499 = ( ~n4028 & n4476 ) | ( ~n4028 & n4497 ) | ( n4476 & n4497 ) ;
  assign n4500 = ( n4028 & ~n4498 ) | ( n4028 & n4499 ) | ( ~n4498 & n4499 ) ;
  assign n4501 = ( n4031 & n4455 ) | ( n4031 & n4500 ) | ( n4455 & n4500 ) ;
  assign n4502 = ( ~n4031 & n4455 ) | ( ~n4031 & n4500 ) | ( n4455 & n4500 ) ;
  assign n4503 = ( n4031 & ~n4501 ) | ( n4031 & n4502 ) | ( ~n4501 & n4502 ) ;
  assign n4504 = ( n4265 & n4412 ) | ( n4265 & n4503 ) | ( n4412 & n4503 ) ;
  assign n4505 = ( n4265 & ~n4412 ) | ( n4265 & n4503 ) | ( ~n4412 & n4503 ) ;
  assign n4506 = ( n4412 & ~n4504 ) | ( n4412 & n4505 ) | ( ~n4504 & n4505 ) ;
  assign n4507 = ( n4269 & n4272 ) | ( n4269 & n4506 ) | ( n4272 & n4506 ) ;
  assign n4508 = ( ~n3840 & n3842 ) | ( ~n3840 & n3844 ) | ( n3842 & n3844 ) ;
  assign n4509 = ( n3840 & ~n3845 ) | ( n3840 & n4508 ) | ( ~n3845 & n4508 ) ;
  assign n4510 = ( ~n4305 & n4307 ) | ( ~n4305 & n4311 ) | ( n4307 & n4311 ) ;
  assign n4511 = ( n4305 & n4307 ) | ( n4305 & n4311 ) | ( n4307 & n4311 ) ;
  assign n4512 = ( n4305 & n4510 ) | ( n4305 & ~n4511 ) | ( n4510 & ~n4511 ) ;
  assign n4513 = ( n4296 & n4298 ) | ( n4296 & ~n4302 ) | ( n4298 & ~n4302 ) ;
  assign n4514 = ( n4296 & n4298 ) | ( n4296 & n4302 ) | ( n4298 & n4302 ) ;
  assign n4515 = ( n4302 & n4513 ) | ( n4302 & ~n4514 ) | ( n4513 & ~n4514 ) ;
  assign n4516 = ( ~n4313 & n4512 ) | ( ~n4313 & n4515 ) | ( n4512 & n4515 ) ;
  assign n4517 = ( n4313 & n4512 ) | ( n4313 & n4515 ) | ( n4512 & n4515 ) ;
  assign n4518 = ( n4313 & n4516 ) | ( n4313 & ~n4517 ) | ( n4516 & ~n4517 ) ;
  assign n4519 = ( n4274 & n4276 ) | ( n4274 & n4279 ) | ( n4276 & n4279 ) ;
  assign n4520 = ( n4274 & n4276 ) | ( n4274 & ~n4279 ) | ( n4276 & ~n4279 ) ;
  assign n4521 = ( n4279 & ~n4519 ) | ( n4279 & n4520 ) | ( ~n4519 & n4520 ) ;
  assign n4522 = ( n4214 & n4289 ) | ( n4214 & ~n4290 ) | ( n4289 & ~n4290 ) ;
  assign n4523 = ( n4196 & n4199 ) | ( n4196 & n4202 ) | ( n4199 & n4202 ) ;
  assign n4524 = ( n4283 & n4522 ) | ( n4283 & n4523 ) | ( n4522 & n4523 ) ;
  assign n4525 = ( n4283 & ~n4522 ) | ( n4283 & n4523 ) | ( ~n4522 & n4523 ) ;
  assign n4526 = ( n4522 & ~n4524 ) | ( n4522 & n4525 ) | ( ~n4524 & n4525 ) ;
  assign n4527 = ( n4292 & n4521 ) | ( n4292 & n4526 ) | ( n4521 & n4526 ) ;
  assign n4528 = ( ~n4292 & n4521 ) | ( ~n4292 & n4526 ) | ( n4521 & n4526 ) ;
  assign n4529 = ( n4292 & ~n4527 ) | ( n4292 & n4528 ) | ( ~n4527 & n4528 ) ;
  assign n4530 = ( ~n4316 & n4518 ) | ( ~n4316 & n4529 ) | ( n4518 & n4529 ) ;
  assign n4531 = ( n4316 & n4518 ) | ( n4316 & n4529 ) | ( n4518 & n4529 ) ;
  assign n4532 = ( n4316 & n4530 ) | ( n4316 & ~n4531 ) | ( n4530 & ~n4531 ) ;
  assign n4533 = n4324 | n4326 ;
  assign n4534 = n4320 & n4330 ;
  assign n4535 = n4320 | n4330 ;
  assign n4536 = ~n4534 & n4535 ;
  assign n4537 = ( n4333 & n4533 ) | ( n4333 & n4536 ) | ( n4533 & n4536 ) ;
  assign n4538 = ( ~n4333 & n4533 ) | ( ~n4333 & n4536 ) | ( n4533 & n4536 ) ;
  assign n4539 = ( n4333 & ~n4537 ) | ( n4333 & n4538 ) | ( ~n4537 & n4538 ) ;
  assign n4540 = n4075 & n4093 ;
  assign n4541 = n4356 & ~n4540 ;
  assign n4542 = ( n4335 & ~n4358 ) | ( n4335 & n4541 ) | ( ~n4358 & n4541 ) ;
  assign n4543 = ( n4346 & n4348 ) | ( n4346 & ~n4351 ) | ( n4348 & ~n4351 ) ;
  assign n4544 = ( n4346 & n4348 ) | ( n4346 & n4351 ) | ( n4348 & n4351 ) ;
  assign n4545 = ( n4351 & n4543 ) | ( n4351 & ~n4544 ) | ( n4543 & ~n4544 ) ;
  assign n4546 = ( n4344 & n4353 ) | ( n4344 & n4540 ) | ( n4353 & n4540 ) ;
  assign n4547 = ( n4337 & n4339 ) | ( n4337 & n4342 ) | ( n4339 & n4342 ) ;
  assign n4548 = ( n4337 & n4339 ) | ( n4337 & ~n4342 ) | ( n4339 & ~n4342 ) ;
  assign n4549 = ( n4342 & ~n4547 ) | ( n4342 & n4548 ) | ( ~n4547 & n4548 ) ;
  assign n4550 = ( ~n4545 & n4546 ) | ( ~n4545 & n4549 ) | ( n4546 & n4549 ) ;
  assign n4551 = ( n4545 & n4546 ) | ( n4545 & n4549 ) | ( n4546 & n4549 ) ;
  assign n4552 = ( n4545 & n4550 ) | ( n4545 & ~n4551 ) | ( n4550 & ~n4551 ) ;
  assign n4553 = ( ~n4539 & n4542 ) | ( ~n4539 & n4552 ) | ( n4542 & n4552 ) ;
  assign n4554 = ( n4539 & n4542 ) | ( n4539 & n4552 ) | ( n4542 & n4552 ) ;
  assign n4555 = ( n4539 & n4553 ) | ( n4539 & ~n4554 ) | ( n4553 & ~n4554 ) ;
  assign n4556 = ( n4371 & n4373 ) | ( n4371 & n4377 ) | ( n4373 & n4377 ) ;
  assign n4557 = ( n4371 & n4373 ) | ( n4371 & ~n4377 ) | ( n4373 & ~n4377 ) ;
  assign n4558 = ( n4377 & ~n4556 ) | ( n4377 & n4557 ) | ( ~n4556 & n4557 ) ;
  assign n4559 = ( n4362 & n4364 ) | ( n4362 & ~n4368 ) | ( n4364 & ~n4368 ) ;
  assign n4560 = ( n4362 & n4364 ) | ( n4362 & n4368 ) | ( n4364 & n4368 ) ;
  assign n4561 = ( n4368 & n4559 ) | ( n4368 & ~n4560 ) | ( n4559 & ~n4560 ) ;
  assign n4562 = ( ~n4379 & n4558 ) | ( ~n4379 & n4561 ) | ( n4558 & n4561 ) ;
  assign n4563 = ( n4379 & n4558 ) | ( n4379 & n4561 ) | ( n4558 & n4561 ) ;
  assign n4564 = ( n4379 & n4562 ) | ( n4379 & ~n4563 ) | ( n4562 & ~n4563 ) ;
  assign n4565 = ( n4383 & n4385 ) | ( n4383 & ~n4388 ) | ( n4385 & ~n4388 ) ;
  assign n4566 = ( n4383 & n4385 ) | ( n4383 & n4388 ) | ( n4385 & n4388 ) ;
  assign n4567 = ( n4388 & n4565 ) | ( n4388 & ~n4566 ) | ( n4565 & ~n4566 ) ;
  assign n4568 = ( n4392 & n4394 ) | ( n4392 & n4398 ) | ( n4394 & n4398 ) ;
  assign n4569 = ( n4392 & n4394 ) | ( n4392 & ~n4398 ) | ( n4394 & ~n4398 ) ;
  assign n4570 = ( n4398 & ~n4568 ) | ( n4398 & n4569 ) | ( ~n4568 & n4569 ) ;
  assign n4571 = ( n4400 & n4567 ) | ( n4400 & n4570 ) | ( n4567 & n4570 ) ;
  assign n4572 = ( ~n4400 & n4567 ) | ( ~n4400 & n4570 ) | ( n4567 & n4570 ) ;
  assign n4573 = ( n4400 & ~n4571 ) | ( n4400 & n4572 ) | ( ~n4571 & n4572 ) ;
  assign n4574 = ( ~n4403 & n4564 ) | ( ~n4403 & n4573 ) | ( n4564 & n4573 ) ;
  assign n4575 = ( n4403 & n4564 ) | ( n4403 & n4573 ) | ( n4564 & n4573 ) ;
  assign n4576 = ( n4403 & n4574 ) | ( n4403 & ~n4575 ) | ( n4574 & ~n4575 ) ;
  assign n4577 = ( n4406 & n4555 ) | ( n4406 & n4576 ) | ( n4555 & n4576 ) ;
  assign n4578 = ( n4406 & ~n4555 ) | ( n4406 & n4576 ) | ( ~n4555 & n4576 ) ;
  assign n4579 = ( n4555 & ~n4577 ) | ( n4555 & n4578 ) | ( ~n4577 & n4578 ) ;
  assign n4580 = ( n4410 & n4532 ) | ( n4410 & n4579 ) | ( n4532 & n4579 ) ;
  assign n4581 = ( ~n4410 & n4532 ) | ( ~n4410 & n4579 ) | ( n4532 & n4579 ) ;
  assign n4582 = ( n4410 & ~n4580 ) | ( n4410 & n4581 ) | ( ~n4580 & n4581 ) ;
  assign n4583 = ( n4442 & n4444 ) | ( n4442 & n4447 ) | ( n4444 & n4447 ) ;
  assign n4584 = ( n4442 & n4444 ) | ( n4442 & ~n4447 ) | ( n4444 & ~n4447 ) ;
  assign n4585 = ( n4447 & ~n4583 ) | ( n4447 & n4584 ) | ( ~n4583 & n4584 ) ;
  assign n4586 = ( n4433 & n4435 ) | ( n4433 & n4439 ) | ( n4435 & n4439 ) ;
  assign n4587 = ( n4433 & n4435 ) | ( n4433 & ~n4439 ) | ( n4435 & ~n4439 ) ;
  assign n4588 = ( n4439 & ~n4586 ) | ( n4439 & n4587 ) | ( ~n4586 & n4587 ) ;
  assign n4589 = ( n4450 & n4585 ) | ( n4450 & n4588 ) | ( n4585 & n4588 ) ;
  assign n4590 = ( ~n4450 & n4585 ) | ( ~n4450 & n4588 ) | ( n4585 & n4588 ) ;
  assign n4591 = ( n4450 & ~n4589 ) | ( n4450 & n4590 ) | ( ~n4589 & n4590 ) ;
  assign n4592 = n3886 & n3907 ;
  assign n4593 = n4431 & ~n4592 ;
  assign n4594 = ( ~n4431 & n4454 ) | ( ~n4431 & n4593 ) | ( n4454 & n4593 ) ;
  assign n4595 = ( n3906 & n4419 ) | ( n3906 & ~n4422 ) | ( n4419 & ~n4422 ) ;
  assign n4596 = ( n3897 & n3900 ) | ( n3897 & n3902 ) | ( n3900 & n3902 ) ;
  assign n4597 = ( n4418 & n4595 ) | ( n4418 & n4596 ) | ( n4595 & n4596 ) ;
  assign n4598 = ( ~n4418 & n4595 ) | ( ~n4418 & n4596 ) | ( n4595 & n4596 ) ;
  assign n4599 = ( n4418 & ~n4597 ) | ( n4418 & n4598 ) | ( ~n4597 & n4598 ) ;
  assign n4600 = ~n3885 & n4428 ;
  assign n4601 = n3879 | n4426 ;
  assign n4602 = n3879 & n4426 ;
  assign n4603 = n4601 & ~n4602 ;
  assign n4604 = ( n4424 & n4600 ) | ( n4424 & n4603 ) | ( n4600 & n4603 ) ;
  assign n4605 = ( ~n4424 & n4600 ) | ( ~n4424 & n4603 ) | ( n4600 & n4603 ) ;
  assign n4606 = ( n4424 & ~n4604 ) | ( n4424 & n4605 ) | ( ~n4604 & n4605 ) ;
  assign n4607 = ( n4431 & n4592 ) | ( n4431 & n4600 ) | ( n4592 & n4600 ) ;
  assign n4608 = ( n4422 & ~n4593 ) | ( n4422 & n4607 ) | ( ~n4593 & n4607 ) ;
  assign n4609 = ( n4599 & n4606 ) | ( n4599 & n4608 ) | ( n4606 & n4608 ) ;
  assign n4610 = ( ~n4599 & n4606 ) | ( ~n4599 & n4608 ) | ( n4606 & n4608 ) ;
  assign n4611 = ( n4599 & ~n4609 ) | ( n4599 & n4610 ) | ( ~n4609 & n4610 ) ;
  assign n4612 = ( n4591 & n4594 ) | ( n4591 & n4611 ) | ( n4594 & n4611 ) ;
  assign n4613 = ( ~n4591 & n4594 ) | ( ~n4591 & n4611 ) | ( n4594 & n4611 ) ;
  assign n4614 = ( n4591 & ~n4612 ) | ( n4591 & n4613 ) | ( ~n4612 & n4613 ) ;
  assign n4615 = ( n4466 & n4468 ) | ( n4466 & ~n4471 ) | ( n4468 & ~n4471 ) ;
  assign n4616 = ( n4466 & n4468 ) | ( n4466 & n4471 ) | ( n4468 & n4471 ) ;
  assign n4617 = ( n4471 & n4615 ) | ( n4471 & ~n4616 ) | ( n4615 & ~n4616 ) ;
  assign n4618 = ( n4457 & n4459 ) | ( n4457 & ~n4463 ) | ( n4459 & ~n4463 ) ;
  assign n4619 = ( n4457 & n4459 ) | ( n4457 & n4463 ) | ( n4459 & n4463 ) ;
  assign n4620 = ( n4463 & n4618 ) | ( n4463 & ~n4619 ) | ( n4618 & ~n4619 ) ;
  assign n4621 = ( ~n4474 & n4617 ) | ( ~n4474 & n4620 ) | ( n4617 & n4620 ) ;
  assign n4622 = ( n4474 & n4617 ) | ( n4474 & n4620 ) | ( n4617 & n4620 ) ;
  assign n4623 = ( n4474 & n4621 ) | ( n4474 & ~n4622 ) | ( n4621 & ~n4622 ) ;
  assign n4624 = ( n4487 & n4489 ) | ( n4487 & n4492 ) | ( n4489 & n4492 ) ;
  assign n4625 = ( n4487 & n4489 ) | ( n4487 & ~n4492 ) | ( n4489 & ~n4492 ) ;
  assign n4626 = ( n4492 & ~n4624 ) | ( n4492 & n4625 ) | ( ~n4624 & n4625 ) ;
  assign n4627 = ( n4478 & n4480 ) | ( n4478 & n4484 ) | ( n4480 & n4484 ) ;
  assign n4628 = ( n4478 & n4480 ) | ( n4478 & ~n4484 ) | ( n4480 & ~n4484 ) ;
  assign n4629 = ( n4484 & ~n4627 ) | ( n4484 & n4628 ) | ( ~n4627 & n4628 ) ;
  assign n4630 = ( n4495 & n4626 ) | ( n4495 & n4629 ) | ( n4626 & n4629 ) ;
  assign n4631 = ( ~n4495 & n4626 ) | ( ~n4495 & n4629 ) | ( n4626 & n4629 ) ;
  assign n4632 = ( n4495 & ~n4630 ) | ( n4495 & n4631 ) | ( ~n4630 & n4631 ) ;
  assign n4633 = ( n4498 & n4623 ) | ( n4498 & n4632 ) | ( n4623 & n4632 ) ;
  assign n4634 = ( n4498 & ~n4623 ) | ( n4498 & n4632 ) | ( ~n4623 & n4632 ) ;
  assign n4635 = ( n4623 & ~n4633 ) | ( n4623 & n4634 ) | ( ~n4633 & n4634 ) ;
  assign n4636 = ( ~n4501 & n4614 ) | ( ~n4501 & n4635 ) | ( n4614 & n4635 ) ;
  assign n4637 = ( n4501 & n4614 ) | ( n4501 & n4635 ) | ( n4614 & n4635 ) ;
  assign n4638 = ( n4501 & n4636 ) | ( n4501 & ~n4637 ) | ( n4636 & ~n4637 ) ;
  assign n4639 = ( n4504 & n4582 ) | ( n4504 & n4638 ) | ( n4582 & n4638 ) ;
  assign n4640 = ( n4504 & ~n4582 ) | ( n4504 & n4638 ) | ( ~n4582 & n4638 ) ;
  assign n4641 = ( n4582 & ~n4639 ) | ( n4582 & n4640 ) | ( ~n4639 & n4640 ) ;
  assign n4642 = ( n4507 & n4509 ) | ( n4507 & n4641 ) | ( n4509 & n4641 ) ;
  assign n4643 = ( ~n3845 & n3847 ) | ( ~n3845 & n3849 ) | ( n3847 & n3849 ) ;
  assign n4644 = ( n3845 & ~n3850 ) | ( n3845 & n4643 ) | ( ~n3850 & n4643 ) ;
  assign n4645 = ( n4519 & n4524 ) | ( n4519 & ~n4527 ) | ( n4524 & ~n4527 ) ;
  assign n4646 = ( n4519 & n4524 ) | ( n4519 & n4527 ) | ( n4524 & n4527 ) ;
  assign n4647 = ( n4527 & n4645 ) | ( n4527 & ~n4646 ) | ( n4645 & ~n4646 ) ;
  assign n4648 = ( n4511 & n4514 ) | ( n4511 & n4517 ) | ( n4514 & n4517 ) ;
  assign n4649 = ( n4511 & n4514 ) | ( n4511 & ~n4517 ) | ( n4514 & ~n4517 ) ;
  assign n4650 = ( n4517 & ~n4648 ) | ( n4517 & n4649 ) | ( ~n4648 & n4649 ) ;
  assign n4651 = ( ~n4531 & n4647 ) | ( ~n4531 & n4650 ) | ( n4647 & n4650 ) ;
  assign n4652 = ( n4531 & n4647 ) | ( n4531 & n4650 ) | ( n4647 & n4650 ) ;
  assign n4653 = ( n4531 & n4651 ) | ( n4531 & ~n4652 ) | ( n4651 & ~n4652 ) ;
  assign n4654 = ( n4544 & n4547 ) | ( n4544 & n4551 ) | ( n4547 & n4551 ) ;
  assign n4655 = ( n4544 & n4547 ) | ( n4544 & ~n4551 ) | ( n4547 & ~n4551 ) ;
  assign n4656 = ( n4551 & ~n4654 ) | ( n4551 & n4655 ) | ( ~n4654 & n4655 ) ;
  assign n4657 = n4534 & ~n4537 ;
  assign n4658 = ~n4534 & n4537 ;
  assign n4659 = n4657 | n4658 ;
  assign n4660 = ( ~n4554 & n4656 ) | ( ~n4554 & n4659 ) | ( n4656 & n4659 ) ;
  assign n4661 = ( n4554 & n4656 ) | ( n4554 & n4659 ) | ( n4656 & n4659 ) ;
  assign n4662 = ( n4554 & n4660 ) | ( n4554 & ~n4661 ) | ( n4660 & ~n4661 ) ;
  assign n4663 = ( ~n4566 & n4568 ) | ( ~n4566 & n4571 ) | ( n4568 & n4571 ) ;
  assign n4664 = ( n4566 & n4568 ) | ( n4566 & n4571 ) | ( n4568 & n4571 ) ;
  assign n4665 = ( n4566 & n4663 ) | ( n4566 & ~n4664 ) | ( n4663 & ~n4664 ) ;
  assign n4666 = ( n4556 & n4560 ) | ( n4556 & ~n4563 ) | ( n4560 & ~n4563 ) ;
  assign n4667 = ( n4556 & n4560 ) | ( n4556 & n4563 ) | ( n4560 & n4563 ) ;
  assign n4668 = ( n4563 & n4666 ) | ( n4563 & ~n4667 ) | ( n4666 & ~n4667 ) ;
  assign n4669 = ( ~n4575 & n4665 ) | ( ~n4575 & n4668 ) | ( n4665 & n4668 ) ;
  assign n4670 = ( n4575 & n4665 ) | ( n4575 & n4668 ) | ( n4665 & n4668 ) ;
  assign n4671 = ( n4575 & n4669 ) | ( n4575 & ~n4670 ) | ( n4669 & ~n4670 ) ;
  assign n4672 = ( n4577 & n4662 ) | ( n4577 & n4671 ) | ( n4662 & n4671 ) ;
  assign n4673 = ( ~n4577 & n4662 ) | ( ~n4577 & n4671 ) | ( n4662 & n4671 ) ;
  assign n4674 = ( n4577 & ~n4672 ) | ( n4577 & n4673 ) | ( ~n4672 & n4673 ) ;
  assign n4675 = ( n4580 & n4653 ) | ( n4580 & n4674 ) | ( n4653 & n4674 ) ;
  assign n4676 = ( ~n4580 & n4653 ) | ( ~n4580 & n4674 ) | ( n4653 & n4674 ) ;
  assign n4677 = ( n4580 & ~n4675 ) | ( n4580 & n4676 ) | ( ~n4675 & n4676 ) ;
  assign n4678 = ( ~n4624 & n4627 ) | ( ~n4624 & n4630 ) | ( n4627 & n4630 ) ;
  assign n4679 = ( n4624 & n4627 ) | ( n4624 & n4630 ) | ( n4627 & n4630 ) ;
  assign n4680 = ( n4624 & n4678 ) | ( n4624 & ~n4679 ) | ( n4678 & ~n4679 ) ;
  assign n4681 = ( n4616 & n4619 ) | ( n4616 & n4622 ) | ( n4619 & n4622 ) ;
  assign n4682 = ( n4616 & n4619 ) | ( n4616 & ~n4622 ) | ( n4619 & ~n4622 ) ;
  assign n4683 = ( n4622 & ~n4681 ) | ( n4622 & n4682 ) | ( ~n4681 & n4682 ) ;
  assign n4684 = ( n4633 & n4680 ) | ( n4633 & n4683 ) | ( n4680 & n4683 ) ;
  assign n4685 = ( n4633 & ~n4680 ) | ( n4633 & n4683 ) | ( ~n4680 & n4683 ) ;
  assign n4686 = ( n4680 & ~n4684 ) | ( n4680 & n4685 ) | ( ~n4684 & n4685 ) ;
  assign n4687 = n3879 & n3882 ;
  assign n4688 = ( n4604 & ~n4605 ) | ( n4604 & n4687 ) | ( ~n4605 & n4687 ) ;
  assign n4689 = ( n4597 & n4609 ) | ( n4597 & n4688 ) | ( n4609 & n4688 ) ;
  assign n4690 = ( ~n4597 & n4609 ) | ( ~n4597 & n4688 ) | ( n4609 & n4688 ) ;
  assign n4691 = ( n4597 & ~n4689 ) | ( n4597 & n4690 ) | ( ~n4689 & n4690 ) ;
  assign n4692 = ( n4583 & n4586 ) | ( n4583 & ~n4589 ) | ( n4586 & ~n4589 ) ;
  assign n4693 = ( n4583 & n4586 ) | ( n4583 & n4589 ) | ( n4586 & n4589 ) ;
  assign n4694 = ( n4589 & n4692 ) | ( n4589 & ~n4693 ) | ( n4692 & ~n4693 ) ;
  assign n4695 = ( n4612 & n4691 ) | ( n4612 & n4694 ) | ( n4691 & n4694 ) ;
  assign n4696 = ( ~n4612 & n4691 ) | ( ~n4612 & n4694 ) | ( n4691 & n4694 ) ;
  assign n4697 = ( n4612 & ~n4695 ) | ( n4612 & n4696 ) | ( ~n4695 & n4696 ) ;
  assign n4698 = ( n4637 & n4686 ) | ( n4637 & n4697 ) | ( n4686 & n4697 ) ;
  assign n4699 = ( n4637 & ~n4686 ) | ( n4637 & n4697 ) | ( ~n4686 & n4697 ) ;
  assign n4700 = ( n4686 & ~n4698 ) | ( n4686 & n4699 ) | ( ~n4698 & n4699 ) ;
  assign n4701 = ( n4639 & n4677 ) | ( n4639 & n4700 ) | ( n4677 & n4700 ) ;
  assign n4702 = ( n4639 & ~n4677 ) | ( n4639 & n4700 ) | ( ~n4677 & n4700 ) ;
  assign n4703 = ( n4677 & ~n4701 ) | ( n4677 & n4702 ) | ( ~n4701 & n4702 ) ;
  assign n4704 = ( n4642 & n4644 ) | ( n4642 & n4703 ) | ( n4644 & n4703 ) ;
  assign n4705 = ( n4689 & n4693 ) | ( n4689 & ~n4695 ) | ( n4693 & ~n4695 ) ;
  assign n4706 = ( n4689 & n4693 ) | ( n4689 & n4695 ) | ( n4693 & n4695 ) ;
  assign n4707 = ( n4695 & n4705 ) | ( n4695 & ~n4706 ) | ( n4705 & ~n4706 ) ;
  assign n4708 = ( n4679 & n4681 ) | ( n4679 & n4684 ) | ( n4681 & n4684 ) ;
  assign n4709 = ( ~n4679 & n4681 ) | ( ~n4679 & n4684 ) | ( n4681 & n4684 ) ;
  assign n4710 = ( n4679 & ~n4708 ) | ( n4679 & n4709 ) | ( ~n4708 & n4709 ) ;
  assign n4711 = ( ~n4698 & n4707 ) | ( ~n4698 & n4710 ) | ( n4707 & n4710 ) ;
  assign n4712 = ( n4698 & n4707 ) | ( n4698 & n4710 ) | ( n4707 & n4710 ) ;
  assign n4713 = ( n4698 & n4711 ) | ( n4698 & ~n4712 ) | ( n4711 & ~n4712 ) ;
  assign n4714 = ( n4646 & n4648 ) | ( n4646 & n4652 ) | ( n4648 & n4652 ) ;
  assign n4715 = ( n4646 & n4648 ) | ( n4646 & ~n4652 ) | ( n4648 & ~n4652 ) ;
  assign n4716 = ( n4652 & ~n4714 ) | ( n4652 & n4715 ) | ( ~n4714 & n4715 ) ;
  assign n4717 = ( n4664 & n4667 ) | ( n4664 & n4670 ) | ( n4667 & n4670 ) ;
  assign n4718 = ( n4664 & n4667 ) | ( n4664 & ~n4670 ) | ( n4667 & ~n4670 ) ;
  assign n4719 = ( n4670 & ~n4717 ) | ( n4670 & n4718 ) | ( ~n4717 & n4718 ) ;
  assign n4720 = n4672 & n4719 ;
  assign n4721 = n4672 | n4719 ;
  assign n4722 = ~n4720 & n4721 ;
  assign n4723 = n4333 & n4533 ;
  assign n4724 = ~n4534 & n4723 ;
  assign n4725 = ( n4661 & n4723 ) | ( n4661 & ~n4724 ) | ( n4723 & ~n4724 ) ;
  assign n4726 = ( n4654 & n4722 ) | ( n4654 & n4725 ) | ( n4722 & n4725 ) ;
  assign n4727 = ( n4654 & ~n4722 ) | ( n4654 & n4725 ) | ( ~n4722 & n4725 ) ;
  assign n4728 = ( n4722 & ~n4726 ) | ( n4722 & n4727 ) | ( ~n4726 & n4727 ) ;
  assign n4729 = ( n4675 & n4716 ) | ( n4675 & n4728 ) | ( n4716 & n4728 ) ;
  assign n4730 = ( ~n4675 & n4716 ) | ( ~n4675 & n4728 ) | ( n4716 & n4728 ) ;
  assign n4731 = ( n4675 & ~n4729 ) | ( n4675 & n4730 ) | ( ~n4729 & n4730 ) ;
  assign n4732 = ( n4701 & n4713 ) | ( n4701 & n4731 ) | ( n4713 & n4731 ) ;
  assign n4733 = ( ~n4701 & n4713 ) | ( ~n4701 & n4731 ) | ( n4713 & n4731 ) ;
  assign n4734 = ( n4701 & ~n4732 ) | ( n4701 & n4733 ) | ( ~n4732 & n4733 ) ;
  assign n4735 = ( n3850 & ~n3852 ) | ( n3850 & n3854 ) | ( ~n3852 & n3854 ) ;
  assign n4736 = ( n3852 & ~n3855 ) | ( n3852 & n4735 ) | ( ~n3855 & n4735 ) ;
  assign n4737 = ( n4704 & n4734 ) | ( n4704 & n4736 ) | ( n4734 & n4736 ) ;
  assign n4738 = ( ~n3855 & n3857 ) | ( ~n3855 & n3859 ) | ( n3857 & n3859 ) ;
  assign n4739 = ( n3855 & ~n3860 ) | ( n3855 & n4738 ) | ( ~n3860 & n4738 ) ;
  assign n4740 = ( n4706 & n4708 ) | ( n4706 & n4712 ) | ( n4708 & n4712 ) ;
  assign n4741 = ( n4706 & n4708 ) | ( n4706 & ~n4712 ) | ( n4708 & ~n4712 ) ;
  assign n4742 = ( n4712 & ~n4740 ) | ( n4712 & n4741 ) | ( ~n4740 & n4741 ) ;
  assign n4743 = n4717 | n4720 ;
  assign n4744 = n4726 & n4743 ;
  assign n4745 = n4726 | n4743 ;
  assign n4746 = ~n4744 & n4745 ;
  assign n4747 = ( n4714 & n4729 ) | ( n4714 & n4746 ) | ( n4729 & n4746 ) ;
  assign n4748 = ( ~n4714 & n4729 ) | ( ~n4714 & n4746 ) | ( n4729 & n4746 ) ;
  assign n4749 = ( n4714 & ~n4747 ) | ( n4714 & n4748 ) | ( ~n4747 & n4748 ) ;
  assign n4750 = ( n4732 & n4742 ) | ( n4732 & n4749 ) | ( n4742 & n4749 ) ;
  assign n4751 = ( ~n4732 & n4742 ) | ( ~n4732 & n4749 ) | ( n4742 & n4749 ) ;
  assign n4752 = ( n4732 & ~n4750 ) | ( n4732 & n4751 ) | ( ~n4750 & n4751 ) ;
  assign n4753 = ( n4737 & n4739 ) | ( n4737 & n4752 ) | ( n4739 & n4752 ) ;
  assign n4754 = ( n3860 & ~n3862 ) | ( n3860 & n3864 ) | ( ~n3862 & n3864 ) ;
  assign n4755 = ( n3862 & ~n3865 ) | ( n3862 & n4754 ) | ( ~n3865 & n4754 ) ;
  assign n4756 = n4740 | n4744 ;
  assign n4757 = n4740 & n4744 ;
  assign n4758 = n4756 & ~n4757 ;
  assign n4759 = ( n4747 & ~n4750 ) | ( n4747 & n4758 ) | ( ~n4750 & n4758 ) ;
  assign n4760 = ( n4747 & n4750 ) | ( n4747 & n4758 ) | ( n4750 & n4758 ) ;
  assign n4761 = ( n4750 & n4759 ) | ( n4750 & ~n4760 ) | ( n4759 & ~n4760 ) ;
  assign n4762 = ( n4753 & n4755 ) | ( n4753 & n4761 ) | ( n4755 & n4761 ) ;
  assign n4763 = n4747 | n4757 ;
  assign n4764 = ( n4750 & n4756 ) | ( n4750 & n4763 ) | ( n4756 & n4763 ) ;
  assign n4765 = ( n3868 & n4762 ) | ( n3868 & n4764 ) | ( n4762 & n4764 ) ;
  assign n4766 = ( ~n3868 & n4762 ) | ( ~n3868 & n4764 ) | ( n4762 & n4764 ) ;
  assign n4767 = ( n3868 & ~n4765 ) | ( n3868 & n4766 ) | ( ~n4765 & n4766 ) ;
  assign n4768 = n2442 & n4767 ;
  assign n4769 = ( ~n4737 & n4739 ) | ( ~n4737 & n4752 ) | ( n4739 & n4752 ) ;
  assign n4770 = ( n4737 & ~n4753 ) | ( n4737 & n4769 ) | ( ~n4753 & n4769 ) ;
  assign n4771 = ( n4753 & ~n4755 ) | ( n4753 & n4761 ) | ( ~n4755 & n4761 ) ;
  assign n4772 = ( n4755 & ~n4762 ) | ( n4755 & n4771 ) | ( ~n4762 & n4771 ) ;
  assign n4773 = ( ~n1711 & n2435 ) | ( ~n1711 & n2438 ) | ( n2435 & n2438 ) ;
  assign n4774 = ( n1711 & ~n2439 ) | ( n1711 & n4773 ) | ( ~n2439 & n4773 ) ;
  assign n4775 = n4772 | n4774 ;
  assign n4776 = ( ~n4704 & n4734 ) | ( ~n4704 & n4736 ) | ( n4734 & n4736 ) ;
  assign n4777 = ( n4704 & ~n4737 ) | ( n4704 & n4776 ) | ( ~n4737 & n4776 ) ;
  assign n4778 = ( ~n2351 & n2396 ) | ( ~n2351 & n2398 ) | ( n2396 & n2398 ) ;
  assign n4779 = ( n2351 & ~n2399 ) | ( n2351 & n4778 ) | ( ~n2399 & n4778 ) ;
  assign n4780 = ( ~n3830 & n3832 ) | ( ~n3830 & n4267 ) | ( n3832 & n4267 ) ;
  assign n4781 = ( n3830 & ~n4268 ) | ( n3830 & n4780 ) | ( ~n4268 & n4780 ) ;
  assign n4782 = n2044 | n2046 ;
  assign n4783 = ~n2047 & n4782 ;
  assign n4784 = n4781 & n4783 ;
  assign n4785 = ( ~n4269 & n4272 ) | ( ~n4269 & n4506 ) | ( n4272 & n4506 ) ;
  assign n4786 = ( n4269 & ~n4507 ) | ( n4269 & n4785 ) | ( ~n4507 & n4785 ) ;
  assign n4787 = ( n2047 & ~n2239 ) | ( n2047 & n2241 ) | ( ~n2239 & n2241 ) ;
  assign n4788 = ( n2239 & ~n2242 ) | ( n2239 & n4787 ) | ( ~n2242 & n4787 ) ;
  assign n4789 = ( n4784 & n4786 ) | ( n4784 & n4788 ) | ( n4786 & n4788 ) ;
  assign n4790 = ( ~n2242 & n2244 ) | ( ~n2242 & n2350 ) | ( n2244 & n2350 ) ;
  assign n4791 = ( n2242 & ~n2351 ) | ( n2242 & n4790 ) | ( ~n2351 & n4790 ) ;
  assign n4792 = ( ~n4507 & n4509 ) | ( ~n4507 & n4641 ) | ( n4509 & n4641 ) ;
  assign n4793 = ( n4507 & ~n4642 ) | ( n4507 & n4792 ) | ( ~n4642 & n4792 ) ;
  assign n4794 = ( n4789 & n4791 ) | ( n4789 & n4793 ) | ( n4791 & n4793 ) ;
  assign n4795 = ( n4642 & ~n4644 ) | ( n4642 & n4703 ) | ( ~n4644 & n4703 ) ;
  assign n4796 = ( n4644 & ~n4704 ) | ( n4644 & n4795 ) | ( ~n4704 & n4795 ) ;
  assign n4797 = ( n4779 & n4794 ) | ( n4779 & n4796 ) | ( n4794 & n4796 ) ;
  assign n4798 = ( n2399 & ~n2401 ) | ( n2399 & n2422 ) | ( ~n2401 & n2422 ) ;
  assign n4799 = ( n2401 & ~n2423 ) | ( n2401 & n4798 ) | ( ~n2423 & n4798 ) ;
  assign n4800 = ( n4777 & n4797 ) | ( n4777 & n4799 ) | ( n4797 & n4799 ) ;
  assign n4801 = ( n2423 & ~n2425 ) | ( n2423 & n2434 ) | ( ~n2425 & n2434 ) ;
  assign n4802 = ( n2425 & ~n2435 ) | ( n2425 & n4801 ) | ( ~n2435 & n4801 ) ;
  assign n4803 = n4800 | n4802 ;
  assign n4804 = ( n4772 & n4774 ) | ( n4772 & ~n4803 ) | ( n4774 & ~n4803 ) ;
  assign n4805 = n4775 & ~n4804 ;
  assign n4806 = n4770 & ~n4805 ;
  assign n4807 = ( n4779 & n4794 ) | ( n4779 & ~n4796 ) | ( n4794 & ~n4796 ) ;
  assign n4808 = ( n4796 & ~n4797 ) | ( n4796 & n4807 ) | ( ~n4797 & n4807 ) ;
  assign n4809 = n4786 | n4788 ;
  assign n4810 = n4786 & n4788 ;
  assign n4811 = n4809 & ~n4810 ;
  assign n4812 = ( x1000 & n4781 ) | ( x1000 & ~n4811 ) | ( n4781 & ~n4811 ) ;
  assign n4813 = n4783 | n4811 ;
  assign n4814 = ( ~n4784 & n4812 ) | ( ~n4784 & n4813 ) | ( n4812 & n4813 ) ;
  assign n4815 = ( n4789 & n4791 ) | ( n4789 & ~n4793 ) | ( n4791 & ~n4793 ) ;
  assign n4816 = ( n4793 & ~n4794 ) | ( n4793 & n4815 ) | ( ~n4794 & n4815 ) ;
  assign n4817 = n4814 & n4816 ;
  assign n4818 = n4808 | n4817 ;
  assign n4819 = n4800 & n4802 ;
  assign n4820 = ( ~n4770 & n4772 ) | ( ~n4770 & n4774 ) | ( n4772 & n4774 ) ;
  assign n4821 = ( n4775 & n4819 ) | ( n4775 & ~n4820 ) | ( n4819 & ~n4820 ) ;
  assign n4822 = n4818 & ~n4821 ;
  assign n4823 = ( n4806 & n4818 ) | ( n4806 & n4822 ) | ( n4818 & n4822 ) ;
  assign n4824 = ( ~n4777 & n4797 ) | ( ~n4777 & n4799 ) | ( n4797 & n4799 ) ;
  assign n4825 = ( n4777 & ~n4800 ) | ( n4777 & n4824 ) | ( ~n4800 & n4824 ) ;
  assign n4826 = n4805 | n4821 ;
  assign n4827 = n4825 & n4826 ;
  assign n4828 = n4823 & n4827 ;
  assign n4829 = ( n4770 & n4800 ) | ( n4770 & n4802 ) | ( n4800 & n4802 ) ;
  assign n4830 = ( n4772 & n4774 ) | ( n4772 & n4829 ) | ( n4774 & n4829 ) ;
  assign n4831 = ( ~n4768 & n4828 ) | ( ~n4768 & n4830 ) | ( n4828 & n4830 ) ;
  assign n4832 = n4768 & n4831 ;
  assign n4833 = ( n2440 & n3866 ) | ( n2440 & n4765 ) | ( n3866 & n4765 ) ;
  assign n4834 = ( n2442 & n4767 ) | ( n2442 & n4830 ) | ( n4767 & n4830 ) ;
  assign n4835 = n4828 | n4834 ;
  assign n4836 = n2440 | n3866 ;
  assign n4837 = n4765 & ~n4836 ;
  assign n4838 = ( n4835 & n4836 ) | ( n4835 & n4837 ) | ( n4836 & n4837 ) ;
  assign n4839 = ( ~n2442 & n4767 ) | ( ~n2442 & n4830 ) | ( n4767 & n4830 ) ;
  assign n4840 = ( n2442 & n4833 ) | ( n2442 & ~n4839 ) | ( n4833 & ~n4839 ) ;
  assign n4841 = n4839 | n4840 ;
  assign n4842 = ( n4833 & n4838 ) | ( n4833 & n4841 ) | ( n4838 & n4841 ) ;
  assign n4843 = n4832 | n4842 ;
  assign y0 = n4843 ;
endmodule
