module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 ;
  assign n11 = x1 & x3 ;
  assign n12 = x2 | n11 ;
  assign n13 = x6 & ~n12 ;
  assign n14 = ( ~x3 & x9 ) | ( ~x3 & n13 ) | ( x9 & n13 ) ;
  assign n15 = x0 & ~x5 ;
  assign n16 = ( x5 & n14 ) | ( x5 & ~n15 ) | ( n14 & ~n15 ) ;
  assign n17 = x2 | x3 ;
  assign n18 = x0 & ~x9 ;
  assign n19 = n17 | n18 ;
  assign n20 = x6 & n19 ;
  assign n21 = ( ~x0 & x1 ) | ( ~x0 & x9 ) | ( x1 & x9 ) ;
  assign n22 = ~x0 & x9 ;
  assign n23 = ( n20 & n21 ) | ( n20 & ~n22 ) | ( n21 & ~n22 ) ;
  assign n24 = x5 & x6 ;
  assign n25 = n23 | n24 ;
  assign n26 = x2 | x6 ;
  assign n27 = ( x3 & x6 ) | ( x3 & n26 ) | ( x6 & n26 ) ;
  assign n28 = n17 & ~n27 ;
  assign n29 = n25 & ~n28 ;
  assign n30 = ( ~x8 & n16 ) | ( ~x8 & n29 ) | ( n16 & n29 ) ;
  assign n31 = x0 | x1 ;
  assign n32 = n17 | n31 ;
  assign n33 = x4 & ~x7 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = x4 | x7 ;
  assign n36 = n23 & ~n35 ;
  assign n37 = n34 | n36 ;
  assign n38 = ( x8 & ~n29 ) | ( x8 & n37 ) | ( ~n29 & n37 ) ;
  assign n39 = n30 & n38 ;
  assign n40 = x2 & n11 ;
  assign n41 = n17 & ~n40 ;
  assign n42 = x2 & ~x8 ;
  assign n43 = x1 & ~n42 ;
  assign n44 = x8 | x9 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = ~n41 & n45 ;
  assign n47 = x1 & x2 ;
  assign n48 = n18 & ~n47 ;
  assign n49 = ~x1 & x3 ;
  assign n50 = n17 & ~n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = n46 | n51 ;
  assign n53 = x0 | x2 ;
  assign n54 = x5 & ~x6 ;
  assign n55 = ( ~x6 & n53 ) | ( ~x6 & n54 ) | ( n53 & n54 ) ;
  assign n56 = n32 & ~n55 ;
  assign n57 = n52 | n56 ;
  assign n58 = ~x6 & x9 ;
  assign n59 = ~x1 & x9 ;
  assign n60 = x2 & x3 ;
  assign n61 = ( x2 & n59 ) | ( x2 & ~n60 ) | ( n59 & ~n60 ) ;
  assign n62 = n58 | n61 ;
  assign n63 = x3 & x6 ;
  assign n64 = ~n53 & n63 ;
  assign n65 = n31 | n64 ;
  assign n66 = n62 | n65 ;
  assign n67 = ~x0 & x1 ;
  assign n68 = x3 | n67 ;
  assign n69 = ( x1 & x3 ) | ( x1 & n21 ) | ( x3 & n21 ) ;
  assign n70 = x5 | x9 ;
  assign n71 = ( ~x2 & x5 ) | ( ~x2 & n70 ) | ( x5 & n70 ) ;
  assign n72 = ( x5 & ~n69 ) | ( x5 & n71 ) | ( ~n69 & n71 ) ;
  assign n73 = x1 | x3 ;
  assign n74 = ( ~x9 & n71 ) | ( ~x9 & n73 ) | ( n71 & n73 ) ;
  assign n75 = ( ~n68 & n72 ) | ( ~n68 & n74 ) | ( n72 & n74 ) ;
  assign n76 = n66 & ~n75 ;
  assign n77 = n57 & ~n76 ;
  assign n78 = x2 & n31 ;
  assign n79 = x5 | x6 ;
  assign n80 = x3 | n79 ;
  assign n81 = n78 | n80 ;
  assign n82 = x4 | n81 ;
  assign n83 = x1 & ~x9 ;
  assign n84 = x0 | x8 ;
  assign n85 = x0 & x8 ;
  assign n86 = ( n83 & n84 ) | ( n83 & ~n85 ) | ( n84 & ~n85 ) ;
  assign n87 = x2 | n86 ;
  assign n88 = ( n42 & n67 ) | ( n42 & n87 ) | ( n67 & n87 ) ;
  assign n89 = n82 | n88 ;
  assign n90 = ~x7 & x9 ;
  assign n91 = ( ~x7 & x9 ) | ( ~x7 & n86 ) | ( x9 & n86 ) ;
  assign n92 = ( n89 & ~n90 ) | ( n89 & n91 ) | ( ~n90 & n91 ) ;
  assign n93 = ~x5 & n60 ;
  assign n94 = n48 & n93 ;
  assign n95 = x8 | n35 ;
  assign n96 = ( n35 & ~n94 ) | ( n35 & n95 ) | ( ~n94 & n95 ) ;
  assign n97 = n92 & n96 ;
  assign n98 = n77 | n97 ;
  assign n99 = ~n39 & n98 ;
  assign n100 = ~x3 & x5 ;
  assign n101 = ~n57 & n100 ;
  assign n102 = ~x2 & x8 ;
  assign n103 = x0 & n102 ;
  assign n104 = n49 & n54 ;
  assign n105 = ( n54 & n103 ) | ( n54 & n104 ) | ( n103 & n104 ) ;
  assign n106 = ~x9 & n105 ;
  assign n107 = ( ~x9 & n101 ) | ( ~x9 & n106 ) | ( n101 & n106 ) ;
  assign n108 = ~x0 & x8 ;
  assign n109 = x6 | n108 ;
  assign n110 = x5 | n73 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = x6 | n70 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = x8 & x9 ;
  assign n115 = n44 & ~n114 ;
  assign n116 = x0 & ~n11 ;
  assign n117 = n115 & n116 ;
  assign n118 = n12 & ~n117 ;
  assign n119 = ~n113 & n118 ;
  assign n120 = x1 & x5 ;
  assign n121 = x3 | n120 ;
  assign n122 = ( ~x6 & n47 ) | ( ~x6 & n78 ) | ( n47 & n78 ) ;
  assign n123 = ~n121 & n122 ;
  assign n124 = ~n11 & n114 ;
  assign n125 = n85 | n124 ;
  assign n126 = n28 & ~n125 ;
  assign n127 = x5 | x8 ;
  assign n128 = ( n71 & ~n124 ) | ( n71 & n127 ) | ( ~n124 & n127 ) ;
  assign n129 = ~n126 & n128 ;
  assign n130 = n123 & ~n129 ;
  assign n131 = ~x8 & x9 ;
  assign n132 = x5 & n131 ;
  assign n133 = ~n41 & n132 ;
  assign n134 = ~x1 & n44 ;
  assign n135 = ( ~x2 & x6 ) | ( ~x2 & n134 ) | ( x6 & n134 ) ;
  assign n136 = ~n70 & n135 ;
  assign n137 = n133 | n136 ;
  assign n138 = n83 & ~n127 ;
  assign n139 = x1 & x8 ;
  assign n140 = x0 & n139 ;
  assign n141 = ( ~n80 & n138 ) | ( ~n80 & n140 ) | ( n138 & n140 ) ;
  assign n142 = n68 | n141 ;
  assign n143 = ( n137 & n141 ) | ( n137 & n142 ) | ( n141 & n142 ) ;
  assign n144 = n123 | n143 ;
  assign n145 = ( n119 & ~n130 ) | ( n119 & n144 ) | ( ~n130 & n144 ) ;
  assign n146 = n107 | n145 ;
  assign n147 = ~n35 & n146 ;
  assign n148 = ( ~x6 & x9 ) | ( ~x6 & n37 ) | ( x9 & n37 ) ;
  assign n149 = n52 | n117 ;
  assign n150 = x5 | n40 ;
  assign n151 = x2 & ~n150 ;
  assign n152 = ( n149 & n150 ) | ( n149 & ~n151 ) | ( n150 & ~n151 ) ;
  assign n153 = ( x6 & ~x9 ) | ( x6 & n152 ) | ( ~x9 & n152 ) ;
  assign n154 = n148 & n153 ;
  assign n155 = n26 | n73 ;
  assign n156 = ( n42 & n102 ) | ( n42 & n155 ) | ( n102 & n155 ) ;
  assign n157 = ~n62 & n156 ;
  assign n158 = x8 & n63 ;
  assign n159 = ( ~x1 & x8 ) | ( ~x1 & x9 ) | ( x8 & x9 ) ;
  assign n160 = n17 | n159 ;
  assign n161 = ( n83 & ~n158 ) | ( n83 & n160 ) | ( ~n158 & n160 ) ;
  assign n162 = n15 & ~n161 ;
  assign n163 = ( n15 & n157 ) | ( n15 & n162 ) | ( n157 & n162 ) ;
  assign n164 = x2 & ~x6 ;
  assign n165 = n70 & ~n121 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = x6 | n42 ;
  assign n168 = n115 | n167 ;
  assign n169 = n73 | n84 ;
  assign n170 = n168 & ~n169 ;
  assign n171 = ( x0 & ~x5 ) | ( x0 & n116 ) | ( ~x5 & n116 ) ;
  assign n172 = ~n168 & n171 ;
  assign n173 = ( ~n166 & n170 ) | ( ~n166 & n172 ) | ( n170 & n172 ) ;
  assign n174 = n64 & ~n139 ;
  assign n175 = n173 | n174 ;
  assign n176 = n163 | n175 ;
  assign n177 = ( x5 & x8 ) | ( x5 & n59 ) | ( x8 & n59 ) ;
  assign n178 = n164 & ~n177 ;
  assign n179 = n114 & ~n178 ;
  assign n180 = ~n58 & n67 ;
  assign n181 = ~x3 & n164 ;
  assign n182 = ( ~x3 & n180 ) | ( ~x3 & n181 ) | ( n180 & n181 ) ;
  assign n183 = ~n179 & n182 ;
  assign n184 = ~n138 & n183 ;
  assign n185 = n176 | n184 ;
  assign n186 = n35 & n82 ;
  assign n187 = n81 & ~n113 ;
  assign n188 = n35 | n187 ;
  assign n189 = ~n186 & n188 ;
  assign n190 = n185 & ~n189 ;
  assign n191 = ( n154 & n185 ) | ( n154 & ~n190 ) | ( n185 & ~n190 ) ;
  assign n192 = n147 | n191 ;
  assign n193 = x7 & n155 ;
  assign n194 = x4 | n193 ;
  assign n195 = x6 & n47 ;
  assign n196 = n44 & ~n195 ;
  assign n197 = ( ~x2 & n42 ) | ( ~x2 & n70 ) | ( n42 & n70 ) ;
  assign n198 = x3 & n197 ;
  assign n199 = n196 & n198 ;
  assign n200 = n47 & ~n70 ;
  assign n201 = x8 & n200 ;
  assign n202 = n199 | n201 ;
  assign n203 = ~x6 & n43 ;
  assign n204 = x2 & x5 ;
  assign n205 = ~n203 & n204 ;
  assign n206 = n141 | n205 ;
  assign n207 = n202 | n206 ;
  assign n208 = x0 | n194 ;
  assign n209 = n207 & ~n208 ;
  assign n210 = ( n185 & ~n194 ) | ( n185 & n209 ) | ( ~n194 & n209 ) ;
  assign n211 = x7 & n114 ;
  assign n212 = n183 | n211 ;
  assign n213 = ( x0 & x1 ) | ( x0 & ~n159 ) | ( x1 & ~n159 ) ;
  assign n214 = ~n82 & n213 ;
  assign n215 = n212 & n214 ;
  assign n216 = x6 & ~x8 ;
  assign n217 = ( ~x5 & n114 ) | ( ~x5 & n216 ) | ( n114 & n216 ) ;
  assign n218 = n34 & ~n217 ;
  assign n219 = n215 | n218 ;
  assign n220 = n210 | n219 ;
  assign n221 = x3 | x6 ;
  assign n222 = ~x2 & n59 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = ~n108 & n200 ;
  assign n225 = ( ~n108 & n223 ) | ( ~n108 & n224 ) | ( n223 & n224 ) ;
  assign n226 = ~n60 & n225 ;
  assign n227 = x9 & n26 ;
  assign n228 = x8 & ~n227 ;
  assign n229 = n49 | n228 ;
  assign n230 = x1 & n221 ;
  assign n231 = n228 & ~n230 ;
  assign n232 = ( n226 & n229 ) | ( n226 & ~n231 ) | ( n229 & ~n231 ) ;
  assign n233 = ~n24 & n232 ;
  assign n234 = n120 & n168 ;
  assign n235 = ~x6 & n59 ;
  assign n236 = ( x0 & n18 ) | ( x0 & n79 ) | ( n18 & n79 ) ;
  assign n237 = n235 | n236 ;
  assign n238 = ( n183 & ~n234 ) | ( n183 & n237 ) | ( ~n234 & n237 ) ;
  assign n239 = n234 & ~n237 ;
  assign n240 = ( n17 & n237 ) | ( n17 & ~n239 ) | ( n237 & ~n239 ) ;
  assign n241 = ~n238 & n240 ;
  assign n242 = n233 | n241 ;
  assign n243 = n18 & n54 ;
  assign n244 = ~n43 & n243 ;
  assign n245 = ~n52 & n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = ~n79 & n114 ;
  assign n248 = n24 | n247 ;
  assign n249 = n34 & n248 ;
  assign n250 = n35 & ~n249 ;
  assign n251 = ( n246 & n249 ) | ( n246 & ~n250 ) | ( n249 & ~n250 ) ;
  assign n252 = ~x7 & n24 ;
  assign n253 = ( x4 & n17 ) | ( x4 & n252 ) | ( n17 & n252 ) ;
  assign n254 = x2 | n31 ;
  assign n255 = ~n78 & n254 ;
  assign n256 = ( x4 & n17 ) | ( x4 & n255 ) | ( n17 & n255 ) ;
  assign n257 = n253 & ~n256 ;
  assign n258 = ~n35 & n60 ;
  assign n259 = ( n31 & ~n35 ) | ( n31 & n258 ) | ( ~n35 & n258 ) ;
  assign n260 = x3 & n259 ;
  assign n261 = ( n24 & n34 ) | ( n24 & n260 ) | ( n34 & n260 ) ;
  assign n262 = ~n15 & n114 ;
  assign n263 = n11 & ~n262 ;
  assign n264 = n70 | n108 ;
  assign n265 = x2 | n264 ;
  assign n266 = n263 & n265 ;
  assign n267 = n242 & n266 ;
  assign n268 = n17 | n100 ;
  assign n269 = ( n100 & n124 ) | ( n100 & n268 ) | ( n124 & n268 ) ;
  assign n270 = ~n53 & n79 ;
  assign n271 = ~x3 & x6 ;
  assign n272 = x0 & ~n271 ;
  assign n273 = n270 | n272 ;
  assign n274 = n269 & ~n273 ;
  assign n275 = n204 | n221 ;
  assign n276 = n48 & ~n275 ;
  assign n277 = n196 & ~n276 ;
  assign n278 = ~n274 & n277 ;
  assign n279 = n84 & n183 ;
  assign n280 = n23 & n100 ;
  assign n281 = n183 | n280 ;
  assign n282 = ( n278 & n279 ) | ( n278 & ~n281 ) | ( n279 & ~n281 ) ;
  assign n283 = ~n87 & n163 ;
  assign n284 = n44 | n165 ;
  assign n285 = n13 | n284 ;
  assign n286 = ( x0 & x1 ) | ( x0 & n26 ) | ( x1 & n26 ) ;
  assign n287 = ( n31 & n285 ) | ( n31 & ~n286 ) | ( n285 & ~n286 ) ;
  assign n288 = n163 | n287 ;
  assign n289 = ( ~n282 & n283 ) | ( ~n282 & n288 ) | ( n283 & n288 ) ;
  assign n290 = n267 | n289 ;
  assign n291 = n34 | n252 ;
  assign n292 = x7 & ~x9 ;
  assign n293 = ( x2 & ~x8 ) | ( x2 & n292 ) | ( ~x8 & n292 ) ;
  assign n294 = ( ~n82 & n215 ) | ( ~n82 & n293 ) | ( n215 & n293 ) ;
  assign n295 = n291 | n294 ;
  assign n296 = n35 & ~n295 ;
  assign n297 = ( n290 & n295 ) | ( n290 & ~n296 ) | ( n295 & ~n296 ) ;
  assign n298 = n47 & ~n114 ;
  assign n299 = n246 & n298 ;
  assign n300 = x1 & ~n114 ;
  assign n301 = x3 & ~n78 ;
  assign n302 = n196 | n301 ;
  assign n303 = ( x6 & x7 ) | ( x6 & ~n164 ) | ( x7 & ~n164 ) ;
  assign n304 = n302 & n303 ;
  assign n305 = ( ~x1 & n53 ) | ( ~x1 & n114 ) | ( n53 & n114 ) ;
  assign n306 = ( n300 & n304 ) | ( n300 & n305 ) | ( n304 & n305 ) ;
  assign n307 = n141 | n306 ;
  assign n308 = ~n72 & n307 ;
  assign n309 = ( x8 & n59 ) | ( x8 & n60 ) | ( n59 & n60 ) ;
  assign n310 = ( ~n159 & n254 ) | ( ~n159 & n309 ) | ( n254 & n309 ) ;
  assign n311 = n17 | n108 ;
  assign n312 = n54 & n311 ;
  assign n313 = x9 & n105 ;
  assign n314 = n129 & ~n313 ;
  assign n315 = ~n310 & n314 ;
  assign n316 = ( n310 & ~n312 ) | ( n310 & n315 ) | ( ~n312 & n315 ) ;
  assign n317 = ~n308 & n316 ;
  assign n318 = ( n299 & ~n308 ) | ( n299 & n317 ) | ( ~n308 & n317 ) ;
  assign n319 = ~n310 & n312 ;
  assign n320 = ( n35 & ~n134 ) | ( n35 & n186 ) | ( ~n134 & n186 ) ;
  assign n321 = n319 | n320 ;
  assign n322 = n318 | n321 ;
  assign n323 = n213 & n258 ;
  assign n324 = ( n34 & ~n79 ) | ( n34 & n323 ) | ( ~n79 & n323 ) ;
  assign n325 = n322 & ~n324 ;
  assign n326 = n225 & ~n319 ;
  assign n327 = ( n242 & ~n319 ) | ( n242 & n326 ) | ( ~n319 & n326 ) ;
  assign n328 = ~n14 & n203 ;
  assign n329 = n179 & n270 ;
  assign n330 = ( x3 & n178 ) | ( x3 & ~n329 ) | ( n178 & ~n329 ) ;
  assign n331 = n328 | n330 ;
  assign n332 = ( n12 & ~n24 ) | ( n12 & n28 ) | ( ~n24 & n28 ) ;
  assign n333 = n264 & ~n332 ;
  assign n334 = n320 | n333 ;
  assign n335 = n331 & ~n334 ;
  assign n336 = n59 | n114 ;
  assign n337 = n87 | n336 ;
  assign n338 = ( n186 & ~n335 ) | ( n186 & n337 ) | ( ~n335 & n337 ) ;
  assign n339 = n327 | n338 ;
  assign n340 = ~n24 & n34 ;
  assign n341 = n335 | n340 ;
  assign n342 = x6 | n324 ;
  assign n343 = ( n324 & n341 ) | ( n324 & n342 ) | ( n341 & n342 ) ;
  assign n344 = n339 & ~n343 ;
  assign n345 = ~n324 & n341 ;
  assign y0 = ~n99 ;
  assign y1 = n192 ;
  assign y2 = n220 ;
  assign y3 = n251 ;
  assign y4 = n257 ;
  assign y5 = n261 ;
  assign y6 = ~n297 ;
  assign y7 = n325 ;
  assign y8 = n344 ;
  assign y9 = n345 ;
  assign y10 = n324 ;
endmodule
