module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 ;
  assign n129 = ~x56 & x64 ;
  assign n130 = ~x57 & x64 ;
  assign n131 = x126 | x127 ;
  assign n132 = x125 | n131 ;
  assign n133 = x124 | n132 ;
  assign n134 = x123 | n133 ;
  assign n135 = x122 | n134 ;
  assign n136 = x121 | n135 ;
  assign n137 = x120 | n136 ;
  assign n138 = x119 | n137 ;
  assign n139 = x118 | n138 ;
  assign n140 = x117 | n139 ;
  assign n141 = x116 | n140 ;
  assign n142 = x115 | n141 ;
  assign n143 = x114 | n142 ;
  assign n144 = x113 | n143 ;
  assign n145 = x112 | n144 ;
  assign n146 = x111 | n145 ;
  assign n147 = x110 | n146 ;
  assign n148 = x109 | n147 ;
  assign n149 = x108 | n148 ;
  assign n150 = x107 | n149 ;
  assign n151 = x106 | n150 ;
  assign n152 = x105 | n151 ;
  assign n153 = x104 | n152 ;
  assign n154 = x103 | n153 ;
  assign n155 = x102 | n154 ;
  assign n156 = x101 | n155 ;
  assign n157 = x100 | n156 ;
  assign n158 = x99 | n157 ;
  assign n159 = x98 | n158 ;
  assign n160 = x97 | n159 ;
  assign n161 = x96 | n160 ;
  assign n162 = x95 | n161 ;
  assign n163 = x94 | n162 ;
  assign n164 = x93 | n163 ;
  assign n165 = x92 | n164 ;
  assign n166 = x91 | n165 ;
  assign n167 = x90 | n166 ;
  assign n168 = x89 | n167 ;
  assign n169 = x88 | n168 ;
  assign n170 = x87 | n169 ;
  assign n171 = x86 | n170 ;
  assign n172 = x85 | n171 ;
  assign n173 = x84 | n172 ;
  assign n174 = x83 | n173 ;
  assign n175 = x82 | n174 ;
  assign n176 = x81 | n175 ;
  assign n177 = x80 | n176 ;
  assign n178 = x79 | n177 ;
  assign n179 = x78 | n178 ;
  assign n180 = x77 | n179 ;
  assign n181 = x76 | n180 ;
  assign n182 = x75 | n181 ;
  assign n183 = x74 | n182 ;
  assign n184 = x73 | n183 ;
  assign n185 = x72 | n184 ;
  assign n186 = x71 | n185 ;
  assign n187 = x70 | n186 ;
  assign n188 = x69 | n187 ;
  assign n189 = x68 | n188 ;
  assign n190 = x67 | n189 ;
  assign n191 = x64 & ~x65 ;
  assign n192 = ~x62 & x64 ;
  assign n193 = x65 & ~n192 ;
  assign n194 = ( ~x66 & n191 ) | ( ~x66 & n193 ) | ( n191 & n193 ) ;
  assign n195 = x63 | x66 ;
  assign n196 = ( x66 & n194 ) | ( x66 & n195 ) | ( n194 & n195 ) ;
  assign n197 = x65 | x66 ;
  assign n198 = ( ~x63 & x66 ) | ( ~x63 & n197 ) | ( x66 & n197 ) ;
  assign n199 = n190 | n198 ;
  assign n200 = x64 & ~n199 ;
  assign n201 = x62 & ~n200 ;
  assign n202 = ~x61 & x64 ;
  assign n203 = ( x65 & ~n201 ) | ( x65 & n202 ) | ( ~n201 & n202 ) ;
  assign n204 = ( ~x63 & n196 ) | ( ~x63 & n203 ) | ( n196 & n203 ) ;
  assign n205 = n190 | n204 ;
  assign n206 = x63 & ~n194 ;
  assign n207 = ( x63 & n190 ) | ( x63 & n206 ) | ( n190 & n206 ) ;
  assign n208 = ~n197 & n207 ;
  assign n209 = ( n205 & n207 ) | ( n205 & n208 ) | ( n207 & n208 ) ;
  assign n210 = ~x60 & x64 ;
  assign n211 = ~x61 & n205 ;
  assign n212 = ( x61 & ~x64 ) | ( x61 & n205 ) | ( ~x64 & n205 ) ;
  assign n213 = ( n202 & ~n211 ) | ( n202 & n212 ) | ( ~n211 & n212 ) ;
  assign n214 = ( x65 & n210 ) | ( x65 & ~n213 ) | ( n210 & ~n213 ) ;
  assign n215 = ( x65 & n202 ) | ( x65 & ~n205 ) | ( n202 & ~n205 ) ;
  assign n216 = x65 & n202 ;
  assign n217 = ( ~n201 & n215 ) | ( ~n201 & n216 ) | ( n215 & n216 ) ;
  assign n218 = ( n201 & n215 ) | ( n201 & n216 ) | ( n215 & n216 ) ;
  assign n219 = ( n201 & n217 ) | ( n201 & ~n218 ) | ( n217 & ~n218 ) ;
  assign n220 = ( x66 & n214 ) | ( x66 & ~n219 ) | ( n214 & ~n219 ) ;
  assign n221 = ( x67 & ~n189 ) | ( x67 & n220 ) | ( ~n189 & n220 ) ;
  assign n222 = x67 & n220 ;
  assign n223 = ( n209 & ~n221 ) | ( n209 & n222 ) | ( ~n221 & n222 ) ;
  assign n224 = ~x59 & x64 ;
  assign n225 = ( x67 & ~n209 ) | ( x67 & n220 ) | ( ~n209 & n220 ) ;
  assign n226 = n189 | n225 ;
  assign n227 = ~x60 & n226 ;
  assign n228 = ( x60 & ~x64 ) | ( x60 & n226 ) | ( ~x64 & n226 ) ;
  assign n229 = ( n210 & ~n227 ) | ( n210 & n228 ) | ( ~n227 & n228 ) ;
  assign n230 = ( x65 & n224 ) | ( x65 & ~n229 ) | ( n224 & ~n229 ) ;
  assign n231 = ( x65 & n210 ) | ( x65 & n226 ) | ( n210 & n226 ) ;
  assign n232 = x65 | n210 ;
  assign n233 = ( ~n213 & n231 ) | ( ~n213 & n232 ) | ( n231 & n232 ) ;
  assign n234 = ( n213 & n231 ) | ( n213 & n232 ) | ( n231 & n232 ) ;
  assign n235 = ( n213 & n233 ) | ( n213 & ~n234 ) | ( n233 & ~n234 ) ;
  assign n236 = ( x66 & n230 ) | ( x66 & ~n235 ) | ( n230 & ~n235 ) ;
  assign n237 = ( x66 & n214 ) | ( x66 & n226 ) | ( n214 & n226 ) ;
  assign n238 = x66 | n214 ;
  assign n239 = ( ~n219 & n237 ) | ( ~n219 & n238 ) | ( n237 & n238 ) ;
  assign n240 = ( n219 & n237 ) | ( n219 & n238 ) | ( n237 & n238 ) ;
  assign n241 = ( n219 & n239 ) | ( n219 & ~n240 ) | ( n239 & ~n240 ) ;
  assign n242 = ( x67 & n236 ) | ( x67 & ~n241 ) | ( n236 & ~n241 ) ;
  assign n243 = ( x68 & n188 ) | ( x68 & n242 ) | ( n188 & n242 ) ;
  assign n244 = x68 | n242 ;
  assign n245 = ( n223 & n243 ) | ( n223 & ~n244 ) | ( n243 & ~n244 ) ;
  assign n246 = ~x58 & x64 ;
  assign n247 = ( x68 & ~n223 ) | ( x68 & n242 ) | ( ~n223 & n242 ) ;
  assign n248 = n188 | n247 ;
  assign n249 = ~x59 & n248 ;
  assign n250 = ( x59 & ~x64 ) | ( x59 & n248 ) | ( ~x64 & n248 ) ;
  assign n251 = ( n224 & ~n249 ) | ( n224 & n250 ) | ( ~n249 & n250 ) ;
  assign n252 = ( x65 & n246 ) | ( x65 & ~n251 ) | ( n246 & ~n251 ) ;
  assign n253 = ( x65 & n224 ) | ( x65 & n248 ) | ( n224 & n248 ) ;
  assign n254 = x65 | n224 ;
  assign n255 = ( ~n229 & n253 ) | ( ~n229 & n254 ) | ( n253 & n254 ) ;
  assign n256 = ( n229 & n253 ) | ( n229 & n254 ) | ( n253 & n254 ) ;
  assign n257 = ( n229 & n255 ) | ( n229 & ~n256 ) | ( n255 & ~n256 ) ;
  assign n258 = ( x66 & n252 ) | ( x66 & ~n257 ) | ( n252 & ~n257 ) ;
  assign n259 = ( x66 & n230 ) | ( x66 & n248 ) | ( n230 & n248 ) ;
  assign n260 = x66 | n230 ;
  assign n261 = ( ~n235 & n259 ) | ( ~n235 & n260 ) | ( n259 & n260 ) ;
  assign n262 = ( n235 & n259 ) | ( n235 & n260 ) | ( n259 & n260 ) ;
  assign n263 = ( n235 & n261 ) | ( n235 & ~n262 ) | ( n261 & ~n262 ) ;
  assign n264 = ( x67 & n258 ) | ( x67 & ~n263 ) | ( n258 & ~n263 ) ;
  assign n265 = ( x67 & n236 ) | ( x67 & ~n248 ) | ( n236 & ~n248 ) ;
  assign n266 = x67 & n236 ;
  assign n267 = ( ~n241 & n265 ) | ( ~n241 & n266 ) | ( n265 & n266 ) ;
  assign n268 = ( n241 & n265 ) | ( n241 & n266 ) | ( n265 & n266 ) ;
  assign n269 = ( n241 & n267 ) | ( n241 & ~n268 ) | ( n267 & ~n268 ) ;
  assign n270 = ( x68 & n264 ) | ( x68 & ~n269 ) | ( n264 & ~n269 ) ;
  assign n271 = ( x69 & n187 ) | ( x69 & n270 ) | ( n187 & n270 ) ;
  assign n272 = x69 | n270 ;
  assign n273 = ( n245 & n271 ) | ( n245 & ~n272 ) | ( n271 & ~n272 ) ;
  assign n274 = ( x69 & ~n245 ) | ( x69 & n270 ) | ( ~n245 & n270 ) ;
  assign n275 = n187 | n274 ;
  assign n276 = ~x58 & n275 ;
  assign n277 = ( x58 & ~x64 ) | ( x58 & n275 ) | ( ~x64 & n275 ) ;
  assign n278 = ( n246 & ~n276 ) | ( n246 & n277 ) | ( ~n276 & n277 ) ;
  assign n279 = ( x65 & n130 ) | ( x65 & ~n278 ) | ( n130 & ~n278 ) ;
  assign n280 = ( x65 & n246 ) | ( x65 & n275 ) | ( n246 & n275 ) ;
  assign n281 = x65 | n246 ;
  assign n282 = ( ~n251 & n280 ) | ( ~n251 & n281 ) | ( n280 & n281 ) ;
  assign n283 = ( n251 & n280 ) | ( n251 & n281 ) | ( n280 & n281 ) ;
  assign n284 = ( n251 & n282 ) | ( n251 & ~n283 ) | ( n282 & ~n283 ) ;
  assign n285 = ( x66 & n279 ) | ( x66 & ~n284 ) | ( n279 & ~n284 ) ;
  assign n286 = ( x66 & n252 ) | ( x66 & n275 ) | ( n252 & n275 ) ;
  assign n287 = x66 | n252 ;
  assign n288 = ( ~n257 & n286 ) | ( ~n257 & n287 ) | ( n286 & n287 ) ;
  assign n289 = ( n257 & n286 ) | ( n257 & n287 ) | ( n286 & n287 ) ;
  assign n290 = ( n257 & n288 ) | ( n257 & ~n289 ) | ( n288 & ~n289 ) ;
  assign n291 = ( x67 & n285 ) | ( x67 & ~n290 ) | ( n285 & ~n290 ) ;
  assign n292 = ( x67 & n258 ) | ( x67 & n275 ) | ( n258 & n275 ) ;
  assign n293 = x67 | n258 ;
  assign n294 = ( ~n263 & n292 ) | ( ~n263 & n293 ) | ( n292 & n293 ) ;
  assign n295 = ( n263 & n292 ) | ( n263 & n293 ) | ( n292 & n293 ) ;
  assign n296 = ( n263 & n294 ) | ( n263 & ~n295 ) | ( n294 & ~n295 ) ;
  assign n297 = ( x68 & n291 ) | ( x68 & ~n296 ) | ( n291 & ~n296 ) ;
  assign n298 = ( x68 & n264 ) | ( x68 & n275 ) | ( n264 & n275 ) ;
  assign n299 = x68 | n264 ;
  assign n300 = ( ~n269 & n298 ) | ( ~n269 & n299 ) | ( n298 & n299 ) ;
  assign n301 = ( n269 & n298 ) | ( n269 & n299 ) | ( n298 & n299 ) ;
  assign n302 = ( n269 & n300 ) | ( n269 & ~n301 ) | ( n300 & ~n301 ) ;
  assign n303 = ( x69 & n297 ) | ( x69 & ~n302 ) | ( n297 & ~n302 ) ;
  assign n304 = ( x70 & ~n273 ) | ( x70 & n303 ) | ( ~n273 & n303 ) ;
  assign n305 = n186 | n304 ;
  assign n306 = ~x57 & n305 ;
  assign n307 = ( x57 & ~x64 ) | ( x57 & n305 ) | ( ~x64 & n305 ) ;
  assign n308 = ( n130 & ~n306 ) | ( n130 & n307 ) | ( ~n306 & n307 ) ;
  assign n309 = ( x65 & n129 ) | ( x65 & ~n308 ) | ( n129 & ~n308 ) ;
  assign n310 = ( x65 & n130 ) | ( x65 & n305 ) | ( n130 & n305 ) ;
  assign n311 = x65 | n130 ;
  assign n312 = ( ~n278 & n310 ) | ( ~n278 & n311 ) | ( n310 & n311 ) ;
  assign n313 = ( n278 & n310 ) | ( n278 & n311 ) | ( n310 & n311 ) ;
  assign n314 = ( n278 & n312 ) | ( n278 & ~n313 ) | ( n312 & ~n313 ) ;
  assign n315 = ( x66 & n309 ) | ( x66 & ~n314 ) | ( n309 & ~n314 ) ;
  assign n316 = ( x66 & n279 ) | ( x66 & n305 ) | ( n279 & n305 ) ;
  assign n317 = x66 | n279 ;
  assign n318 = ( ~n284 & n316 ) | ( ~n284 & n317 ) | ( n316 & n317 ) ;
  assign n319 = ( n284 & n316 ) | ( n284 & n317 ) | ( n316 & n317 ) ;
  assign n320 = ( n284 & n318 ) | ( n284 & ~n319 ) | ( n318 & ~n319 ) ;
  assign n321 = ( x67 & n315 ) | ( x67 & ~n320 ) | ( n315 & ~n320 ) ;
  assign n322 = ( x67 & n285 ) | ( x67 & n305 ) | ( n285 & n305 ) ;
  assign n323 = x67 | n285 ;
  assign n324 = ( ~n290 & n322 ) | ( ~n290 & n323 ) | ( n322 & n323 ) ;
  assign n325 = ( n290 & n322 ) | ( n290 & n323 ) | ( n322 & n323 ) ;
  assign n326 = ( n290 & n324 ) | ( n290 & ~n325 ) | ( n324 & ~n325 ) ;
  assign n327 = ( x68 & n321 ) | ( x68 & ~n326 ) | ( n321 & ~n326 ) ;
  assign n328 = ( x68 & n291 ) | ( x68 & ~n305 ) | ( n291 & ~n305 ) ;
  assign n329 = x68 & n291 ;
  assign n330 = ( ~n296 & n328 ) | ( ~n296 & n329 ) | ( n328 & n329 ) ;
  assign n331 = ( n296 & n328 ) | ( n296 & n329 ) | ( n328 & n329 ) ;
  assign n332 = ( n296 & n330 ) | ( n296 & ~n331 ) | ( n330 & ~n331 ) ;
  assign n333 = ( x69 & n327 ) | ( x69 & ~n332 ) | ( n327 & ~n332 ) ;
  assign n334 = ( x69 & n297 ) | ( x69 & ~n305 ) | ( n297 & ~n305 ) ;
  assign n335 = x69 & n297 ;
  assign n336 = ( ~n302 & n334 ) | ( ~n302 & n335 ) | ( n334 & n335 ) ;
  assign n337 = ( n302 & n334 ) | ( n302 & n335 ) | ( n334 & n335 ) ;
  assign n338 = ( n302 & n336 ) | ( n302 & ~n337 ) | ( n336 & ~n337 ) ;
  assign n339 = ( x70 & n333 ) | ( x70 & ~n338 ) | ( n333 & ~n338 ) ;
  assign n340 = ( x70 & n186 ) | ( x70 & n303 ) | ( n186 & n303 ) ;
  assign n341 = x70 | n303 ;
  assign n342 = ( n273 & n340 ) | ( n273 & ~n341 ) | ( n340 & ~n341 ) ;
  assign n343 = ( ~x71 & n339 ) | ( ~x71 & n342 ) | ( n339 & n342 ) ;
  assign n344 = ( ~x71 & n185 ) | ( ~x71 & n339 ) | ( n185 & n339 ) ;
  assign n345 = n343 & ~n344 ;
  assign n346 = ~x55 & x64 ;
  assign n347 = ( x71 & n339 ) | ( x71 & ~n342 ) | ( n339 & ~n342 ) ;
  assign n348 = n185 | n347 ;
  assign n349 = ~x56 & n348 ;
  assign n350 = ( x56 & ~x64 ) | ( x56 & n348 ) | ( ~x64 & n348 ) ;
  assign n351 = ( n129 & ~n349 ) | ( n129 & n350 ) | ( ~n349 & n350 ) ;
  assign n352 = ( x65 & n346 ) | ( x65 & ~n351 ) | ( n346 & ~n351 ) ;
  assign n353 = ( x65 & n129 ) | ( x65 & n348 ) | ( n129 & n348 ) ;
  assign n354 = x65 | n129 ;
  assign n355 = ( ~n308 & n353 ) | ( ~n308 & n354 ) | ( n353 & n354 ) ;
  assign n356 = ( n308 & n353 ) | ( n308 & n354 ) | ( n353 & n354 ) ;
  assign n357 = ( n308 & n355 ) | ( n308 & ~n356 ) | ( n355 & ~n356 ) ;
  assign n358 = ( x66 & n352 ) | ( x66 & ~n357 ) | ( n352 & ~n357 ) ;
  assign n359 = ( x66 & n309 ) | ( x66 & n348 ) | ( n309 & n348 ) ;
  assign n360 = x66 | n309 ;
  assign n361 = ( ~n314 & n359 ) | ( ~n314 & n360 ) | ( n359 & n360 ) ;
  assign n362 = ( n314 & n359 ) | ( n314 & n360 ) | ( n359 & n360 ) ;
  assign n363 = ( n314 & n361 ) | ( n314 & ~n362 ) | ( n361 & ~n362 ) ;
  assign n364 = ( x67 & n358 ) | ( x67 & ~n363 ) | ( n358 & ~n363 ) ;
  assign n365 = ( x67 & n315 ) | ( x67 & ~n348 ) | ( n315 & ~n348 ) ;
  assign n366 = x67 & n315 ;
  assign n367 = ( ~n320 & n365 ) | ( ~n320 & n366 ) | ( n365 & n366 ) ;
  assign n368 = ( n320 & n365 ) | ( n320 & n366 ) | ( n365 & n366 ) ;
  assign n369 = ( n320 & n367 ) | ( n320 & ~n368 ) | ( n367 & ~n368 ) ;
  assign n370 = ( x68 & n364 ) | ( x68 & ~n369 ) | ( n364 & ~n369 ) ;
  assign n371 = ( x68 & n321 ) | ( x68 & ~n348 ) | ( n321 & ~n348 ) ;
  assign n372 = x68 & n321 ;
  assign n373 = ( ~n326 & n371 ) | ( ~n326 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( n326 & n371 ) | ( n326 & n372 ) | ( n371 & n372 ) ;
  assign n375 = ( n326 & n373 ) | ( n326 & ~n374 ) | ( n373 & ~n374 ) ;
  assign n376 = ( x69 & n370 ) | ( x69 & ~n375 ) | ( n370 & ~n375 ) ;
  assign n377 = ( x69 & n327 ) | ( x69 & ~n348 ) | ( n327 & ~n348 ) ;
  assign n378 = x69 & n327 ;
  assign n379 = ( ~n332 & n377 ) | ( ~n332 & n378 ) | ( n377 & n378 ) ;
  assign n380 = ( n332 & n377 ) | ( n332 & n378 ) | ( n377 & n378 ) ;
  assign n381 = ( n332 & n379 ) | ( n332 & ~n380 ) | ( n379 & ~n380 ) ;
  assign n382 = ( x70 & n376 ) | ( x70 & ~n381 ) | ( n376 & ~n381 ) ;
  assign n383 = ( x70 & n333 ) | ( x70 & ~n348 ) | ( n333 & ~n348 ) ;
  assign n384 = x70 & n333 ;
  assign n385 = ( ~n338 & n383 ) | ( ~n338 & n384 ) | ( n383 & n384 ) ;
  assign n386 = ( n338 & n383 ) | ( n338 & n384 ) | ( n383 & n384 ) ;
  assign n387 = ( n338 & n385 ) | ( n338 & ~n386 ) | ( n385 & ~n386 ) ;
  assign n388 = ( x71 & n382 ) | ( x71 & ~n387 ) | ( n382 & ~n387 ) ;
  assign n389 = n345 & ~n388 ;
  assign n390 = ~x1 & x64 ;
  assign n391 = ~x2 & x64 ;
  assign n392 = ( n184 & n185 ) | ( n184 & ~n342 ) | ( n185 & ~n342 ) ;
  assign n393 = ( ~n345 & n388 ) | ( ~n345 & n392 ) | ( n388 & n392 ) ;
  assign n394 = ( x71 & n382 ) | ( x71 & ~n393 ) | ( n382 & ~n393 ) ;
  assign n395 = x71 & n382 ;
  assign n396 = ( ~n387 & n394 ) | ( ~n387 & n395 ) | ( n394 & n395 ) ;
  assign n397 = ( n387 & n394 ) | ( n387 & n395 ) | ( n394 & n395 ) ;
  assign n398 = ( n387 & n396 ) | ( n387 & ~n397 ) | ( n396 & ~n397 ) ;
  assign n399 = ~x54 & x64 ;
  assign n400 = ~x55 & n393 ;
  assign n401 = ( x55 & ~x64 ) | ( x55 & n393 ) | ( ~x64 & n393 ) ;
  assign n402 = ( n346 & ~n400 ) | ( n346 & n401 ) | ( ~n400 & n401 ) ;
  assign n403 = ( x65 & n399 ) | ( x65 & ~n402 ) | ( n399 & ~n402 ) ;
  assign n404 = ( x65 & n346 ) | ( x65 & n393 ) | ( n346 & n393 ) ;
  assign n405 = x65 | n346 ;
  assign n406 = ( ~n351 & n404 ) | ( ~n351 & n405 ) | ( n404 & n405 ) ;
  assign n407 = ( n351 & n404 ) | ( n351 & n405 ) | ( n404 & n405 ) ;
  assign n408 = ( n351 & n406 ) | ( n351 & ~n407 ) | ( n406 & ~n407 ) ;
  assign n409 = ( x66 & n403 ) | ( x66 & ~n408 ) | ( n403 & ~n408 ) ;
  assign n410 = ( x66 & n352 ) | ( x66 & n393 ) | ( n352 & n393 ) ;
  assign n411 = x66 | n352 ;
  assign n412 = ( ~n357 & n410 ) | ( ~n357 & n411 ) | ( n410 & n411 ) ;
  assign n413 = ( n357 & n410 ) | ( n357 & n411 ) | ( n410 & n411 ) ;
  assign n414 = ( n357 & n412 ) | ( n357 & ~n413 ) | ( n412 & ~n413 ) ;
  assign n415 = ( x67 & n409 ) | ( x67 & ~n414 ) | ( n409 & ~n414 ) ;
  assign n416 = ( x67 & n358 ) | ( x67 & ~n393 ) | ( n358 & ~n393 ) ;
  assign n417 = x67 & n358 ;
  assign n418 = ( ~n363 & n416 ) | ( ~n363 & n417 ) | ( n416 & n417 ) ;
  assign n419 = ( n363 & n416 ) | ( n363 & n417 ) | ( n416 & n417 ) ;
  assign n420 = ( n363 & n418 ) | ( n363 & ~n419 ) | ( n418 & ~n419 ) ;
  assign n421 = ( x68 & n415 ) | ( x68 & ~n420 ) | ( n415 & ~n420 ) ;
  assign n422 = ( x68 & n364 ) | ( x68 & ~n393 ) | ( n364 & ~n393 ) ;
  assign n423 = x68 & n364 ;
  assign n424 = ( ~n369 & n422 ) | ( ~n369 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ( n369 & n422 ) | ( n369 & n423 ) | ( n422 & n423 ) ;
  assign n426 = ( n369 & n424 ) | ( n369 & ~n425 ) | ( n424 & ~n425 ) ;
  assign n427 = ( x69 & n421 ) | ( x69 & ~n426 ) | ( n421 & ~n426 ) ;
  assign n428 = ( x69 & n370 ) | ( x69 & ~n393 ) | ( n370 & ~n393 ) ;
  assign n429 = x69 & n370 ;
  assign n430 = ( ~n375 & n428 ) | ( ~n375 & n429 ) | ( n428 & n429 ) ;
  assign n431 = ( n375 & n428 ) | ( n375 & n429 ) | ( n428 & n429 ) ;
  assign n432 = ( n375 & n430 ) | ( n375 & ~n431 ) | ( n430 & ~n431 ) ;
  assign n433 = ( x70 & n427 ) | ( x70 & ~n432 ) | ( n427 & ~n432 ) ;
  assign n434 = ( x70 & n376 ) | ( x70 & ~n393 ) | ( n376 & ~n393 ) ;
  assign n435 = x70 & n376 ;
  assign n436 = ( ~n381 & n434 ) | ( ~n381 & n435 ) | ( n434 & n435 ) ;
  assign n437 = ( n381 & n434 ) | ( n381 & n435 ) | ( n434 & n435 ) ;
  assign n438 = ( n381 & n436 ) | ( n381 & ~n437 ) | ( n436 & ~n437 ) ;
  assign n439 = ( x71 & n433 ) | ( x71 & ~n438 ) | ( n433 & ~n438 ) ;
  assign n440 = ( x72 & ~n398 ) | ( x72 & n439 ) | ( ~n398 & n439 ) ;
  assign n441 = ( n184 & n185 ) | ( n184 & n388 ) | ( n185 & n388 ) ;
  assign n442 = n342 & n441 ;
  assign n443 = n389 | n442 ;
  assign n444 = ( x73 & n440 ) | ( x73 & ~n443 ) | ( n440 & ~n443 ) ;
  assign n445 = n183 | n444 ;
  assign n446 = ( x72 & n439 ) | ( x72 & n445 ) | ( n439 & n445 ) ;
  assign n447 = x72 | n439 ;
  assign n448 = ( ~n398 & n446 ) | ( ~n398 & n447 ) | ( n446 & n447 ) ;
  assign n449 = ( n398 & n446 ) | ( n398 & n447 ) | ( n446 & n447 ) ;
  assign n450 = ( n398 & n448 ) | ( n398 & ~n449 ) | ( n448 & ~n449 ) ;
  assign n451 = ~x53 & x64 ;
  assign n452 = ~x54 & n445 ;
  assign n453 = ( x54 & ~x64 ) | ( x54 & n445 ) | ( ~x64 & n445 ) ;
  assign n454 = ( n399 & ~n452 ) | ( n399 & n453 ) | ( ~n452 & n453 ) ;
  assign n455 = ( x65 & n451 ) | ( x65 & ~n454 ) | ( n451 & ~n454 ) ;
  assign n456 = ( x65 & n399 ) | ( x65 & n445 ) | ( n399 & n445 ) ;
  assign n457 = x65 | n399 ;
  assign n458 = ( ~n402 & n456 ) | ( ~n402 & n457 ) | ( n456 & n457 ) ;
  assign n459 = ( n402 & n456 ) | ( n402 & n457 ) | ( n456 & n457 ) ;
  assign n460 = ( n402 & n458 ) | ( n402 & ~n459 ) | ( n458 & ~n459 ) ;
  assign n461 = ( x66 & n455 ) | ( x66 & ~n460 ) | ( n455 & ~n460 ) ;
  assign n462 = ( x66 & n403 ) | ( x66 & n445 ) | ( n403 & n445 ) ;
  assign n463 = x66 | n403 ;
  assign n464 = ( ~n408 & n462 ) | ( ~n408 & n463 ) | ( n462 & n463 ) ;
  assign n465 = ( n408 & n462 ) | ( n408 & n463 ) | ( n462 & n463 ) ;
  assign n466 = ( n408 & n464 ) | ( n408 & ~n465 ) | ( n464 & ~n465 ) ;
  assign n467 = ( x67 & n461 ) | ( x67 & ~n466 ) | ( n461 & ~n466 ) ;
  assign n468 = ( x67 & n409 ) | ( x67 & ~n445 ) | ( n409 & ~n445 ) ;
  assign n469 = x67 & n409 ;
  assign n470 = ( ~n414 & n468 ) | ( ~n414 & n469 ) | ( n468 & n469 ) ;
  assign n471 = ( n414 & n468 ) | ( n414 & n469 ) | ( n468 & n469 ) ;
  assign n472 = ( n414 & n470 ) | ( n414 & ~n471 ) | ( n470 & ~n471 ) ;
  assign n473 = ( x68 & n467 ) | ( x68 & ~n472 ) | ( n467 & ~n472 ) ;
  assign n474 = ( x68 & n415 ) | ( x68 & ~n445 ) | ( n415 & ~n445 ) ;
  assign n475 = x68 & n415 ;
  assign n476 = ( ~n420 & n474 ) | ( ~n420 & n475 ) | ( n474 & n475 ) ;
  assign n477 = ( n420 & n474 ) | ( n420 & n475 ) | ( n474 & n475 ) ;
  assign n478 = ( n420 & n476 ) | ( n420 & ~n477 ) | ( n476 & ~n477 ) ;
  assign n479 = ( x69 & n473 ) | ( x69 & ~n478 ) | ( n473 & ~n478 ) ;
  assign n480 = ( x69 & n421 ) | ( x69 & ~n445 ) | ( n421 & ~n445 ) ;
  assign n481 = x69 & n421 ;
  assign n482 = ( ~n426 & n480 ) | ( ~n426 & n481 ) | ( n480 & n481 ) ;
  assign n483 = ( n426 & n480 ) | ( n426 & n481 ) | ( n480 & n481 ) ;
  assign n484 = ( n426 & n482 ) | ( n426 & ~n483 ) | ( n482 & ~n483 ) ;
  assign n485 = ( x70 & n479 ) | ( x70 & ~n484 ) | ( n479 & ~n484 ) ;
  assign n486 = ( x70 & n427 ) | ( x70 & ~n445 ) | ( n427 & ~n445 ) ;
  assign n487 = x70 & n427 ;
  assign n488 = ( ~n432 & n486 ) | ( ~n432 & n487 ) | ( n486 & n487 ) ;
  assign n489 = ( n432 & n486 ) | ( n432 & n487 ) | ( n486 & n487 ) ;
  assign n490 = ( n432 & n488 ) | ( n432 & ~n489 ) | ( n488 & ~n489 ) ;
  assign n491 = ( x71 & n485 ) | ( x71 & ~n490 ) | ( n485 & ~n490 ) ;
  assign n492 = ( x71 & n433 ) | ( x71 & ~n445 ) | ( n433 & ~n445 ) ;
  assign n493 = x71 & n433 ;
  assign n494 = ( ~n438 & n492 ) | ( ~n438 & n493 ) | ( n492 & n493 ) ;
  assign n495 = ( n438 & n492 ) | ( n438 & n493 ) | ( n492 & n493 ) ;
  assign n496 = ( n438 & n494 ) | ( n438 & ~n495 ) | ( n494 & ~n495 ) ;
  assign n497 = ( x72 & n491 ) | ( x72 & ~n496 ) | ( n491 & ~n496 ) ;
  assign n498 = ( x73 & n183 ) | ( x73 & n440 ) | ( n183 & n440 ) ;
  assign n499 = x73 | n440 ;
  assign n500 = ( n443 & n498 ) | ( n443 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = ( x73 & ~n450 ) | ( x73 & n497 ) | ( ~n450 & n497 ) ;
  assign n502 = ( x74 & ~n500 ) | ( x74 & n501 ) | ( ~n500 & n501 ) ;
  assign n503 = n182 | n502 ;
  assign n504 = ( x73 & n497 ) | ( x73 & n503 ) | ( n497 & n503 ) ;
  assign n505 = x73 | n497 ;
  assign n506 = ( ~n450 & n504 ) | ( ~n450 & n505 ) | ( n504 & n505 ) ;
  assign n507 = ( n450 & n504 ) | ( n450 & n505 ) | ( n504 & n505 ) ;
  assign n508 = ( n450 & n506 ) | ( n450 & ~n507 ) | ( n506 & ~n507 ) ;
  assign n509 = ~x52 & x64 ;
  assign n510 = ~x53 & n503 ;
  assign n511 = ( x53 & ~x64 ) | ( x53 & n503 ) | ( ~x64 & n503 ) ;
  assign n512 = ( n451 & ~n510 ) | ( n451 & n511 ) | ( ~n510 & n511 ) ;
  assign n513 = ( x65 & n509 ) | ( x65 & ~n512 ) | ( n509 & ~n512 ) ;
  assign n514 = ( x65 & n451 ) | ( x65 & n503 ) | ( n451 & n503 ) ;
  assign n515 = x65 | n451 ;
  assign n516 = ( ~n454 & n514 ) | ( ~n454 & n515 ) | ( n514 & n515 ) ;
  assign n517 = ( n454 & n514 ) | ( n454 & n515 ) | ( n514 & n515 ) ;
  assign n518 = ( n454 & n516 ) | ( n454 & ~n517 ) | ( n516 & ~n517 ) ;
  assign n519 = ( x66 & n513 ) | ( x66 & ~n518 ) | ( n513 & ~n518 ) ;
  assign n520 = ( x66 & n455 ) | ( x66 & n503 ) | ( n455 & n503 ) ;
  assign n521 = x66 | n455 ;
  assign n522 = ( ~n460 & n520 ) | ( ~n460 & n521 ) | ( n520 & n521 ) ;
  assign n523 = ( n460 & n520 ) | ( n460 & n521 ) | ( n520 & n521 ) ;
  assign n524 = ( n460 & n522 ) | ( n460 & ~n523 ) | ( n522 & ~n523 ) ;
  assign n525 = ( x67 & n519 ) | ( x67 & ~n524 ) | ( n519 & ~n524 ) ;
  assign n526 = ( x67 & n461 ) | ( x67 & ~n503 ) | ( n461 & ~n503 ) ;
  assign n527 = x67 & n461 ;
  assign n528 = ( ~n466 & n526 ) | ( ~n466 & n527 ) | ( n526 & n527 ) ;
  assign n529 = ( n466 & n526 ) | ( n466 & n527 ) | ( n526 & n527 ) ;
  assign n530 = ( n466 & n528 ) | ( n466 & ~n529 ) | ( n528 & ~n529 ) ;
  assign n531 = ( x68 & n525 ) | ( x68 & ~n530 ) | ( n525 & ~n530 ) ;
  assign n532 = ( x68 & n467 ) | ( x68 & ~n503 ) | ( n467 & ~n503 ) ;
  assign n533 = x68 & n467 ;
  assign n534 = ( ~n472 & n532 ) | ( ~n472 & n533 ) | ( n532 & n533 ) ;
  assign n535 = ( n472 & n532 ) | ( n472 & n533 ) | ( n532 & n533 ) ;
  assign n536 = ( n472 & n534 ) | ( n472 & ~n535 ) | ( n534 & ~n535 ) ;
  assign n537 = ( x69 & n531 ) | ( x69 & ~n536 ) | ( n531 & ~n536 ) ;
  assign n538 = ( x69 & n473 ) | ( x69 & ~n503 ) | ( n473 & ~n503 ) ;
  assign n539 = x69 & n473 ;
  assign n540 = ( ~n478 & n538 ) | ( ~n478 & n539 ) | ( n538 & n539 ) ;
  assign n541 = ( n478 & n538 ) | ( n478 & n539 ) | ( n538 & n539 ) ;
  assign n542 = ( n478 & n540 ) | ( n478 & ~n541 ) | ( n540 & ~n541 ) ;
  assign n543 = ( x70 & n537 ) | ( x70 & ~n542 ) | ( n537 & ~n542 ) ;
  assign n544 = ( x70 & n479 ) | ( x70 & ~n503 ) | ( n479 & ~n503 ) ;
  assign n545 = x70 & n479 ;
  assign n546 = ( ~n484 & n544 ) | ( ~n484 & n545 ) | ( n544 & n545 ) ;
  assign n547 = ( n484 & n544 ) | ( n484 & n545 ) | ( n544 & n545 ) ;
  assign n548 = ( n484 & n546 ) | ( n484 & ~n547 ) | ( n546 & ~n547 ) ;
  assign n549 = ( x71 & n543 ) | ( x71 & ~n548 ) | ( n543 & ~n548 ) ;
  assign n550 = ( x71 & n485 ) | ( x71 & ~n503 ) | ( n485 & ~n503 ) ;
  assign n551 = x71 & n485 ;
  assign n552 = ( ~n490 & n550 ) | ( ~n490 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( n490 & n550 ) | ( n490 & n551 ) | ( n550 & n551 ) ;
  assign n554 = ( n490 & n552 ) | ( n490 & ~n553 ) | ( n552 & ~n553 ) ;
  assign n555 = ( x72 & n549 ) | ( x72 & ~n554 ) | ( n549 & ~n554 ) ;
  assign n556 = ( x72 & n491 ) | ( x72 & ~n503 ) | ( n491 & ~n503 ) ;
  assign n557 = x72 & n491 ;
  assign n558 = ( ~n496 & n556 ) | ( ~n496 & n557 ) | ( n556 & n557 ) ;
  assign n559 = ( n496 & n556 ) | ( n496 & n557 ) | ( n556 & n557 ) ;
  assign n560 = ( n496 & n558 ) | ( n496 & ~n559 ) | ( n558 & ~n559 ) ;
  assign n561 = ( x73 & n555 ) | ( x73 & ~n560 ) | ( n555 & ~n560 ) ;
  assign n562 = ( n181 & n182 ) | ( n181 & ~n500 ) | ( n182 & ~n500 ) ;
  assign n563 = ( x74 & ~n508 ) | ( x74 & n561 ) | ( ~n508 & n561 ) ;
  assign n564 = ( ~x74 & n182 ) | ( ~x74 & n501 ) | ( n182 & n501 ) ;
  assign n565 = ( ~x74 & n500 ) | ( ~x74 & n501 ) | ( n500 & n501 ) ;
  assign n566 = ~n564 & n565 ;
  assign n567 = ~n562 & n566 ;
  assign n568 = ( n562 & n563 ) | ( n562 & ~n567 ) | ( n563 & ~n567 ) ;
  assign n569 = ( x74 & n561 ) | ( x74 & n568 ) | ( n561 & n568 ) ;
  assign n570 = x74 | n561 ;
  assign n571 = ( ~n508 & n569 ) | ( ~n508 & n570 ) | ( n569 & n570 ) ;
  assign n572 = ( n508 & n569 ) | ( n508 & n570 ) | ( n569 & n570 ) ;
  assign n573 = ( n508 & n571 ) | ( n508 & ~n572 ) | ( n571 & ~n572 ) ;
  assign n574 = ~x51 & x64 ;
  assign n575 = ~x52 & n568 ;
  assign n576 = ( x52 & ~x64 ) | ( x52 & n568 ) | ( ~x64 & n568 ) ;
  assign n577 = ( n509 & ~n575 ) | ( n509 & n576 ) | ( ~n575 & n576 ) ;
  assign n578 = ( x65 & n574 ) | ( x65 & ~n577 ) | ( n574 & ~n577 ) ;
  assign n579 = ( x65 & n509 ) | ( x65 & n568 ) | ( n509 & n568 ) ;
  assign n580 = x65 | n509 ;
  assign n581 = ( ~n512 & n579 ) | ( ~n512 & n580 ) | ( n579 & n580 ) ;
  assign n582 = ( n512 & n579 ) | ( n512 & n580 ) | ( n579 & n580 ) ;
  assign n583 = ( n512 & n581 ) | ( n512 & ~n582 ) | ( n581 & ~n582 ) ;
  assign n584 = ( x66 & n578 ) | ( x66 & ~n583 ) | ( n578 & ~n583 ) ;
  assign n585 = ( x66 & n513 ) | ( x66 & n568 ) | ( n513 & n568 ) ;
  assign n586 = x66 | n513 ;
  assign n587 = ( ~n518 & n585 ) | ( ~n518 & n586 ) | ( n585 & n586 ) ;
  assign n588 = ( n518 & n585 ) | ( n518 & n586 ) | ( n585 & n586 ) ;
  assign n589 = ( n518 & n587 ) | ( n518 & ~n588 ) | ( n587 & ~n588 ) ;
  assign n590 = ( x67 & n584 ) | ( x67 & ~n589 ) | ( n584 & ~n589 ) ;
  assign n591 = ( x67 & n519 ) | ( x67 & n568 ) | ( n519 & n568 ) ;
  assign n592 = x67 | n519 ;
  assign n593 = ( ~n524 & n591 ) | ( ~n524 & n592 ) | ( n591 & n592 ) ;
  assign n594 = ( n524 & n591 ) | ( n524 & n592 ) | ( n591 & n592 ) ;
  assign n595 = ( n524 & n593 ) | ( n524 & ~n594 ) | ( n593 & ~n594 ) ;
  assign n596 = ( x68 & n590 ) | ( x68 & ~n595 ) | ( n590 & ~n595 ) ;
  assign n597 = ( x68 & n525 ) | ( x68 & ~n568 ) | ( n525 & ~n568 ) ;
  assign n598 = x68 & n525 ;
  assign n599 = ( ~n530 & n597 ) | ( ~n530 & n598 ) | ( n597 & n598 ) ;
  assign n600 = ( n530 & n597 ) | ( n530 & n598 ) | ( n597 & n598 ) ;
  assign n601 = ( n530 & n599 ) | ( n530 & ~n600 ) | ( n599 & ~n600 ) ;
  assign n602 = ( x69 & n596 ) | ( x69 & ~n601 ) | ( n596 & ~n601 ) ;
  assign n603 = ( x69 & n531 ) | ( x69 & ~n568 ) | ( n531 & ~n568 ) ;
  assign n604 = x69 & n531 ;
  assign n605 = ( ~n536 & n603 ) | ( ~n536 & n604 ) | ( n603 & n604 ) ;
  assign n606 = ( n536 & n603 ) | ( n536 & n604 ) | ( n603 & n604 ) ;
  assign n607 = ( n536 & n605 ) | ( n536 & ~n606 ) | ( n605 & ~n606 ) ;
  assign n608 = ( x70 & n602 ) | ( x70 & ~n607 ) | ( n602 & ~n607 ) ;
  assign n609 = ( x70 & n537 ) | ( x70 & ~n568 ) | ( n537 & ~n568 ) ;
  assign n610 = x70 & n537 ;
  assign n611 = ( ~n542 & n609 ) | ( ~n542 & n610 ) | ( n609 & n610 ) ;
  assign n612 = ( n542 & n609 ) | ( n542 & n610 ) | ( n609 & n610 ) ;
  assign n613 = ( n542 & n611 ) | ( n542 & ~n612 ) | ( n611 & ~n612 ) ;
  assign n614 = ( x71 & n608 ) | ( x71 & ~n613 ) | ( n608 & ~n613 ) ;
  assign n615 = ( x71 & n543 ) | ( x71 & ~n568 ) | ( n543 & ~n568 ) ;
  assign n616 = x71 & n543 ;
  assign n617 = ( ~n548 & n615 ) | ( ~n548 & n616 ) | ( n615 & n616 ) ;
  assign n618 = ( n548 & n615 ) | ( n548 & n616 ) | ( n615 & n616 ) ;
  assign n619 = ( n548 & n617 ) | ( n548 & ~n618 ) | ( n617 & ~n618 ) ;
  assign n620 = ( x72 & n614 ) | ( x72 & ~n619 ) | ( n614 & ~n619 ) ;
  assign n621 = ( x72 & n549 ) | ( x72 & ~n568 ) | ( n549 & ~n568 ) ;
  assign n622 = x72 & n549 ;
  assign n623 = ( ~n554 & n621 ) | ( ~n554 & n622 ) | ( n621 & n622 ) ;
  assign n624 = ( n554 & n621 ) | ( n554 & n622 ) | ( n621 & n622 ) ;
  assign n625 = ( n554 & n623 ) | ( n554 & ~n624 ) | ( n623 & ~n624 ) ;
  assign n626 = ( x73 & n620 ) | ( x73 & ~n625 ) | ( n620 & ~n625 ) ;
  assign n627 = ( x73 & n555 ) | ( x73 & ~n568 ) | ( n555 & ~n568 ) ;
  assign n628 = x73 & n555 ;
  assign n629 = ( ~n560 & n627 ) | ( ~n560 & n628 ) | ( n627 & n628 ) ;
  assign n630 = ( n560 & n627 ) | ( n560 & n628 ) | ( n627 & n628 ) ;
  assign n631 = ( n560 & n629 ) | ( n560 & ~n630 ) | ( n629 & ~n630 ) ;
  assign n632 = ( x74 & n626 ) | ( x74 & ~n631 ) | ( n626 & ~n631 ) ;
  assign n633 = ( x75 & ~n573 ) | ( x75 & n632 ) | ( ~n573 & n632 ) ;
  assign n634 = ( n181 & n182 ) | ( n181 & n563 ) | ( n182 & n563 ) ;
  assign n635 = n500 & n634 ;
  assign n636 = n389 | n635 ;
  assign n637 = ( x76 & n633 ) | ( x76 & ~n636 ) | ( n633 & ~n636 ) ;
  assign n638 = n180 | n637 ;
  assign n639 = ( x75 & n632 ) | ( x75 & n638 ) | ( n632 & n638 ) ;
  assign n640 = x75 | n632 ;
  assign n641 = ( ~n573 & n639 ) | ( ~n573 & n640 ) | ( n639 & n640 ) ;
  assign n642 = ( n573 & n639 ) | ( n573 & n640 ) | ( n639 & n640 ) ;
  assign n643 = ( n573 & n641 ) | ( n573 & ~n642 ) | ( n641 & ~n642 ) ;
  assign n644 = ~x50 & x64 ;
  assign n645 = ~x51 & n638 ;
  assign n646 = ( x51 & ~x64 ) | ( x51 & n638 ) | ( ~x64 & n638 ) ;
  assign n647 = ( n574 & ~n645 ) | ( n574 & n646 ) | ( ~n645 & n646 ) ;
  assign n648 = ( x65 & n644 ) | ( x65 & ~n647 ) | ( n644 & ~n647 ) ;
  assign n649 = ( x65 & n574 ) | ( x65 & n638 ) | ( n574 & n638 ) ;
  assign n650 = x65 | n574 ;
  assign n651 = ( ~n577 & n649 ) | ( ~n577 & n650 ) | ( n649 & n650 ) ;
  assign n652 = ( n577 & n649 ) | ( n577 & n650 ) | ( n649 & n650 ) ;
  assign n653 = ( n577 & n651 ) | ( n577 & ~n652 ) | ( n651 & ~n652 ) ;
  assign n654 = ( x66 & n648 ) | ( x66 & ~n653 ) | ( n648 & ~n653 ) ;
  assign n655 = ( x66 & n578 ) | ( x66 & n638 ) | ( n578 & n638 ) ;
  assign n656 = x66 | n578 ;
  assign n657 = ( ~n583 & n655 ) | ( ~n583 & n656 ) | ( n655 & n656 ) ;
  assign n658 = ( n583 & n655 ) | ( n583 & n656 ) | ( n655 & n656 ) ;
  assign n659 = ( n583 & n657 ) | ( n583 & ~n658 ) | ( n657 & ~n658 ) ;
  assign n660 = ( x67 & n654 ) | ( x67 & ~n659 ) | ( n654 & ~n659 ) ;
  assign n661 = ( x67 & n584 ) | ( x67 & n638 ) | ( n584 & n638 ) ;
  assign n662 = x67 | n584 ;
  assign n663 = ( ~n589 & n661 ) | ( ~n589 & n662 ) | ( n661 & n662 ) ;
  assign n664 = ( n589 & n661 ) | ( n589 & n662 ) | ( n661 & n662 ) ;
  assign n665 = ( n589 & n663 ) | ( n589 & ~n664 ) | ( n663 & ~n664 ) ;
  assign n666 = ( x68 & n660 ) | ( x68 & ~n665 ) | ( n660 & ~n665 ) ;
  assign n667 = ( x68 & n590 ) | ( x68 & ~n638 ) | ( n590 & ~n638 ) ;
  assign n668 = x68 & n590 ;
  assign n669 = ( ~n595 & n667 ) | ( ~n595 & n668 ) | ( n667 & n668 ) ;
  assign n670 = ( n595 & n667 ) | ( n595 & n668 ) | ( n667 & n668 ) ;
  assign n671 = ( n595 & n669 ) | ( n595 & ~n670 ) | ( n669 & ~n670 ) ;
  assign n672 = ( x69 & n666 ) | ( x69 & ~n671 ) | ( n666 & ~n671 ) ;
  assign n673 = ( x69 & n596 ) | ( x69 & ~n638 ) | ( n596 & ~n638 ) ;
  assign n674 = x69 & n596 ;
  assign n675 = ( ~n601 & n673 ) | ( ~n601 & n674 ) | ( n673 & n674 ) ;
  assign n676 = ( n601 & n673 ) | ( n601 & n674 ) | ( n673 & n674 ) ;
  assign n677 = ( n601 & n675 ) | ( n601 & ~n676 ) | ( n675 & ~n676 ) ;
  assign n678 = ( x70 & n672 ) | ( x70 & ~n677 ) | ( n672 & ~n677 ) ;
  assign n679 = ( x70 & n602 ) | ( x70 & ~n638 ) | ( n602 & ~n638 ) ;
  assign n680 = x70 & n602 ;
  assign n681 = ( ~n607 & n679 ) | ( ~n607 & n680 ) | ( n679 & n680 ) ;
  assign n682 = ( n607 & n679 ) | ( n607 & n680 ) | ( n679 & n680 ) ;
  assign n683 = ( n607 & n681 ) | ( n607 & ~n682 ) | ( n681 & ~n682 ) ;
  assign n684 = ( x71 & n678 ) | ( x71 & ~n683 ) | ( n678 & ~n683 ) ;
  assign n685 = ( x71 & n608 ) | ( x71 & ~n638 ) | ( n608 & ~n638 ) ;
  assign n686 = x71 & n608 ;
  assign n687 = ( ~n613 & n685 ) | ( ~n613 & n686 ) | ( n685 & n686 ) ;
  assign n688 = ( n613 & n685 ) | ( n613 & n686 ) | ( n685 & n686 ) ;
  assign n689 = ( n613 & n687 ) | ( n613 & ~n688 ) | ( n687 & ~n688 ) ;
  assign n690 = ( x72 & n684 ) | ( x72 & ~n689 ) | ( n684 & ~n689 ) ;
  assign n691 = ( x72 & n614 ) | ( x72 & ~n638 ) | ( n614 & ~n638 ) ;
  assign n692 = x72 & n614 ;
  assign n693 = ( ~n619 & n691 ) | ( ~n619 & n692 ) | ( n691 & n692 ) ;
  assign n694 = ( n619 & n691 ) | ( n619 & n692 ) | ( n691 & n692 ) ;
  assign n695 = ( n619 & n693 ) | ( n619 & ~n694 ) | ( n693 & ~n694 ) ;
  assign n696 = ( x73 & n690 ) | ( x73 & ~n695 ) | ( n690 & ~n695 ) ;
  assign n697 = ( x73 & n620 ) | ( x73 & ~n638 ) | ( n620 & ~n638 ) ;
  assign n698 = x73 & n620 ;
  assign n699 = ( ~n625 & n697 ) | ( ~n625 & n698 ) | ( n697 & n698 ) ;
  assign n700 = ( n625 & n697 ) | ( n625 & n698 ) | ( n697 & n698 ) ;
  assign n701 = ( n625 & n699 ) | ( n625 & ~n700 ) | ( n699 & ~n700 ) ;
  assign n702 = ( x74 & n696 ) | ( x74 & ~n701 ) | ( n696 & ~n701 ) ;
  assign n703 = ( x74 & n626 ) | ( x74 & ~n638 ) | ( n626 & ~n638 ) ;
  assign n704 = x74 & n626 ;
  assign n705 = ( ~n631 & n703 ) | ( ~n631 & n704 ) | ( n703 & n704 ) ;
  assign n706 = ( n631 & n703 ) | ( n631 & n704 ) | ( n703 & n704 ) ;
  assign n707 = ( n631 & n705 ) | ( n631 & ~n706 ) | ( n705 & ~n706 ) ;
  assign n708 = ( x75 & n702 ) | ( x75 & ~n707 ) | ( n702 & ~n707 ) ;
  assign n709 = ( x76 & n180 ) | ( x76 & n633 ) | ( n180 & n633 ) ;
  assign n710 = x76 | n633 ;
  assign n711 = ( n636 & n709 ) | ( n636 & ~n710 ) | ( n709 & ~n710 ) ;
  assign n712 = ( x76 & ~n643 ) | ( x76 & n708 ) | ( ~n643 & n708 ) ;
  assign n713 = ( x77 & ~n711 ) | ( x77 & n712 ) | ( ~n711 & n712 ) ;
  assign n714 = n179 | n713 ;
  assign n715 = ( x76 & n708 ) | ( x76 & n714 ) | ( n708 & n714 ) ;
  assign n716 = x76 | n708 ;
  assign n717 = ( ~n643 & n715 ) | ( ~n643 & n716 ) | ( n715 & n716 ) ;
  assign n718 = ( n643 & n715 ) | ( n643 & n716 ) | ( n715 & n716 ) ;
  assign n719 = ( n643 & n717 ) | ( n643 & ~n718 ) | ( n717 & ~n718 ) ;
  assign n720 = ~x49 & x64 ;
  assign n721 = ~x50 & n714 ;
  assign n722 = ( x50 & ~x64 ) | ( x50 & n714 ) | ( ~x64 & n714 ) ;
  assign n723 = ( n644 & ~n721 ) | ( n644 & n722 ) | ( ~n721 & n722 ) ;
  assign n724 = ( x65 & n720 ) | ( x65 & ~n723 ) | ( n720 & ~n723 ) ;
  assign n725 = ( x65 & n644 ) | ( x65 & n714 ) | ( n644 & n714 ) ;
  assign n726 = x65 | n644 ;
  assign n727 = ( ~n647 & n725 ) | ( ~n647 & n726 ) | ( n725 & n726 ) ;
  assign n728 = ( n647 & n725 ) | ( n647 & n726 ) | ( n725 & n726 ) ;
  assign n729 = ( n647 & n727 ) | ( n647 & ~n728 ) | ( n727 & ~n728 ) ;
  assign n730 = ( x66 & n724 ) | ( x66 & ~n729 ) | ( n724 & ~n729 ) ;
  assign n731 = ( x66 & n648 ) | ( x66 & n714 ) | ( n648 & n714 ) ;
  assign n732 = x66 | n648 ;
  assign n733 = ( ~n653 & n731 ) | ( ~n653 & n732 ) | ( n731 & n732 ) ;
  assign n734 = ( n653 & n731 ) | ( n653 & n732 ) | ( n731 & n732 ) ;
  assign n735 = ( n653 & n733 ) | ( n653 & ~n734 ) | ( n733 & ~n734 ) ;
  assign n736 = ( x67 & n730 ) | ( x67 & ~n735 ) | ( n730 & ~n735 ) ;
  assign n737 = ( x67 & n654 ) | ( x67 & n714 ) | ( n654 & n714 ) ;
  assign n738 = x67 | n654 ;
  assign n739 = ( ~n659 & n737 ) | ( ~n659 & n738 ) | ( n737 & n738 ) ;
  assign n740 = ( n659 & n737 ) | ( n659 & n738 ) | ( n737 & n738 ) ;
  assign n741 = ( n659 & n739 ) | ( n659 & ~n740 ) | ( n739 & ~n740 ) ;
  assign n742 = ( x68 & n736 ) | ( x68 & ~n741 ) | ( n736 & ~n741 ) ;
  assign n743 = ( x68 & n660 ) | ( x68 & ~n714 ) | ( n660 & ~n714 ) ;
  assign n744 = x68 & n660 ;
  assign n745 = ( ~n665 & n743 ) | ( ~n665 & n744 ) | ( n743 & n744 ) ;
  assign n746 = ( n665 & n743 ) | ( n665 & n744 ) | ( n743 & n744 ) ;
  assign n747 = ( n665 & n745 ) | ( n665 & ~n746 ) | ( n745 & ~n746 ) ;
  assign n748 = ( x69 & n742 ) | ( x69 & ~n747 ) | ( n742 & ~n747 ) ;
  assign n749 = ( x69 & n666 ) | ( x69 & ~n714 ) | ( n666 & ~n714 ) ;
  assign n750 = x69 & n666 ;
  assign n751 = ( ~n671 & n749 ) | ( ~n671 & n750 ) | ( n749 & n750 ) ;
  assign n752 = ( n671 & n749 ) | ( n671 & n750 ) | ( n749 & n750 ) ;
  assign n753 = ( n671 & n751 ) | ( n671 & ~n752 ) | ( n751 & ~n752 ) ;
  assign n754 = ( x70 & n748 ) | ( x70 & ~n753 ) | ( n748 & ~n753 ) ;
  assign n755 = ( x70 & n672 ) | ( x70 & ~n714 ) | ( n672 & ~n714 ) ;
  assign n756 = x70 & n672 ;
  assign n757 = ( ~n677 & n755 ) | ( ~n677 & n756 ) | ( n755 & n756 ) ;
  assign n758 = ( n677 & n755 ) | ( n677 & n756 ) | ( n755 & n756 ) ;
  assign n759 = ( n677 & n757 ) | ( n677 & ~n758 ) | ( n757 & ~n758 ) ;
  assign n760 = ( x71 & n754 ) | ( x71 & ~n759 ) | ( n754 & ~n759 ) ;
  assign n761 = ( x71 & n678 ) | ( x71 & ~n714 ) | ( n678 & ~n714 ) ;
  assign n762 = x71 & n678 ;
  assign n763 = ( ~n683 & n761 ) | ( ~n683 & n762 ) | ( n761 & n762 ) ;
  assign n764 = ( n683 & n761 ) | ( n683 & n762 ) | ( n761 & n762 ) ;
  assign n765 = ( n683 & n763 ) | ( n683 & ~n764 ) | ( n763 & ~n764 ) ;
  assign n766 = ( x72 & n760 ) | ( x72 & ~n765 ) | ( n760 & ~n765 ) ;
  assign n767 = ( x72 & n684 ) | ( x72 & ~n714 ) | ( n684 & ~n714 ) ;
  assign n768 = x72 & n684 ;
  assign n769 = ( ~n689 & n767 ) | ( ~n689 & n768 ) | ( n767 & n768 ) ;
  assign n770 = ( n689 & n767 ) | ( n689 & n768 ) | ( n767 & n768 ) ;
  assign n771 = ( n689 & n769 ) | ( n689 & ~n770 ) | ( n769 & ~n770 ) ;
  assign n772 = ( x73 & n766 ) | ( x73 & ~n771 ) | ( n766 & ~n771 ) ;
  assign n773 = ( x73 & n690 ) | ( x73 & ~n714 ) | ( n690 & ~n714 ) ;
  assign n774 = x73 & n690 ;
  assign n775 = ( ~n695 & n773 ) | ( ~n695 & n774 ) | ( n773 & n774 ) ;
  assign n776 = ( n695 & n773 ) | ( n695 & n774 ) | ( n773 & n774 ) ;
  assign n777 = ( n695 & n775 ) | ( n695 & ~n776 ) | ( n775 & ~n776 ) ;
  assign n778 = ( x74 & n772 ) | ( x74 & ~n777 ) | ( n772 & ~n777 ) ;
  assign n779 = ( x74 & n696 ) | ( x74 & ~n714 ) | ( n696 & ~n714 ) ;
  assign n780 = x74 & n696 ;
  assign n781 = ( ~n701 & n779 ) | ( ~n701 & n780 ) | ( n779 & n780 ) ;
  assign n782 = ( n701 & n779 ) | ( n701 & n780 ) | ( n779 & n780 ) ;
  assign n783 = ( n701 & n781 ) | ( n701 & ~n782 ) | ( n781 & ~n782 ) ;
  assign n784 = ( x75 & n778 ) | ( x75 & ~n783 ) | ( n778 & ~n783 ) ;
  assign n785 = ( x75 & n702 ) | ( x75 & ~n714 ) | ( n702 & ~n714 ) ;
  assign n786 = x75 & n702 ;
  assign n787 = ( ~n707 & n785 ) | ( ~n707 & n786 ) | ( n785 & n786 ) ;
  assign n788 = ( n707 & n785 ) | ( n707 & n786 ) | ( n785 & n786 ) ;
  assign n789 = ( n707 & n787 ) | ( n707 & ~n788 ) | ( n787 & ~n788 ) ;
  assign n790 = ( x76 & n784 ) | ( x76 & ~n789 ) | ( n784 & ~n789 ) ;
  assign n791 = ( n178 & n179 ) | ( n178 & ~n711 ) | ( n179 & ~n711 ) ;
  assign n792 = ( x77 & ~n719 ) | ( x77 & n790 ) | ( ~n719 & n790 ) ;
  assign n793 = n791 | n792 ;
  assign n794 = ( ~x77 & n179 ) | ( ~x77 & n712 ) | ( n179 & n712 ) ;
  assign n795 = ( ~x77 & n711 ) | ( ~x77 & n712 ) | ( n711 & n712 ) ;
  assign n796 = ~n794 & n795 ;
  assign n797 = n793 & ~n796 ;
  assign n798 = ( x77 & n790 ) | ( x77 & ~n797 ) | ( n790 & ~n797 ) ;
  assign n799 = x77 & n790 ;
  assign n800 = ( ~n719 & n798 ) | ( ~n719 & n799 ) | ( n798 & n799 ) ;
  assign n801 = ( n719 & n798 ) | ( n719 & n799 ) | ( n798 & n799 ) ;
  assign n802 = ( n719 & n800 ) | ( n719 & ~n801 ) | ( n800 & ~n801 ) ;
  assign n803 = ~x48 & x64 ;
  assign n804 = x49 & n797 ;
  assign n805 = ( x49 & x64 ) | ( x49 & ~n797 ) | ( x64 & ~n797 ) ;
  assign n806 = x49 & x64 ;
  assign n807 = ( n804 & n805 ) | ( n804 & ~n806 ) | ( n805 & ~n806 ) ;
  assign n808 = ( x65 & n803 ) | ( x65 & ~n807 ) | ( n803 & ~n807 ) ;
  assign n809 = ( x65 & n720 ) | ( x65 & n797 ) | ( n720 & n797 ) ;
  assign n810 = x65 | n720 ;
  assign n811 = ( ~n723 & n809 ) | ( ~n723 & n810 ) | ( n809 & n810 ) ;
  assign n812 = ( n723 & n809 ) | ( n723 & n810 ) | ( n809 & n810 ) ;
  assign n813 = ( n723 & n811 ) | ( n723 & ~n812 ) | ( n811 & ~n812 ) ;
  assign n814 = ( x66 & n808 ) | ( x66 & ~n813 ) | ( n808 & ~n813 ) ;
  assign n815 = ( x66 & n724 ) | ( x66 & n797 ) | ( n724 & n797 ) ;
  assign n816 = x66 | n724 ;
  assign n817 = ( ~n729 & n815 ) | ( ~n729 & n816 ) | ( n815 & n816 ) ;
  assign n818 = ( n729 & n815 ) | ( n729 & n816 ) | ( n815 & n816 ) ;
  assign n819 = ( n729 & n817 ) | ( n729 & ~n818 ) | ( n817 & ~n818 ) ;
  assign n820 = ( x67 & n814 ) | ( x67 & ~n819 ) | ( n814 & ~n819 ) ;
  assign n821 = ( x67 & n730 ) | ( x67 & ~n797 ) | ( n730 & ~n797 ) ;
  assign n822 = x67 & n730 ;
  assign n823 = ( ~n735 & n821 ) | ( ~n735 & n822 ) | ( n821 & n822 ) ;
  assign n824 = ( n735 & n821 ) | ( n735 & n822 ) | ( n821 & n822 ) ;
  assign n825 = ( n735 & n823 ) | ( n735 & ~n824 ) | ( n823 & ~n824 ) ;
  assign n826 = ( x68 & n820 ) | ( x68 & ~n825 ) | ( n820 & ~n825 ) ;
  assign n827 = ( x68 & n736 ) | ( x68 & ~n797 ) | ( n736 & ~n797 ) ;
  assign n828 = x68 & n736 ;
  assign n829 = ( ~n741 & n827 ) | ( ~n741 & n828 ) | ( n827 & n828 ) ;
  assign n830 = ( n741 & n827 ) | ( n741 & n828 ) | ( n827 & n828 ) ;
  assign n831 = ( n741 & n829 ) | ( n741 & ~n830 ) | ( n829 & ~n830 ) ;
  assign n832 = ( x69 & n826 ) | ( x69 & ~n831 ) | ( n826 & ~n831 ) ;
  assign n833 = ( x69 & n742 ) | ( x69 & ~n797 ) | ( n742 & ~n797 ) ;
  assign n834 = x69 & n742 ;
  assign n835 = ( ~n747 & n833 ) | ( ~n747 & n834 ) | ( n833 & n834 ) ;
  assign n836 = ( n747 & n833 ) | ( n747 & n834 ) | ( n833 & n834 ) ;
  assign n837 = ( n747 & n835 ) | ( n747 & ~n836 ) | ( n835 & ~n836 ) ;
  assign n838 = ( x70 & n832 ) | ( x70 & ~n837 ) | ( n832 & ~n837 ) ;
  assign n839 = ( x70 & n748 ) | ( x70 & ~n797 ) | ( n748 & ~n797 ) ;
  assign n840 = x70 & n748 ;
  assign n841 = ( ~n753 & n839 ) | ( ~n753 & n840 ) | ( n839 & n840 ) ;
  assign n842 = ( n753 & n839 ) | ( n753 & n840 ) | ( n839 & n840 ) ;
  assign n843 = ( n753 & n841 ) | ( n753 & ~n842 ) | ( n841 & ~n842 ) ;
  assign n844 = ( x71 & n838 ) | ( x71 & ~n843 ) | ( n838 & ~n843 ) ;
  assign n845 = ( x71 & n754 ) | ( x71 & ~n797 ) | ( n754 & ~n797 ) ;
  assign n846 = x71 & n754 ;
  assign n847 = ( ~n759 & n845 ) | ( ~n759 & n846 ) | ( n845 & n846 ) ;
  assign n848 = ( n759 & n845 ) | ( n759 & n846 ) | ( n845 & n846 ) ;
  assign n849 = ( n759 & n847 ) | ( n759 & ~n848 ) | ( n847 & ~n848 ) ;
  assign n850 = ( x72 & n844 ) | ( x72 & ~n849 ) | ( n844 & ~n849 ) ;
  assign n851 = ( x72 & n760 ) | ( x72 & ~n797 ) | ( n760 & ~n797 ) ;
  assign n852 = x72 & n760 ;
  assign n853 = ( ~n765 & n851 ) | ( ~n765 & n852 ) | ( n851 & n852 ) ;
  assign n854 = ( n765 & n851 ) | ( n765 & n852 ) | ( n851 & n852 ) ;
  assign n855 = ( n765 & n853 ) | ( n765 & ~n854 ) | ( n853 & ~n854 ) ;
  assign n856 = ( x73 & n850 ) | ( x73 & ~n855 ) | ( n850 & ~n855 ) ;
  assign n857 = ( x73 & n766 ) | ( x73 & ~n797 ) | ( n766 & ~n797 ) ;
  assign n858 = x73 & n766 ;
  assign n859 = ( ~n771 & n857 ) | ( ~n771 & n858 ) | ( n857 & n858 ) ;
  assign n860 = ( n771 & n857 ) | ( n771 & n858 ) | ( n857 & n858 ) ;
  assign n861 = ( n771 & n859 ) | ( n771 & ~n860 ) | ( n859 & ~n860 ) ;
  assign n862 = ( x74 & n856 ) | ( x74 & ~n861 ) | ( n856 & ~n861 ) ;
  assign n863 = ( x74 & n772 ) | ( x74 & ~n797 ) | ( n772 & ~n797 ) ;
  assign n864 = x74 & n772 ;
  assign n865 = ( ~n777 & n863 ) | ( ~n777 & n864 ) | ( n863 & n864 ) ;
  assign n866 = ( n777 & n863 ) | ( n777 & n864 ) | ( n863 & n864 ) ;
  assign n867 = ( n777 & n865 ) | ( n777 & ~n866 ) | ( n865 & ~n866 ) ;
  assign n868 = ( x75 & n862 ) | ( x75 & ~n867 ) | ( n862 & ~n867 ) ;
  assign n869 = ( x75 & n778 ) | ( x75 & ~n797 ) | ( n778 & ~n797 ) ;
  assign n870 = x75 & n778 ;
  assign n871 = ( ~n783 & n869 ) | ( ~n783 & n870 ) | ( n869 & n870 ) ;
  assign n872 = ( n783 & n869 ) | ( n783 & n870 ) | ( n869 & n870 ) ;
  assign n873 = ( n783 & n871 ) | ( n783 & ~n872 ) | ( n871 & ~n872 ) ;
  assign n874 = ( x76 & n868 ) | ( x76 & ~n873 ) | ( n868 & ~n873 ) ;
  assign n875 = ( x76 & n784 ) | ( x76 & ~n797 ) | ( n784 & ~n797 ) ;
  assign n876 = x76 & n784 ;
  assign n877 = ( ~n789 & n875 ) | ( ~n789 & n876 ) | ( n875 & n876 ) ;
  assign n878 = ( n789 & n875 ) | ( n789 & n876 ) | ( n875 & n876 ) ;
  assign n879 = ( n789 & n877 ) | ( n789 & ~n878 ) | ( n877 & ~n878 ) ;
  assign n880 = ( x77 & n874 ) | ( x77 & ~n879 ) | ( n874 & ~n879 ) ;
  assign n881 = ( n179 & n389 ) | ( n179 & n636 ) | ( n389 & n636 ) ;
  assign n882 = ( n389 & n793 ) | ( n389 & n881 ) | ( n793 & n881 ) ;
  assign n883 = ( x78 & ~n802 ) | ( x78 & n880 ) | ( ~n802 & n880 ) ;
  assign n884 = ( x79 & ~n882 ) | ( x79 & n883 ) | ( ~n882 & n883 ) ;
  assign n885 = n177 | n884 ;
  assign n886 = ( x78 & n880 ) | ( x78 & n885 ) | ( n880 & n885 ) ;
  assign n887 = x78 | n880 ;
  assign n888 = ( ~n802 & n886 ) | ( ~n802 & n887 ) | ( n886 & n887 ) ;
  assign n889 = ( n802 & n886 ) | ( n802 & n887 ) | ( n886 & n887 ) ;
  assign n890 = ( n802 & n888 ) | ( n802 & ~n889 ) | ( n888 & ~n889 ) ;
  assign n891 = ~x47 & x64 ;
  assign n892 = ~x48 & n885 ;
  assign n893 = ( x48 & ~x64 ) | ( x48 & n885 ) | ( ~x64 & n885 ) ;
  assign n894 = ( n803 & ~n892 ) | ( n803 & n893 ) | ( ~n892 & n893 ) ;
  assign n895 = ( x65 & n891 ) | ( x65 & ~n894 ) | ( n891 & ~n894 ) ;
  assign n896 = ( x65 & n803 ) | ( x65 & n885 ) | ( n803 & n885 ) ;
  assign n897 = x65 | n803 ;
  assign n898 = ( ~n807 & n896 ) | ( ~n807 & n897 ) | ( n896 & n897 ) ;
  assign n899 = ( n807 & n896 ) | ( n807 & n897 ) | ( n896 & n897 ) ;
  assign n900 = ( n807 & n898 ) | ( n807 & ~n899 ) | ( n898 & ~n899 ) ;
  assign n901 = ( x66 & n895 ) | ( x66 & ~n900 ) | ( n895 & ~n900 ) ;
  assign n902 = ( x66 & n808 ) | ( x66 & n885 ) | ( n808 & n885 ) ;
  assign n903 = x66 | n808 ;
  assign n904 = ( ~n813 & n902 ) | ( ~n813 & n903 ) | ( n902 & n903 ) ;
  assign n905 = ( n813 & n902 ) | ( n813 & n903 ) | ( n902 & n903 ) ;
  assign n906 = ( n813 & n904 ) | ( n813 & ~n905 ) | ( n904 & ~n905 ) ;
  assign n907 = ( x67 & n901 ) | ( x67 & ~n906 ) | ( n901 & ~n906 ) ;
  assign n908 = ( x67 & n814 ) | ( x67 & n885 ) | ( n814 & n885 ) ;
  assign n909 = x67 | n814 ;
  assign n910 = ( ~n819 & n908 ) | ( ~n819 & n909 ) | ( n908 & n909 ) ;
  assign n911 = ( n819 & n908 ) | ( n819 & n909 ) | ( n908 & n909 ) ;
  assign n912 = ( n819 & n910 ) | ( n819 & ~n911 ) | ( n910 & ~n911 ) ;
  assign n913 = ( x68 & n907 ) | ( x68 & ~n912 ) | ( n907 & ~n912 ) ;
  assign n914 = ( x68 & n820 ) | ( x68 & ~n885 ) | ( n820 & ~n885 ) ;
  assign n915 = x68 & n820 ;
  assign n916 = ( ~n825 & n914 ) | ( ~n825 & n915 ) | ( n914 & n915 ) ;
  assign n917 = ( n825 & n914 ) | ( n825 & n915 ) | ( n914 & n915 ) ;
  assign n918 = ( n825 & n916 ) | ( n825 & ~n917 ) | ( n916 & ~n917 ) ;
  assign n919 = ( x69 & n913 ) | ( x69 & ~n918 ) | ( n913 & ~n918 ) ;
  assign n920 = ( x69 & n826 ) | ( x69 & ~n885 ) | ( n826 & ~n885 ) ;
  assign n921 = x69 & n826 ;
  assign n922 = ( ~n831 & n920 ) | ( ~n831 & n921 ) | ( n920 & n921 ) ;
  assign n923 = ( n831 & n920 ) | ( n831 & n921 ) | ( n920 & n921 ) ;
  assign n924 = ( n831 & n922 ) | ( n831 & ~n923 ) | ( n922 & ~n923 ) ;
  assign n925 = ( x70 & n919 ) | ( x70 & ~n924 ) | ( n919 & ~n924 ) ;
  assign n926 = ( x70 & n832 ) | ( x70 & ~n885 ) | ( n832 & ~n885 ) ;
  assign n927 = x70 & n832 ;
  assign n928 = ( ~n837 & n926 ) | ( ~n837 & n927 ) | ( n926 & n927 ) ;
  assign n929 = ( n837 & n926 ) | ( n837 & n927 ) | ( n926 & n927 ) ;
  assign n930 = ( n837 & n928 ) | ( n837 & ~n929 ) | ( n928 & ~n929 ) ;
  assign n931 = ( x71 & n925 ) | ( x71 & ~n930 ) | ( n925 & ~n930 ) ;
  assign n932 = ( x71 & n838 ) | ( x71 & ~n885 ) | ( n838 & ~n885 ) ;
  assign n933 = x71 & n838 ;
  assign n934 = ( ~n843 & n932 ) | ( ~n843 & n933 ) | ( n932 & n933 ) ;
  assign n935 = ( n843 & n932 ) | ( n843 & n933 ) | ( n932 & n933 ) ;
  assign n936 = ( n843 & n934 ) | ( n843 & ~n935 ) | ( n934 & ~n935 ) ;
  assign n937 = ( x72 & n931 ) | ( x72 & ~n936 ) | ( n931 & ~n936 ) ;
  assign n938 = ( x72 & n844 ) | ( x72 & ~n885 ) | ( n844 & ~n885 ) ;
  assign n939 = x72 & n844 ;
  assign n940 = ( ~n849 & n938 ) | ( ~n849 & n939 ) | ( n938 & n939 ) ;
  assign n941 = ( n849 & n938 ) | ( n849 & n939 ) | ( n938 & n939 ) ;
  assign n942 = ( n849 & n940 ) | ( n849 & ~n941 ) | ( n940 & ~n941 ) ;
  assign n943 = ( x73 & n937 ) | ( x73 & ~n942 ) | ( n937 & ~n942 ) ;
  assign n944 = ( x73 & n850 ) | ( x73 & ~n885 ) | ( n850 & ~n885 ) ;
  assign n945 = x73 & n850 ;
  assign n946 = ( ~n855 & n944 ) | ( ~n855 & n945 ) | ( n944 & n945 ) ;
  assign n947 = ( n855 & n944 ) | ( n855 & n945 ) | ( n944 & n945 ) ;
  assign n948 = ( n855 & n946 ) | ( n855 & ~n947 ) | ( n946 & ~n947 ) ;
  assign n949 = ( x74 & n943 ) | ( x74 & ~n948 ) | ( n943 & ~n948 ) ;
  assign n950 = ( x74 & n856 ) | ( x74 & ~n885 ) | ( n856 & ~n885 ) ;
  assign n951 = x74 & n856 ;
  assign n952 = ( ~n861 & n950 ) | ( ~n861 & n951 ) | ( n950 & n951 ) ;
  assign n953 = ( n861 & n950 ) | ( n861 & n951 ) | ( n950 & n951 ) ;
  assign n954 = ( n861 & n952 ) | ( n861 & ~n953 ) | ( n952 & ~n953 ) ;
  assign n955 = ( x75 & n949 ) | ( x75 & ~n954 ) | ( n949 & ~n954 ) ;
  assign n956 = ( x75 & n862 ) | ( x75 & ~n885 ) | ( n862 & ~n885 ) ;
  assign n957 = x75 & n862 ;
  assign n958 = ( ~n867 & n956 ) | ( ~n867 & n957 ) | ( n956 & n957 ) ;
  assign n959 = ( n867 & n956 ) | ( n867 & n957 ) | ( n956 & n957 ) ;
  assign n960 = ( n867 & n958 ) | ( n867 & ~n959 ) | ( n958 & ~n959 ) ;
  assign n961 = ( x76 & n955 ) | ( x76 & ~n960 ) | ( n955 & ~n960 ) ;
  assign n962 = ( x76 & n868 ) | ( x76 & ~n885 ) | ( n868 & ~n885 ) ;
  assign n963 = x76 & n868 ;
  assign n964 = ( ~n873 & n962 ) | ( ~n873 & n963 ) | ( n962 & n963 ) ;
  assign n965 = ( n873 & n962 ) | ( n873 & n963 ) | ( n962 & n963 ) ;
  assign n966 = ( n873 & n964 ) | ( n873 & ~n965 ) | ( n964 & ~n965 ) ;
  assign n967 = ( x77 & n961 ) | ( x77 & ~n966 ) | ( n961 & ~n966 ) ;
  assign n968 = ( x77 & n874 ) | ( x77 & ~n885 ) | ( n874 & ~n885 ) ;
  assign n969 = x77 & n874 ;
  assign n970 = ( ~n879 & n968 ) | ( ~n879 & n969 ) | ( n968 & n969 ) ;
  assign n971 = ( n879 & n968 ) | ( n879 & n969 ) | ( n968 & n969 ) ;
  assign n972 = ( n879 & n970 ) | ( n879 & ~n971 ) | ( n970 & ~n971 ) ;
  assign n973 = ( x78 & n967 ) | ( x78 & ~n972 ) | ( n967 & ~n972 ) ;
  assign n974 = ( x79 & n177 ) | ( x79 & n883 ) | ( n177 & n883 ) ;
  assign n975 = x79 | n883 ;
  assign n976 = ( n882 & n974 ) | ( n882 & ~n975 ) | ( n974 & ~n975 ) ;
  assign n977 = ( x79 & ~n890 ) | ( x79 & n973 ) | ( ~n890 & n973 ) ;
  assign n978 = ( x80 & ~n976 ) | ( x80 & n977 ) | ( ~n976 & n977 ) ;
  assign n979 = n176 | n978 ;
  assign n980 = ( x79 & n973 ) | ( x79 & n979 ) | ( n973 & n979 ) ;
  assign n981 = x79 | n973 ;
  assign n982 = ( ~n890 & n980 ) | ( ~n890 & n981 ) | ( n980 & n981 ) ;
  assign n983 = ( n890 & n980 ) | ( n890 & n981 ) | ( n980 & n981 ) ;
  assign n984 = ( n890 & n982 ) | ( n890 & ~n983 ) | ( n982 & ~n983 ) ;
  assign n985 = ~x46 & x64 ;
  assign n986 = ~x47 & n979 ;
  assign n987 = ( x47 & ~x64 ) | ( x47 & n979 ) | ( ~x64 & n979 ) ;
  assign n988 = ( n891 & ~n986 ) | ( n891 & n987 ) | ( ~n986 & n987 ) ;
  assign n989 = ( x65 & n985 ) | ( x65 & ~n988 ) | ( n985 & ~n988 ) ;
  assign n990 = ( x65 & n891 ) | ( x65 & n979 ) | ( n891 & n979 ) ;
  assign n991 = x65 | n891 ;
  assign n992 = ( ~n894 & n990 ) | ( ~n894 & n991 ) | ( n990 & n991 ) ;
  assign n993 = ( n894 & n990 ) | ( n894 & n991 ) | ( n990 & n991 ) ;
  assign n994 = ( n894 & n992 ) | ( n894 & ~n993 ) | ( n992 & ~n993 ) ;
  assign n995 = ( x66 & n989 ) | ( x66 & ~n994 ) | ( n989 & ~n994 ) ;
  assign n996 = ( x66 & n895 ) | ( x66 & n979 ) | ( n895 & n979 ) ;
  assign n997 = x66 | n895 ;
  assign n998 = ( ~n900 & n996 ) | ( ~n900 & n997 ) | ( n996 & n997 ) ;
  assign n999 = ( n900 & n996 ) | ( n900 & n997 ) | ( n996 & n997 ) ;
  assign n1000 = ( n900 & n998 ) | ( n900 & ~n999 ) | ( n998 & ~n999 ) ;
  assign n1001 = ( x67 & n995 ) | ( x67 & ~n1000 ) | ( n995 & ~n1000 ) ;
  assign n1002 = ( x67 & n901 ) | ( x67 & n979 ) | ( n901 & n979 ) ;
  assign n1003 = x67 | n901 ;
  assign n1004 = ( ~n906 & n1002 ) | ( ~n906 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1005 = ( n906 & n1002 ) | ( n906 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1006 = ( n906 & n1004 ) | ( n906 & ~n1005 ) | ( n1004 & ~n1005 ) ;
  assign n1007 = ( x68 & n1001 ) | ( x68 & ~n1006 ) | ( n1001 & ~n1006 ) ;
  assign n1008 = ( x68 & n907 ) | ( x68 & n979 ) | ( n907 & n979 ) ;
  assign n1009 = x68 | n907 ;
  assign n1010 = ( ~n912 & n1008 ) | ( ~n912 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1011 = ( n912 & n1008 ) | ( n912 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1012 = ( n912 & n1010 ) | ( n912 & ~n1011 ) | ( n1010 & ~n1011 ) ;
  assign n1013 = ( x69 & n1007 ) | ( x69 & ~n1012 ) | ( n1007 & ~n1012 ) ;
  assign n1014 = ( x69 & n913 ) | ( x69 & ~n979 ) | ( n913 & ~n979 ) ;
  assign n1015 = x69 & n913 ;
  assign n1016 = ( ~n918 & n1014 ) | ( ~n918 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = ( n918 & n1014 ) | ( n918 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1018 = ( n918 & n1016 ) | ( n918 & ~n1017 ) | ( n1016 & ~n1017 ) ;
  assign n1019 = ( x70 & n1013 ) | ( x70 & ~n1018 ) | ( n1013 & ~n1018 ) ;
  assign n1020 = ( x70 & n919 ) | ( x70 & ~n979 ) | ( n919 & ~n979 ) ;
  assign n1021 = x70 & n919 ;
  assign n1022 = ( ~n924 & n1020 ) | ( ~n924 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1023 = ( n924 & n1020 ) | ( n924 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1024 = ( n924 & n1022 ) | ( n924 & ~n1023 ) | ( n1022 & ~n1023 ) ;
  assign n1025 = ( x71 & n1019 ) | ( x71 & ~n1024 ) | ( n1019 & ~n1024 ) ;
  assign n1026 = ( x71 & n925 ) | ( x71 & ~n979 ) | ( n925 & ~n979 ) ;
  assign n1027 = x71 & n925 ;
  assign n1028 = ( ~n930 & n1026 ) | ( ~n930 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1029 = ( n930 & n1026 ) | ( n930 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1030 = ( n930 & n1028 ) | ( n930 & ~n1029 ) | ( n1028 & ~n1029 ) ;
  assign n1031 = ( x72 & n1025 ) | ( x72 & ~n1030 ) | ( n1025 & ~n1030 ) ;
  assign n1032 = ( x72 & n931 ) | ( x72 & ~n979 ) | ( n931 & ~n979 ) ;
  assign n1033 = x72 & n931 ;
  assign n1034 = ( ~n936 & n1032 ) | ( ~n936 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1035 = ( n936 & n1032 ) | ( n936 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1036 = ( n936 & n1034 ) | ( n936 & ~n1035 ) | ( n1034 & ~n1035 ) ;
  assign n1037 = ( x73 & n1031 ) | ( x73 & ~n1036 ) | ( n1031 & ~n1036 ) ;
  assign n1038 = ( x73 & n937 ) | ( x73 & ~n979 ) | ( n937 & ~n979 ) ;
  assign n1039 = x73 & n937 ;
  assign n1040 = ( ~n942 & n1038 ) | ( ~n942 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1041 = ( n942 & n1038 ) | ( n942 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1042 = ( n942 & n1040 ) | ( n942 & ~n1041 ) | ( n1040 & ~n1041 ) ;
  assign n1043 = ( x74 & n1037 ) | ( x74 & ~n1042 ) | ( n1037 & ~n1042 ) ;
  assign n1044 = ( x74 & n943 ) | ( x74 & ~n979 ) | ( n943 & ~n979 ) ;
  assign n1045 = x74 & n943 ;
  assign n1046 = ( ~n948 & n1044 ) | ( ~n948 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1047 = ( n948 & n1044 ) | ( n948 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1048 = ( n948 & n1046 ) | ( n948 & ~n1047 ) | ( n1046 & ~n1047 ) ;
  assign n1049 = ( x75 & n1043 ) | ( x75 & ~n1048 ) | ( n1043 & ~n1048 ) ;
  assign n1050 = ( x75 & n949 ) | ( x75 & ~n979 ) | ( n949 & ~n979 ) ;
  assign n1051 = x75 & n949 ;
  assign n1052 = ( ~n954 & n1050 ) | ( ~n954 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1053 = ( n954 & n1050 ) | ( n954 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1054 = ( n954 & n1052 ) | ( n954 & ~n1053 ) | ( n1052 & ~n1053 ) ;
  assign n1055 = ( x76 & n1049 ) | ( x76 & ~n1054 ) | ( n1049 & ~n1054 ) ;
  assign n1056 = ( x76 & n955 ) | ( x76 & ~n979 ) | ( n955 & ~n979 ) ;
  assign n1057 = x76 & n955 ;
  assign n1058 = ( ~n960 & n1056 ) | ( ~n960 & n1057 ) | ( n1056 & n1057 ) ;
  assign n1059 = ( n960 & n1056 ) | ( n960 & n1057 ) | ( n1056 & n1057 ) ;
  assign n1060 = ( n960 & n1058 ) | ( n960 & ~n1059 ) | ( n1058 & ~n1059 ) ;
  assign n1061 = ( x77 & n1055 ) | ( x77 & ~n1060 ) | ( n1055 & ~n1060 ) ;
  assign n1062 = ( x77 & n961 ) | ( x77 & ~n979 ) | ( n961 & ~n979 ) ;
  assign n1063 = x77 & n961 ;
  assign n1064 = ( ~n966 & n1062 ) | ( ~n966 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1065 = ( n966 & n1062 ) | ( n966 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1066 = ( n966 & n1064 ) | ( n966 & ~n1065 ) | ( n1064 & ~n1065 ) ;
  assign n1067 = ( x78 & n1061 ) | ( x78 & ~n1066 ) | ( n1061 & ~n1066 ) ;
  assign n1068 = ( x78 & n967 ) | ( x78 & ~n979 ) | ( n967 & ~n979 ) ;
  assign n1069 = x78 & n967 ;
  assign n1070 = ( ~n972 & n1068 ) | ( ~n972 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1071 = ( n972 & n1068 ) | ( n972 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1072 = ( n972 & n1070 ) | ( n972 & ~n1071 ) | ( n1070 & ~n1071 ) ;
  assign n1073 = ( x79 & n1067 ) | ( x79 & ~n1072 ) | ( n1067 & ~n1072 ) ;
  assign n1074 = ( n175 & n176 ) | ( n175 & ~n976 ) | ( n176 & ~n976 ) ;
  assign n1075 = ( x80 & ~n984 ) | ( x80 & n1073 ) | ( ~n984 & n1073 ) ;
  assign n1076 = ( ~x80 & x81 ) | ( ~x80 & n977 ) | ( x81 & n977 ) ;
  assign n1077 = ( ~x80 & n976 ) | ( ~x80 & n977 ) | ( n976 & n977 ) ;
  assign n1078 = ~n1076 & n1077 ;
  assign n1079 = ~n1074 & n1078 ;
  assign n1080 = ( n1074 & n1075 ) | ( n1074 & ~n1079 ) | ( n1075 & ~n1079 ) ;
  assign n1081 = ( x80 & n1073 ) | ( x80 & n1080 ) | ( n1073 & n1080 ) ;
  assign n1082 = x80 | n1073 ;
  assign n1083 = ( ~n984 & n1081 ) | ( ~n984 & n1082 ) | ( n1081 & n1082 ) ;
  assign n1084 = ( n984 & n1081 ) | ( n984 & n1082 ) | ( n1081 & n1082 ) ;
  assign n1085 = ( n984 & n1083 ) | ( n984 & ~n1084 ) | ( n1083 & ~n1084 ) ;
  assign n1086 = ~x45 & x64 ;
  assign n1087 = ~x46 & n1080 ;
  assign n1088 = ( x46 & ~x64 ) | ( x46 & n1080 ) | ( ~x64 & n1080 ) ;
  assign n1089 = ( n985 & ~n1087 ) | ( n985 & n1088 ) | ( ~n1087 & n1088 ) ;
  assign n1090 = ( x65 & n1086 ) | ( x65 & ~n1089 ) | ( n1086 & ~n1089 ) ;
  assign n1091 = ( x65 & n985 ) | ( x65 & n1080 ) | ( n985 & n1080 ) ;
  assign n1092 = x65 | n985 ;
  assign n1093 = ( ~n988 & n1091 ) | ( ~n988 & n1092 ) | ( n1091 & n1092 ) ;
  assign n1094 = ( n988 & n1091 ) | ( n988 & n1092 ) | ( n1091 & n1092 ) ;
  assign n1095 = ( n988 & n1093 ) | ( n988 & ~n1094 ) | ( n1093 & ~n1094 ) ;
  assign n1096 = ( x66 & n1090 ) | ( x66 & ~n1095 ) | ( n1090 & ~n1095 ) ;
  assign n1097 = ( x66 & n989 ) | ( x66 & n1080 ) | ( n989 & n1080 ) ;
  assign n1098 = x66 | n989 ;
  assign n1099 = ( ~n994 & n1097 ) | ( ~n994 & n1098 ) | ( n1097 & n1098 ) ;
  assign n1100 = ( n994 & n1097 ) | ( n994 & n1098 ) | ( n1097 & n1098 ) ;
  assign n1101 = ( n994 & n1099 ) | ( n994 & ~n1100 ) | ( n1099 & ~n1100 ) ;
  assign n1102 = ( x67 & n1096 ) | ( x67 & ~n1101 ) | ( n1096 & ~n1101 ) ;
  assign n1103 = ( x67 & n995 ) | ( x67 & n1080 ) | ( n995 & n1080 ) ;
  assign n1104 = x67 | n995 ;
  assign n1105 = ( ~n1000 & n1103 ) | ( ~n1000 & n1104 ) | ( n1103 & n1104 ) ;
  assign n1106 = ( n1000 & n1103 ) | ( n1000 & n1104 ) | ( n1103 & n1104 ) ;
  assign n1107 = ( n1000 & n1105 ) | ( n1000 & ~n1106 ) | ( n1105 & ~n1106 ) ;
  assign n1108 = ( x68 & n1102 ) | ( x68 & ~n1107 ) | ( n1102 & ~n1107 ) ;
  assign n1109 = ( x68 & n1001 ) | ( x68 & ~n1080 ) | ( n1001 & ~n1080 ) ;
  assign n1110 = x68 & n1001 ;
  assign n1111 = ( ~n1006 & n1109 ) | ( ~n1006 & n1110 ) | ( n1109 & n1110 ) ;
  assign n1112 = ( n1006 & n1109 ) | ( n1006 & n1110 ) | ( n1109 & n1110 ) ;
  assign n1113 = ( n1006 & n1111 ) | ( n1006 & ~n1112 ) | ( n1111 & ~n1112 ) ;
  assign n1114 = ( x69 & n1108 ) | ( x69 & ~n1113 ) | ( n1108 & ~n1113 ) ;
  assign n1115 = ( x69 & n1007 ) | ( x69 & ~n1080 ) | ( n1007 & ~n1080 ) ;
  assign n1116 = x69 & n1007 ;
  assign n1117 = ( ~n1012 & n1115 ) | ( ~n1012 & n1116 ) | ( n1115 & n1116 ) ;
  assign n1118 = ( n1012 & n1115 ) | ( n1012 & n1116 ) | ( n1115 & n1116 ) ;
  assign n1119 = ( n1012 & n1117 ) | ( n1012 & ~n1118 ) | ( n1117 & ~n1118 ) ;
  assign n1120 = ( x70 & n1114 ) | ( x70 & ~n1119 ) | ( n1114 & ~n1119 ) ;
  assign n1121 = ( x70 & n1013 ) | ( x70 & ~n1080 ) | ( n1013 & ~n1080 ) ;
  assign n1122 = x70 & n1013 ;
  assign n1123 = ( ~n1018 & n1121 ) | ( ~n1018 & n1122 ) | ( n1121 & n1122 ) ;
  assign n1124 = ( n1018 & n1121 ) | ( n1018 & n1122 ) | ( n1121 & n1122 ) ;
  assign n1125 = ( n1018 & n1123 ) | ( n1018 & ~n1124 ) | ( n1123 & ~n1124 ) ;
  assign n1126 = ( x71 & n1120 ) | ( x71 & ~n1125 ) | ( n1120 & ~n1125 ) ;
  assign n1127 = ( x71 & n1019 ) | ( x71 & ~n1080 ) | ( n1019 & ~n1080 ) ;
  assign n1128 = x71 & n1019 ;
  assign n1129 = ( ~n1024 & n1127 ) | ( ~n1024 & n1128 ) | ( n1127 & n1128 ) ;
  assign n1130 = ( n1024 & n1127 ) | ( n1024 & n1128 ) | ( n1127 & n1128 ) ;
  assign n1131 = ( n1024 & n1129 ) | ( n1024 & ~n1130 ) | ( n1129 & ~n1130 ) ;
  assign n1132 = ( x72 & n1126 ) | ( x72 & ~n1131 ) | ( n1126 & ~n1131 ) ;
  assign n1133 = ( x72 & n1025 ) | ( x72 & ~n1080 ) | ( n1025 & ~n1080 ) ;
  assign n1134 = x72 & n1025 ;
  assign n1135 = ( ~n1030 & n1133 ) | ( ~n1030 & n1134 ) | ( n1133 & n1134 ) ;
  assign n1136 = ( n1030 & n1133 ) | ( n1030 & n1134 ) | ( n1133 & n1134 ) ;
  assign n1137 = ( n1030 & n1135 ) | ( n1030 & ~n1136 ) | ( n1135 & ~n1136 ) ;
  assign n1138 = ( x73 & n1132 ) | ( x73 & ~n1137 ) | ( n1132 & ~n1137 ) ;
  assign n1139 = ( x73 & n1031 ) | ( x73 & ~n1080 ) | ( n1031 & ~n1080 ) ;
  assign n1140 = x73 & n1031 ;
  assign n1141 = ( ~n1036 & n1139 ) | ( ~n1036 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = ( n1036 & n1139 ) | ( n1036 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1143 = ( n1036 & n1141 ) | ( n1036 & ~n1142 ) | ( n1141 & ~n1142 ) ;
  assign n1144 = ( x74 & n1138 ) | ( x74 & ~n1143 ) | ( n1138 & ~n1143 ) ;
  assign n1145 = ( x74 & n1037 ) | ( x74 & ~n1080 ) | ( n1037 & ~n1080 ) ;
  assign n1146 = x74 & n1037 ;
  assign n1147 = ( ~n1042 & n1145 ) | ( ~n1042 & n1146 ) | ( n1145 & n1146 ) ;
  assign n1148 = ( n1042 & n1145 ) | ( n1042 & n1146 ) | ( n1145 & n1146 ) ;
  assign n1149 = ( n1042 & n1147 ) | ( n1042 & ~n1148 ) | ( n1147 & ~n1148 ) ;
  assign n1150 = ( x75 & n1144 ) | ( x75 & ~n1149 ) | ( n1144 & ~n1149 ) ;
  assign n1151 = ( x75 & n1043 ) | ( x75 & ~n1080 ) | ( n1043 & ~n1080 ) ;
  assign n1152 = x75 & n1043 ;
  assign n1153 = ( ~n1048 & n1151 ) | ( ~n1048 & n1152 ) | ( n1151 & n1152 ) ;
  assign n1154 = ( n1048 & n1151 ) | ( n1048 & n1152 ) | ( n1151 & n1152 ) ;
  assign n1155 = ( n1048 & n1153 ) | ( n1048 & ~n1154 ) | ( n1153 & ~n1154 ) ;
  assign n1156 = ( x76 & n1150 ) | ( x76 & ~n1155 ) | ( n1150 & ~n1155 ) ;
  assign n1157 = ( x76 & n1049 ) | ( x76 & ~n1080 ) | ( n1049 & ~n1080 ) ;
  assign n1158 = x76 & n1049 ;
  assign n1159 = ( ~n1054 & n1157 ) | ( ~n1054 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1160 = ( n1054 & n1157 ) | ( n1054 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1161 = ( n1054 & n1159 ) | ( n1054 & ~n1160 ) | ( n1159 & ~n1160 ) ;
  assign n1162 = ( x77 & n1156 ) | ( x77 & ~n1161 ) | ( n1156 & ~n1161 ) ;
  assign n1163 = ( x77 & n1055 ) | ( x77 & ~n1080 ) | ( n1055 & ~n1080 ) ;
  assign n1164 = x77 & n1055 ;
  assign n1165 = ( ~n1060 & n1163 ) | ( ~n1060 & n1164 ) | ( n1163 & n1164 ) ;
  assign n1166 = ( n1060 & n1163 ) | ( n1060 & n1164 ) | ( n1163 & n1164 ) ;
  assign n1167 = ( n1060 & n1165 ) | ( n1060 & ~n1166 ) | ( n1165 & ~n1166 ) ;
  assign n1168 = ( x78 & n1162 ) | ( x78 & ~n1167 ) | ( n1162 & ~n1167 ) ;
  assign n1169 = ( x78 & n1061 ) | ( x78 & ~n1080 ) | ( n1061 & ~n1080 ) ;
  assign n1170 = x78 & n1061 ;
  assign n1171 = ( ~n1066 & n1169 ) | ( ~n1066 & n1170 ) | ( n1169 & n1170 ) ;
  assign n1172 = ( n1066 & n1169 ) | ( n1066 & n1170 ) | ( n1169 & n1170 ) ;
  assign n1173 = ( n1066 & n1171 ) | ( n1066 & ~n1172 ) | ( n1171 & ~n1172 ) ;
  assign n1174 = ( x79 & n1168 ) | ( x79 & ~n1173 ) | ( n1168 & ~n1173 ) ;
  assign n1175 = ( x79 & n1067 ) | ( x79 & ~n1080 ) | ( n1067 & ~n1080 ) ;
  assign n1176 = x79 & n1067 ;
  assign n1177 = ( ~n1072 & n1175 ) | ( ~n1072 & n1176 ) | ( n1175 & n1176 ) ;
  assign n1178 = ( n1072 & n1175 ) | ( n1072 & n1176 ) | ( n1175 & n1176 ) ;
  assign n1179 = ( n1072 & n1177 ) | ( n1072 & ~n1178 ) | ( n1177 & ~n1178 ) ;
  assign n1180 = ( x80 & n1174 ) | ( x80 & ~n1179 ) | ( n1174 & ~n1179 ) ;
  assign n1181 = ~n176 & n1075 ;
  assign n1182 = n175 & n976 ;
  assign n1183 = ( n976 & n1075 ) | ( n976 & n1182 ) | ( n1075 & n1182 ) ;
  assign n1184 = n1078 | n1183 ;
  assign n1185 = ~n1181 & n1184 ;
  assign n1186 = ( x81 & ~n1085 ) | ( x81 & n1180 ) | ( ~n1085 & n1180 ) ;
  assign n1187 = ( x82 & ~n1185 ) | ( x82 & n1186 ) | ( ~n1185 & n1186 ) ;
  assign n1188 = n174 | n1187 ;
  assign n1189 = ( x81 & n1180 ) | ( x81 & n1188 ) | ( n1180 & n1188 ) ;
  assign n1190 = x81 | n1180 ;
  assign n1191 = ( ~n1085 & n1189 ) | ( ~n1085 & n1190 ) | ( n1189 & n1190 ) ;
  assign n1192 = ( n1085 & n1189 ) | ( n1085 & n1190 ) | ( n1189 & n1190 ) ;
  assign n1193 = ( n1085 & n1191 ) | ( n1085 & ~n1192 ) | ( n1191 & ~n1192 ) ;
  assign n1194 = ~x44 & x64 ;
  assign n1195 = ~x45 & n1188 ;
  assign n1196 = ( x45 & ~x64 ) | ( x45 & n1188 ) | ( ~x64 & n1188 ) ;
  assign n1197 = ( n1086 & ~n1195 ) | ( n1086 & n1196 ) | ( ~n1195 & n1196 ) ;
  assign n1198 = ( x65 & n1194 ) | ( x65 & ~n1197 ) | ( n1194 & ~n1197 ) ;
  assign n1199 = ( x65 & n1086 ) | ( x65 & n1188 ) | ( n1086 & n1188 ) ;
  assign n1200 = x65 | n1086 ;
  assign n1201 = ( ~n1089 & n1199 ) | ( ~n1089 & n1200 ) | ( n1199 & n1200 ) ;
  assign n1202 = ( n1089 & n1199 ) | ( n1089 & n1200 ) | ( n1199 & n1200 ) ;
  assign n1203 = ( n1089 & n1201 ) | ( n1089 & ~n1202 ) | ( n1201 & ~n1202 ) ;
  assign n1204 = ( x66 & n1198 ) | ( x66 & ~n1203 ) | ( n1198 & ~n1203 ) ;
  assign n1205 = ( x66 & n1090 ) | ( x66 & n1188 ) | ( n1090 & n1188 ) ;
  assign n1206 = x66 | n1090 ;
  assign n1207 = ( ~n1095 & n1205 ) | ( ~n1095 & n1206 ) | ( n1205 & n1206 ) ;
  assign n1208 = ( n1095 & n1205 ) | ( n1095 & n1206 ) | ( n1205 & n1206 ) ;
  assign n1209 = ( n1095 & n1207 ) | ( n1095 & ~n1208 ) | ( n1207 & ~n1208 ) ;
  assign n1210 = ( x67 & n1204 ) | ( x67 & ~n1209 ) | ( n1204 & ~n1209 ) ;
  assign n1211 = ( x67 & n1096 ) | ( x67 & n1188 ) | ( n1096 & n1188 ) ;
  assign n1212 = x67 | n1096 ;
  assign n1213 = ( ~n1101 & n1211 ) | ( ~n1101 & n1212 ) | ( n1211 & n1212 ) ;
  assign n1214 = ( n1101 & n1211 ) | ( n1101 & n1212 ) | ( n1211 & n1212 ) ;
  assign n1215 = ( n1101 & n1213 ) | ( n1101 & ~n1214 ) | ( n1213 & ~n1214 ) ;
  assign n1216 = ( x68 & n1210 ) | ( x68 & ~n1215 ) | ( n1210 & ~n1215 ) ;
  assign n1217 = ( x68 & n1102 ) | ( x68 & ~n1188 ) | ( n1102 & ~n1188 ) ;
  assign n1218 = x68 & n1102 ;
  assign n1219 = ( ~n1107 & n1217 ) | ( ~n1107 & n1218 ) | ( n1217 & n1218 ) ;
  assign n1220 = ( n1107 & n1217 ) | ( n1107 & n1218 ) | ( n1217 & n1218 ) ;
  assign n1221 = ( n1107 & n1219 ) | ( n1107 & ~n1220 ) | ( n1219 & ~n1220 ) ;
  assign n1222 = ( x69 & n1216 ) | ( x69 & ~n1221 ) | ( n1216 & ~n1221 ) ;
  assign n1223 = ( x69 & n1108 ) | ( x69 & ~n1188 ) | ( n1108 & ~n1188 ) ;
  assign n1224 = x69 & n1108 ;
  assign n1225 = ( ~n1113 & n1223 ) | ( ~n1113 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = ( n1113 & n1223 ) | ( n1113 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1227 = ( n1113 & n1225 ) | ( n1113 & ~n1226 ) | ( n1225 & ~n1226 ) ;
  assign n1228 = ( x70 & n1222 ) | ( x70 & ~n1227 ) | ( n1222 & ~n1227 ) ;
  assign n1229 = ( x70 & n1114 ) | ( x70 & ~n1188 ) | ( n1114 & ~n1188 ) ;
  assign n1230 = x70 & n1114 ;
  assign n1231 = ( ~n1119 & n1229 ) | ( ~n1119 & n1230 ) | ( n1229 & n1230 ) ;
  assign n1232 = ( n1119 & n1229 ) | ( n1119 & n1230 ) | ( n1229 & n1230 ) ;
  assign n1233 = ( n1119 & n1231 ) | ( n1119 & ~n1232 ) | ( n1231 & ~n1232 ) ;
  assign n1234 = ( x71 & n1228 ) | ( x71 & ~n1233 ) | ( n1228 & ~n1233 ) ;
  assign n1235 = ( x71 & n1120 ) | ( x71 & ~n1188 ) | ( n1120 & ~n1188 ) ;
  assign n1236 = x71 & n1120 ;
  assign n1237 = ( ~n1125 & n1235 ) | ( ~n1125 & n1236 ) | ( n1235 & n1236 ) ;
  assign n1238 = ( n1125 & n1235 ) | ( n1125 & n1236 ) | ( n1235 & n1236 ) ;
  assign n1239 = ( n1125 & n1237 ) | ( n1125 & ~n1238 ) | ( n1237 & ~n1238 ) ;
  assign n1240 = ( x72 & n1234 ) | ( x72 & ~n1239 ) | ( n1234 & ~n1239 ) ;
  assign n1241 = ( x72 & n1126 ) | ( x72 & ~n1188 ) | ( n1126 & ~n1188 ) ;
  assign n1242 = x72 & n1126 ;
  assign n1243 = ( ~n1131 & n1241 ) | ( ~n1131 & n1242 ) | ( n1241 & n1242 ) ;
  assign n1244 = ( n1131 & n1241 ) | ( n1131 & n1242 ) | ( n1241 & n1242 ) ;
  assign n1245 = ( n1131 & n1243 ) | ( n1131 & ~n1244 ) | ( n1243 & ~n1244 ) ;
  assign n1246 = ( x73 & n1240 ) | ( x73 & ~n1245 ) | ( n1240 & ~n1245 ) ;
  assign n1247 = ( x73 & n1132 ) | ( x73 & ~n1188 ) | ( n1132 & ~n1188 ) ;
  assign n1248 = x73 & n1132 ;
  assign n1249 = ( ~n1137 & n1247 ) | ( ~n1137 & n1248 ) | ( n1247 & n1248 ) ;
  assign n1250 = ( n1137 & n1247 ) | ( n1137 & n1248 ) | ( n1247 & n1248 ) ;
  assign n1251 = ( n1137 & n1249 ) | ( n1137 & ~n1250 ) | ( n1249 & ~n1250 ) ;
  assign n1252 = ( x74 & n1246 ) | ( x74 & ~n1251 ) | ( n1246 & ~n1251 ) ;
  assign n1253 = ( x74 & n1138 ) | ( x74 & ~n1188 ) | ( n1138 & ~n1188 ) ;
  assign n1254 = x74 & n1138 ;
  assign n1255 = ( ~n1143 & n1253 ) | ( ~n1143 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1256 = ( n1143 & n1253 ) | ( n1143 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1257 = ( n1143 & n1255 ) | ( n1143 & ~n1256 ) | ( n1255 & ~n1256 ) ;
  assign n1258 = ( x75 & n1252 ) | ( x75 & ~n1257 ) | ( n1252 & ~n1257 ) ;
  assign n1259 = ( x75 & n1144 ) | ( x75 & ~n1188 ) | ( n1144 & ~n1188 ) ;
  assign n1260 = x75 & n1144 ;
  assign n1261 = ( ~n1149 & n1259 ) | ( ~n1149 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1262 = ( n1149 & n1259 ) | ( n1149 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1263 = ( n1149 & n1261 ) | ( n1149 & ~n1262 ) | ( n1261 & ~n1262 ) ;
  assign n1264 = ( x76 & n1258 ) | ( x76 & ~n1263 ) | ( n1258 & ~n1263 ) ;
  assign n1265 = ( x76 & n1150 ) | ( x76 & ~n1188 ) | ( n1150 & ~n1188 ) ;
  assign n1266 = x76 & n1150 ;
  assign n1267 = ( ~n1155 & n1265 ) | ( ~n1155 & n1266 ) | ( n1265 & n1266 ) ;
  assign n1268 = ( n1155 & n1265 ) | ( n1155 & n1266 ) | ( n1265 & n1266 ) ;
  assign n1269 = ( n1155 & n1267 ) | ( n1155 & ~n1268 ) | ( n1267 & ~n1268 ) ;
  assign n1270 = ( x77 & n1264 ) | ( x77 & ~n1269 ) | ( n1264 & ~n1269 ) ;
  assign n1271 = ( x77 & n1156 ) | ( x77 & ~n1188 ) | ( n1156 & ~n1188 ) ;
  assign n1272 = x77 & n1156 ;
  assign n1273 = ( ~n1161 & n1271 ) | ( ~n1161 & n1272 ) | ( n1271 & n1272 ) ;
  assign n1274 = ( n1161 & n1271 ) | ( n1161 & n1272 ) | ( n1271 & n1272 ) ;
  assign n1275 = ( n1161 & n1273 ) | ( n1161 & ~n1274 ) | ( n1273 & ~n1274 ) ;
  assign n1276 = ( x78 & n1270 ) | ( x78 & ~n1275 ) | ( n1270 & ~n1275 ) ;
  assign n1277 = ( x78 & n1162 ) | ( x78 & ~n1188 ) | ( n1162 & ~n1188 ) ;
  assign n1278 = x78 & n1162 ;
  assign n1279 = ( ~n1167 & n1277 ) | ( ~n1167 & n1278 ) | ( n1277 & n1278 ) ;
  assign n1280 = ( n1167 & n1277 ) | ( n1167 & n1278 ) | ( n1277 & n1278 ) ;
  assign n1281 = ( n1167 & n1279 ) | ( n1167 & ~n1280 ) | ( n1279 & ~n1280 ) ;
  assign n1282 = ( x79 & n1276 ) | ( x79 & ~n1281 ) | ( n1276 & ~n1281 ) ;
  assign n1283 = ( x79 & n1168 ) | ( x79 & ~n1188 ) | ( n1168 & ~n1188 ) ;
  assign n1284 = x79 & n1168 ;
  assign n1285 = ( ~n1173 & n1283 ) | ( ~n1173 & n1284 ) | ( n1283 & n1284 ) ;
  assign n1286 = ( n1173 & n1283 ) | ( n1173 & n1284 ) | ( n1283 & n1284 ) ;
  assign n1287 = ( n1173 & n1285 ) | ( n1173 & ~n1286 ) | ( n1285 & ~n1286 ) ;
  assign n1288 = ( x80 & n1282 ) | ( x80 & ~n1287 ) | ( n1282 & ~n1287 ) ;
  assign n1289 = ( x80 & n1174 ) | ( x80 & ~n1188 ) | ( n1174 & ~n1188 ) ;
  assign n1290 = x80 & n1174 ;
  assign n1291 = ( ~n1179 & n1289 ) | ( ~n1179 & n1290 ) | ( n1289 & n1290 ) ;
  assign n1292 = ( n1179 & n1289 ) | ( n1179 & n1290 ) | ( n1289 & n1290 ) ;
  assign n1293 = ( n1179 & n1291 ) | ( n1179 & ~n1292 ) | ( n1291 & ~n1292 ) ;
  assign n1294 = ( x81 & n1288 ) | ( x81 & ~n1293 ) | ( n1288 & ~n1293 ) ;
  assign n1295 = ( x82 & n174 ) | ( x82 & n1186 ) | ( n174 & n1186 ) ;
  assign n1296 = x82 | n1186 ;
  assign n1297 = ( n1185 & n1295 ) | ( n1185 & ~n1296 ) | ( n1295 & ~n1296 ) ;
  assign n1298 = ( x82 & ~n1193 ) | ( x82 & n1294 ) | ( ~n1193 & n1294 ) ;
  assign n1299 = ( x83 & ~n1297 ) | ( x83 & n1298 ) | ( ~n1297 & n1298 ) ;
  assign n1300 = n173 | n1299 ;
  assign n1301 = ( x82 & n1294 ) | ( x82 & n1300 ) | ( n1294 & n1300 ) ;
  assign n1302 = x82 | n1294 ;
  assign n1303 = ( ~n1193 & n1301 ) | ( ~n1193 & n1302 ) | ( n1301 & n1302 ) ;
  assign n1304 = ( n1193 & n1301 ) | ( n1193 & n1302 ) | ( n1301 & n1302 ) ;
  assign n1305 = ( n1193 & n1303 ) | ( n1193 & ~n1304 ) | ( n1303 & ~n1304 ) ;
  assign n1306 = ~x43 & x64 ;
  assign n1307 = ~x44 & n1300 ;
  assign n1308 = ( x44 & ~x64 ) | ( x44 & n1300 ) | ( ~x64 & n1300 ) ;
  assign n1309 = ( n1194 & ~n1307 ) | ( n1194 & n1308 ) | ( ~n1307 & n1308 ) ;
  assign n1310 = ( x65 & n1306 ) | ( x65 & ~n1309 ) | ( n1306 & ~n1309 ) ;
  assign n1311 = ( x65 & n1194 ) | ( x65 & n1300 ) | ( n1194 & n1300 ) ;
  assign n1312 = x65 | n1194 ;
  assign n1313 = ( ~n1197 & n1311 ) | ( ~n1197 & n1312 ) | ( n1311 & n1312 ) ;
  assign n1314 = ( n1197 & n1311 ) | ( n1197 & n1312 ) | ( n1311 & n1312 ) ;
  assign n1315 = ( n1197 & n1313 ) | ( n1197 & ~n1314 ) | ( n1313 & ~n1314 ) ;
  assign n1316 = ( x66 & n1310 ) | ( x66 & ~n1315 ) | ( n1310 & ~n1315 ) ;
  assign n1317 = ( x66 & n1198 ) | ( x66 & n1300 ) | ( n1198 & n1300 ) ;
  assign n1318 = x66 | n1198 ;
  assign n1319 = ( ~n1203 & n1317 ) | ( ~n1203 & n1318 ) | ( n1317 & n1318 ) ;
  assign n1320 = ( n1203 & n1317 ) | ( n1203 & n1318 ) | ( n1317 & n1318 ) ;
  assign n1321 = ( n1203 & n1319 ) | ( n1203 & ~n1320 ) | ( n1319 & ~n1320 ) ;
  assign n1322 = ( x67 & n1316 ) | ( x67 & ~n1321 ) | ( n1316 & ~n1321 ) ;
  assign n1323 = ( x67 & n1204 ) | ( x67 & ~n1300 ) | ( n1204 & ~n1300 ) ;
  assign n1324 = x67 & n1204 ;
  assign n1325 = ( ~n1209 & n1323 ) | ( ~n1209 & n1324 ) | ( n1323 & n1324 ) ;
  assign n1326 = ( n1209 & n1323 ) | ( n1209 & n1324 ) | ( n1323 & n1324 ) ;
  assign n1327 = ( n1209 & n1325 ) | ( n1209 & ~n1326 ) | ( n1325 & ~n1326 ) ;
  assign n1328 = ( x68 & n1322 ) | ( x68 & ~n1327 ) | ( n1322 & ~n1327 ) ;
  assign n1329 = ( x68 & n1210 ) | ( x68 & ~n1300 ) | ( n1210 & ~n1300 ) ;
  assign n1330 = x68 & n1210 ;
  assign n1331 = ( ~n1215 & n1329 ) | ( ~n1215 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1332 = ( n1215 & n1329 ) | ( n1215 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1333 = ( n1215 & n1331 ) | ( n1215 & ~n1332 ) | ( n1331 & ~n1332 ) ;
  assign n1334 = ( x69 & n1328 ) | ( x69 & ~n1333 ) | ( n1328 & ~n1333 ) ;
  assign n1335 = ( x69 & n1216 ) | ( x69 & ~n1300 ) | ( n1216 & ~n1300 ) ;
  assign n1336 = x69 & n1216 ;
  assign n1337 = ( ~n1221 & n1335 ) | ( ~n1221 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1338 = ( n1221 & n1335 ) | ( n1221 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1339 = ( n1221 & n1337 ) | ( n1221 & ~n1338 ) | ( n1337 & ~n1338 ) ;
  assign n1340 = ( x70 & n1334 ) | ( x70 & ~n1339 ) | ( n1334 & ~n1339 ) ;
  assign n1341 = ( x70 & n1222 ) | ( x70 & ~n1300 ) | ( n1222 & ~n1300 ) ;
  assign n1342 = x70 & n1222 ;
  assign n1343 = ( ~n1227 & n1341 ) | ( ~n1227 & n1342 ) | ( n1341 & n1342 ) ;
  assign n1344 = ( n1227 & n1341 ) | ( n1227 & n1342 ) | ( n1341 & n1342 ) ;
  assign n1345 = ( n1227 & n1343 ) | ( n1227 & ~n1344 ) | ( n1343 & ~n1344 ) ;
  assign n1346 = ( x71 & n1340 ) | ( x71 & ~n1345 ) | ( n1340 & ~n1345 ) ;
  assign n1347 = ( x71 & n1228 ) | ( x71 & ~n1300 ) | ( n1228 & ~n1300 ) ;
  assign n1348 = x71 & n1228 ;
  assign n1349 = ( ~n1233 & n1347 ) | ( ~n1233 & n1348 ) | ( n1347 & n1348 ) ;
  assign n1350 = ( n1233 & n1347 ) | ( n1233 & n1348 ) | ( n1347 & n1348 ) ;
  assign n1351 = ( n1233 & n1349 ) | ( n1233 & ~n1350 ) | ( n1349 & ~n1350 ) ;
  assign n1352 = ( x72 & n1346 ) | ( x72 & ~n1351 ) | ( n1346 & ~n1351 ) ;
  assign n1353 = ( x72 & n1234 ) | ( x72 & ~n1300 ) | ( n1234 & ~n1300 ) ;
  assign n1354 = x72 & n1234 ;
  assign n1355 = ( ~n1239 & n1353 ) | ( ~n1239 & n1354 ) | ( n1353 & n1354 ) ;
  assign n1356 = ( n1239 & n1353 ) | ( n1239 & n1354 ) | ( n1353 & n1354 ) ;
  assign n1357 = ( n1239 & n1355 ) | ( n1239 & ~n1356 ) | ( n1355 & ~n1356 ) ;
  assign n1358 = ( x73 & n1352 ) | ( x73 & ~n1357 ) | ( n1352 & ~n1357 ) ;
  assign n1359 = ( x73 & n1240 ) | ( x73 & ~n1300 ) | ( n1240 & ~n1300 ) ;
  assign n1360 = x73 & n1240 ;
  assign n1361 = ( ~n1245 & n1359 ) | ( ~n1245 & n1360 ) | ( n1359 & n1360 ) ;
  assign n1362 = ( n1245 & n1359 ) | ( n1245 & n1360 ) | ( n1359 & n1360 ) ;
  assign n1363 = ( n1245 & n1361 ) | ( n1245 & ~n1362 ) | ( n1361 & ~n1362 ) ;
  assign n1364 = ( x74 & n1358 ) | ( x74 & ~n1363 ) | ( n1358 & ~n1363 ) ;
  assign n1365 = ( x74 & n1246 ) | ( x74 & ~n1300 ) | ( n1246 & ~n1300 ) ;
  assign n1366 = x74 & n1246 ;
  assign n1367 = ( ~n1251 & n1365 ) | ( ~n1251 & n1366 ) | ( n1365 & n1366 ) ;
  assign n1368 = ( n1251 & n1365 ) | ( n1251 & n1366 ) | ( n1365 & n1366 ) ;
  assign n1369 = ( n1251 & n1367 ) | ( n1251 & ~n1368 ) | ( n1367 & ~n1368 ) ;
  assign n1370 = ( x75 & n1364 ) | ( x75 & ~n1369 ) | ( n1364 & ~n1369 ) ;
  assign n1371 = ( x75 & n1252 ) | ( x75 & ~n1300 ) | ( n1252 & ~n1300 ) ;
  assign n1372 = x75 & n1252 ;
  assign n1373 = ( ~n1257 & n1371 ) | ( ~n1257 & n1372 ) | ( n1371 & n1372 ) ;
  assign n1374 = ( n1257 & n1371 ) | ( n1257 & n1372 ) | ( n1371 & n1372 ) ;
  assign n1375 = ( n1257 & n1373 ) | ( n1257 & ~n1374 ) | ( n1373 & ~n1374 ) ;
  assign n1376 = ( x76 & n1370 ) | ( x76 & ~n1375 ) | ( n1370 & ~n1375 ) ;
  assign n1377 = ( x76 & n1258 ) | ( x76 & ~n1300 ) | ( n1258 & ~n1300 ) ;
  assign n1378 = x76 & n1258 ;
  assign n1379 = ( ~n1263 & n1377 ) | ( ~n1263 & n1378 ) | ( n1377 & n1378 ) ;
  assign n1380 = ( n1263 & n1377 ) | ( n1263 & n1378 ) | ( n1377 & n1378 ) ;
  assign n1381 = ( n1263 & n1379 ) | ( n1263 & ~n1380 ) | ( n1379 & ~n1380 ) ;
  assign n1382 = ( x77 & n1376 ) | ( x77 & ~n1381 ) | ( n1376 & ~n1381 ) ;
  assign n1383 = ( x77 & n1264 ) | ( x77 & ~n1300 ) | ( n1264 & ~n1300 ) ;
  assign n1384 = x77 & n1264 ;
  assign n1385 = ( ~n1269 & n1383 ) | ( ~n1269 & n1384 ) | ( n1383 & n1384 ) ;
  assign n1386 = ( n1269 & n1383 ) | ( n1269 & n1384 ) | ( n1383 & n1384 ) ;
  assign n1387 = ( n1269 & n1385 ) | ( n1269 & ~n1386 ) | ( n1385 & ~n1386 ) ;
  assign n1388 = ( x78 & n1382 ) | ( x78 & ~n1387 ) | ( n1382 & ~n1387 ) ;
  assign n1389 = ( x78 & n1270 ) | ( x78 & ~n1300 ) | ( n1270 & ~n1300 ) ;
  assign n1390 = x78 & n1270 ;
  assign n1391 = ( ~n1275 & n1389 ) | ( ~n1275 & n1390 ) | ( n1389 & n1390 ) ;
  assign n1392 = ( n1275 & n1389 ) | ( n1275 & n1390 ) | ( n1389 & n1390 ) ;
  assign n1393 = ( n1275 & n1391 ) | ( n1275 & ~n1392 ) | ( n1391 & ~n1392 ) ;
  assign n1394 = ( x79 & n1388 ) | ( x79 & ~n1393 ) | ( n1388 & ~n1393 ) ;
  assign n1395 = ( x79 & n1276 ) | ( x79 & ~n1300 ) | ( n1276 & ~n1300 ) ;
  assign n1396 = x79 & n1276 ;
  assign n1397 = ( ~n1281 & n1395 ) | ( ~n1281 & n1396 ) | ( n1395 & n1396 ) ;
  assign n1398 = ( n1281 & n1395 ) | ( n1281 & n1396 ) | ( n1395 & n1396 ) ;
  assign n1399 = ( n1281 & n1397 ) | ( n1281 & ~n1398 ) | ( n1397 & ~n1398 ) ;
  assign n1400 = ( x80 & n1394 ) | ( x80 & ~n1399 ) | ( n1394 & ~n1399 ) ;
  assign n1401 = ( x80 & n1282 ) | ( x80 & ~n1300 ) | ( n1282 & ~n1300 ) ;
  assign n1402 = x80 & n1282 ;
  assign n1403 = ( ~n1287 & n1401 ) | ( ~n1287 & n1402 ) | ( n1401 & n1402 ) ;
  assign n1404 = ( n1287 & n1401 ) | ( n1287 & n1402 ) | ( n1401 & n1402 ) ;
  assign n1405 = ( n1287 & n1403 ) | ( n1287 & ~n1404 ) | ( n1403 & ~n1404 ) ;
  assign n1406 = ( x81 & n1400 ) | ( x81 & ~n1405 ) | ( n1400 & ~n1405 ) ;
  assign n1407 = ( x81 & n1288 ) | ( x81 & ~n1300 ) | ( n1288 & ~n1300 ) ;
  assign n1408 = x81 & n1288 ;
  assign n1409 = ( ~n1293 & n1407 ) | ( ~n1293 & n1408 ) | ( n1407 & n1408 ) ;
  assign n1410 = ( n1293 & n1407 ) | ( n1293 & n1408 ) | ( n1407 & n1408 ) ;
  assign n1411 = ( n1293 & n1409 ) | ( n1293 & ~n1410 ) | ( n1409 & ~n1410 ) ;
  assign n1412 = ( x82 & n1406 ) | ( x82 & ~n1411 ) | ( n1406 & ~n1411 ) ;
  assign n1413 = ( x83 & ~n1305 ) | ( x83 & n1412 ) | ( ~n1305 & n1412 ) ;
  assign n1414 = n172 | n1413 ;
  assign n1415 = ( ~x83 & n173 ) | ( ~x83 & n1298 ) | ( n173 & n1298 ) ;
  assign n1416 = ( ~x83 & n1297 ) | ( ~x83 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1417 = ~n1415 & n1416 ;
  assign n1418 = x84 & ~n1297 ;
  assign n1419 = ( n1414 & ~n1417 ) | ( n1414 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = ( x83 & n1412 ) | ( x83 & ~n1419 ) | ( n1412 & ~n1419 ) ;
  assign n1421 = x83 & n1412 ;
  assign n1422 = ( ~n1305 & n1420 ) | ( ~n1305 & n1421 ) | ( n1420 & n1421 ) ;
  assign n1423 = ( n1305 & n1420 ) | ( n1305 & n1421 ) | ( n1420 & n1421 ) ;
  assign n1424 = ( n1305 & n1422 ) | ( n1305 & ~n1423 ) | ( n1422 & ~n1423 ) ;
  assign n1425 = ~x42 & x64 ;
  assign n1426 = x43 & n1419 ;
  assign n1427 = ( x43 & x64 ) | ( x43 & ~n1419 ) | ( x64 & ~n1419 ) ;
  assign n1428 = x43 & x64 ;
  assign n1429 = ( n1426 & n1427 ) | ( n1426 & ~n1428 ) | ( n1427 & ~n1428 ) ;
  assign n1430 = ( x65 & n1425 ) | ( x65 & ~n1429 ) | ( n1425 & ~n1429 ) ;
  assign n1431 = ( x65 & n1306 ) | ( x65 & n1419 ) | ( n1306 & n1419 ) ;
  assign n1432 = x65 | n1306 ;
  assign n1433 = ( ~n1309 & n1431 ) | ( ~n1309 & n1432 ) | ( n1431 & n1432 ) ;
  assign n1434 = ( n1309 & n1431 ) | ( n1309 & n1432 ) | ( n1431 & n1432 ) ;
  assign n1435 = ( n1309 & n1433 ) | ( n1309 & ~n1434 ) | ( n1433 & ~n1434 ) ;
  assign n1436 = ( x66 & n1430 ) | ( x66 & ~n1435 ) | ( n1430 & ~n1435 ) ;
  assign n1437 = ( x66 & n1310 ) | ( x66 & n1419 ) | ( n1310 & n1419 ) ;
  assign n1438 = x66 | n1310 ;
  assign n1439 = ( ~n1315 & n1437 ) | ( ~n1315 & n1438 ) | ( n1437 & n1438 ) ;
  assign n1440 = ( n1315 & n1437 ) | ( n1315 & n1438 ) | ( n1437 & n1438 ) ;
  assign n1441 = ( n1315 & n1439 ) | ( n1315 & ~n1440 ) | ( n1439 & ~n1440 ) ;
  assign n1442 = ( x67 & n1436 ) | ( x67 & ~n1441 ) | ( n1436 & ~n1441 ) ;
  assign n1443 = ( x67 & n1316 ) | ( x67 & ~n1419 ) | ( n1316 & ~n1419 ) ;
  assign n1444 = x67 & n1316 ;
  assign n1445 = ( ~n1321 & n1443 ) | ( ~n1321 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1446 = ( n1321 & n1443 ) | ( n1321 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1447 = ( n1321 & n1445 ) | ( n1321 & ~n1446 ) | ( n1445 & ~n1446 ) ;
  assign n1448 = ( x68 & n1442 ) | ( x68 & ~n1447 ) | ( n1442 & ~n1447 ) ;
  assign n1449 = ( x68 & n1322 ) | ( x68 & ~n1419 ) | ( n1322 & ~n1419 ) ;
  assign n1450 = x68 & n1322 ;
  assign n1451 = ( ~n1327 & n1449 ) | ( ~n1327 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1452 = ( n1327 & n1449 ) | ( n1327 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1453 = ( n1327 & n1451 ) | ( n1327 & ~n1452 ) | ( n1451 & ~n1452 ) ;
  assign n1454 = ( x69 & n1448 ) | ( x69 & ~n1453 ) | ( n1448 & ~n1453 ) ;
  assign n1455 = ( x69 & n1328 ) | ( x69 & ~n1419 ) | ( n1328 & ~n1419 ) ;
  assign n1456 = x69 & n1328 ;
  assign n1457 = ( ~n1333 & n1455 ) | ( ~n1333 & n1456 ) | ( n1455 & n1456 ) ;
  assign n1458 = ( n1333 & n1455 ) | ( n1333 & n1456 ) | ( n1455 & n1456 ) ;
  assign n1459 = ( n1333 & n1457 ) | ( n1333 & ~n1458 ) | ( n1457 & ~n1458 ) ;
  assign n1460 = ( x70 & n1454 ) | ( x70 & ~n1459 ) | ( n1454 & ~n1459 ) ;
  assign n1461 = ( x70 & n1334 ) | ( x70 & ~n1419 ) | ( n1334 & ~n1419 ) ;
  assign n1462 = x70 & n1334 ;
  assign n1463 = ( ~n1339 & n1461 ) | ( ~n1339 & n1462 ) | ( n1461 & n1462 ) ;
  assign n1464 = ( n1339 & n1461 ) | ( n1339 & n1462 ) | ( n1461 & n1462 ) ;
  assign n1465 = ( n1339 & n1463 ) | ( n1339 & ~n1464 ) | ( n1463 & ~n1464 ) ;
  assign n1466 = ( x71 & n1460 ) | ( x71 & ~n1465 ) | ( n1460 & ~n1465 ) ;
  assign n1467 = ( x71 & n1340 ) | ( x71 & ~n1419 ) | ( n1340 & ~n1419 ) ;
  assign n1468 = x71 & n1340 ;
  assign n1469 = ( ~n1345 & n1467 ) | ( ~n1345 & n1468 ) | ( n1467 & n1468 ) ;
  assign n1470 = ( n1345 & n1467 ) | ( n1345 & n1468 ) | ( n1467 & n1468 ) ;
  assign n1471 = ( n1345 & n1469 ) | ( n1345 & ~n1470 ) | ( n1469 & ~n1470 ) ;
  assign n1472 = ( x72 & n1466 ) | ( x72 & ~n1471 ) | ( n1466 & ~n1471 ) ;
  assign n1473 = ( x72 & n1346 ) | ( x72 & ~n1419 ) | ( n1346 & ~n1419 ) ;
  assign n1474 = x72 & n1346 ;
  assign n1475 = ( ~n1351 & n1473 ) | ( ~n1351 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ( n1351 & n1473 ) | ( n1351 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1477 = ( n1351 & n1475 ) | ( n1351 & ~n1476 ) | ( n1475 & ~n1476 ) ;
  assign n1478 = ( x73 & n1472 ) | ( x73 & ~n1477 ) | ( n1472 & ~n1477 ) ;
  assign n1479 = ( x73 & n1352 ) | ( x73 & ~n1419 ) | ( n1352 & ~n1419 ) ;
  assign n1480 = x73 & n1352 ;
  assign n1481 = ( ~n1357 & n1479 ) | ( ~n1357 & n1480 ) | ( n1479 & n1480 ) ;
  assign n1482 = ( n1357 & n1479 ) | ( n1357 & n1480 ) | ( n1479 & n1480 ) ;
  assign n1483 = ( n1357 & n1481 ) | ( n1357 & ~n1482 ) | ( n1481 & ~n1482 ) ;
  assign n1484 = ( x74 & n1478 ) | ( x74 & ~n1483 ) | ( n1478 & ~n1483 ) ;
  assign n1485 = ( x74 & n1358 ) | ( x74 & ~n1419 ) | ( n1358 & ~n1419 ) ;
  assign n1486 = x74 & n1358 ;
  assign n1487 = ( ~n1363 & n1485 ) | ( ~n1363 & n1486 ) | ( n1485 & n1486 ) ;
  assign n1488 = ( n1363 & n1485 ) | ( n1363 & n1486 ) | ( n1485 & n1486 ) ;
  assign n1489 = ( n1363 & n1487 ) | ( n1363 & ~n1488 ) | ( n1487 & ~n1488 ) ;
  assign n1490 = ( x75 & n1484 ) | ( x75 & ~n1489 ) | ( n1484 & ~n1489 ) ;
  assign n1491 = ( x75 & n1364 ) | ( x75 & ~n1419 ) | ( n1364 & ~n1419 ) ;
  assign n1492 = x75 & n1364 ;
  assign n1493 = ( ~n1369 & n1491 ) | ( ~n1369 & n1492 ) | ( n1491 & n1492 ) ;
  assign n1494 = ( n1369 & n1491 ) | ( n1369 & n1492 ) | ( n1491 & n1492 ) ;
  assign n1495 = ( n1369 & n1493 ) | ( n1369 & ~n1494 ) | ( n1493 & ~n1494 ) ;
  assign n1496 = ( x76 & n1490 ) | ( x76 & ~n1495 ) | ( n1490 & ~n1495 ) ;
  assign n1497 = ( x76 & n1370 ) | ( x76 & ~n1419 ) | ( n1370 & ~n1419 ) ;
  assign n1498 = x76 & n1370 ;
  assign n1499 = ( ~n1375 & n1497 ) | ( ~n1375 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1500 = ( n1375 & n1497 ) | ( n1375 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1501 = ( n1375 & n1499 ) | ( n1375 & ~n1500 ) | ( n1499 & ~n1500 ) ;
  assign n1502 = ( x77 & n1496 ) | ( x77 & ~n1501 ) | ( n1496 & ~n1501 ) ;
  assign n1503 = ( x77 & n1376 ) | ( x77 & ~n1419 ) | ( n1376 & ~n1419 ) ;
  assign n1504 = x77 & n1376 ;
  assign n1505 = ( ~n1381 & n1503 ) | ( ~n1381 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1506 = ( n1381 & n1503 ) | ( n1381 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1507 = ( n1381 & n1505 ) | ( n1381 & ~n1506 ) | ( n1505 & ~n1506 ) ;
  assign n1508 = ( x78 & n1502 ) | ( x78 & ~n1507 ) | ( n1502 & ~n1507 ) ;
  assign n1509 = ( x78 & n1382 ) | ( x78 & ~n1419 ) | ( n1382 & ~n1419 ) ;
  assign n1510 = x78 & n1382 ;
  assign n1511 = ( ~n1387 & n1509 ) | ( ~n1387 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = ( n1387 & n1509 ) | ( n1387 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1513 = ( n1387 & n1511 ) | ( n1387 & ~n1512 ) | ( n1511 & ~n1512 ) ;
  assign n1514 = ( x79 & n1508 ) | ( x79 & ~n1513 ) | ( n1508 & ~n1513 ) ;
  assign n1515 = ( x79 & n1388 ) | ( x79 & ~n1419 ) | ( n1388 & ~n1419 ) ;
  assign n1516 = x79 & n1388 ;
  assign n1517 = ( ~n1393 & n1515 ) | ( ~n1393 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = ( n1393 & n1515 ) | ( n1393 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1519 = ( n1393 & n1517 ) | ( n1393 & ~n1518 ) | ( n1517 & ~n1518 ) ;
  assign n1520 = ( x80 & n1514 ) | ( x80 & ~n1519 ) | ( n1514 & ~n1519 ) ;
  assign n1521 = ( x80 & n1394 ) | ( x80 & ~n1419 ) | ( n1394 & ~n1419 ) ;
  assign n1522 = x80 & n1394 ;
  assign n1523 = ( ~n1399 & n1521 ) | ( ~n1399 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1524 = ( n1399 & n1521 ) | ( n1399 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1525 = ( n1399 & n1523 ) | ( n1399 & ~n1524 ) | ( n1523 & ~n1524 ) ;
  assign n1526 = ( x81 & n1520 ) | ( x81 & ~n1525 ) | ( n1520 & ~n1525 ) ;
  assign n1527 = ( x81 & n1400 ) | ( x81 & ~n1419 ) | ( n1400 & ~n1419 ) ;
  assign n1528 = x81 & n1400 ;
  assign n1529 = ( ~n1405 & n1527 ) | ( ~n1405 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1530 = ( n1405 & n1527 ) | ( n1405 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1531 = ( n1405 & n1529 ) | ( n1405 & ~n1530 ) | ( n1529 & ~n1530 ) ;
  assign n1532 = ( x82 & n1526 ) | ( x82 & ~n1531 ) | ( n1526 & ~n1531 ) ;
  assign n1533 = ( x82 & n1406 ) | ( x82 & ~n1419 ) | ( n1406 & ~n1419 ) ;
  assign n1534 = x82 & n1406 ;
  assign n1535 = ( ~n1411 & n1533 ) | ( ~n1411 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = ( n1411 & n1533 ) | ( n1411 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1537 = ( n1411 & n1535 ) | ( n1411 & ~n1536 ) | ( n1535 & ~n1536 ) ;
  assign n1538 = ( x83 & n1532 ) | ( x83 & ~n1537 ) | ( n1532 & ~n1537 ) ;
  assign n1539 = n173 & n1185 ;
  assign n1540 = n1414 & n1539 ;
  assign n1541 = n389 | n1540 ;
  assign n1542 = ( x84 & ~n1424 ) | ( x84 & n1538 ) | ( ~n1424 & n1538 ) ;
  assign n1543 = ( x85 & ~n1541 ) | ( x85 & n1542 ) | ( ~n1541 & n1542 ) ;
  assign n1544 = n171 | n1543 ;
  assign n1545 = ( x84 & n1538 ) | ( x84 & n1544 ) | ( n1538 & n1544 ) ;
  assign n1546 = x84 | n1538 ;
  assign n1547 = ( ~n1424 & n1545 ) | ( ~n1424 & n1546 ) | ( n1545 & n1546 ) ;
  assign n1548 = ( n1424 & n1545 ) | ( n1424 & n1546 ) | ( n1545 & n1546 ) ;
  assign n1549 = ( n1424 & n1547 ) | ( n1424 & ~n1548 ) | ( n1547 & ~n1548 ) ;
  assign n1550 = ~x41 & x64 ;
  assign n1551 = ~x42 & n1544 ;
  assign n1552 = ( x42 & ~x64 ) | ( x42 & n1544 ) | ( ~x64 & n1544 ) ;
  assign n1553 = ( n1425 & ~n1551 ) | ( n1425 & n1552 ) | ( ~n1551 & n1552 ) ;
  assign n1554 = ( x65 & n1550 ) | ( x65 & ~n1553 ) | ( n1550 & ~n1553 ) ;
  assign n1555 = ( x65 & n1425 ) | ( x65 & n1544 ) | ( n1425 & n1544 ) ;
  assign n1556 = x65 | n1425 ;
  assign n1557 = ( ~n1429 & n1555 ) | ( ~n1429 & n1556 ) | ( n1555 & n1556 ) ;
  assign n1558 = ( n1429 & n1555 ) | ( n1429 & n1556 ) | ( n1555 & n1556 ) ;
  assign n1559 = ( n1429 & n1557 ) | ( n1429 & ~n1558 ) | ( n1557 & ~n1558 ) ;
  assign n1560 = ( x66 & n1554 ) | ( x66 & ~n1559 ) | ( n1554 & ~n1559 ) ;
  assign n1561 = ( x66 & n1430 ) | ( x66 & n1544 ) | ( n1430 & n1544 ) ;
  assign n1562 = x66 | n1430 ;
  assign n1563 = ( ~n1435 & n1561 ) | ( ~n1435 & n1562 ) | ( n1561 & n1562 ) ;
  assign n1564 = ( n1435 & n1561 ) | ( n1435 & n1562 ) | ( n1561 & n1562 ) ;
  assign n1565 = ( n1435 & n1563 ) | ( n1435 & ~n1564 ) | ( n1563 & ~n1564 ) ;
  assign n1566 = ( x67 & n1560 ) | ( x67 & ~n1565 ) | ( n1560 & ~n1565 ) ;
  assign n1567 = ( x67 & n1436 ) | ( x67 & ~n1544 ) | ( n1436 & ~n1544 ) ;
  assign n1568 = x67 & n1436 ;
  assign n1569 = ( ~n1441 & n1567 ) | ( ~n1441 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1570 = ( n1441 & n1567 ) | ( n1441 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1571 = ( n1441 & n1569 ) | ( n1441 & ~n1570 ) | ( n1569 & ~n1570 ) ;
  assign n1572 = ( x68 & n1566 ) | ( x68 & ~n1571 ) | ( n1566 & ~n1571 ) ;
  assign n1573 = ( x68 & n1442 ) | ( x68 & ~n1544 ) | ( n1442 & ~n1544 ) ;
  assign n1574 = x68 & n1442 ;
  assign n1575 = ( ~n1447 & n1573 ) | ( ~n1447 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1576 = ( n1447 & n1573 ) | ( n1447 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1577 = ( n1447 & n1575 ) | ( n1447 & ~n1576 ) | ( n1575 & ~n1576 ) ;
  assign n1578 = ( x69 & n1572 ) | ( x69 & ~n1577 ) | ( n1572 & ~n1577 ) ;
  assign n1579 = ( x69 & n1448 ) | ( x69 & ~n1544 ) | ( n1448 & ~n1544 ) ;
  assign n1580 = x69 & n1448 ;
  assign n1581 = ( ~n1453 & n1579 ) | ( ~n1453 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = ( n1453 & n1579 ) | ( n1453 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1583 = ( n1453 & n1581 ) | ( n1453 & ~n1582 ) | ( n1581 & ~n1582 ) ;
  assign n1584 = ( x70 & n1578 ) | ( x70 & ~n1583 ) | ( n1578 & ~n1583 ) ;
  assign n1585 = ( x70 & n1454 ) | ( x70 & ~n1544 ) | ( n1454 & ~n1544 ) ;
  assign n1586 = x70 & n1454 ;
  assign n1587 = ( ~n1459 & n1585 ) | ( ~n1459 & n1586 ) | ( n1585 & n1586 ) ;
  assign n1588 = ( n1459 & n1585 ) | ( n1459 & n1586 ) | ( n1585 & n1586 ) ;
  assign n1589 = ( n1459 & n1587 ) | ( n1459 & ~n1588 ) | ( n1587 & ~n1588 ) ;
  assign n1590 = ( x71 & n1584 ) | ( x71 & ~n1589 ) | ( n1584 & ~n1589 ) ;
  assign n1591 = ( x71 & n1460 ) | ( x71 & ~n1544 ) | ( n1460 & ~n1544 ) ;
  assign n1592 = x71 & n1460 ;
  assign n1593 = ( ~n1465 & n1591 ) | ( ~n1465 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = ( n1465 & n1591 ) | ( n1465 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1595 = ( n1465 & n1593 ) | ( n1465 & ~n1594 ) | ( n1593 & ~n1594 ) ;
  assign n1596 = ( x72 & n1590 ) | ( x72 & ~n1595 ) | ( n1590 & ~n1595 ) ;
  assign n1597 = ( x72 & n1466 ) | ( x72 & ~n1544 ) | ( n1466 & ~n1544 ) ;
  assign n1598 = x72 & n1466 ;
  assign n1599 = ( ~n1471 & n1597 ) | ( ~n1471 & n1598 ) | ( n1597 & n1598 ) ;
  assign n1600 = ( n1471 & n1597 ) | ( n1471 & n1598 ) | ( n1597 & n1598 ) ;
  assign n1601 = ( n1471 & n1599 ) | ( n1471 & ~n1600 ) | ( n1599 & ~n1600 ) ;
  assign n1602 = ( x73 & n1596 ) | ( x73 & ~n1601 ) | ( n1596 & ~n1601 ) ;
  assign n1603 = ( x73 & n1472 ) | ( x73 & ~n1544 ) | ( n1472 & ~n1544 ) ;
  assign n1604 = x73 & n1472 ;
  assign n1605 = ( ~n1477 & n1603 ) | ( ~n1477 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = ( n1477 & n1603 ) | ( n1477 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1607 = ( n1477 & n1605 ) | ( n1477 & ~n1606 ) | ( n1605 & ~n1606 ) ;
  assign n1608 = ( x74 & n1602 ) | ( x74 & ~n1607 ) | ( n1602 & ~n1607 ) ;
  assign n1609 = ( x74 & n1478 ) | ( x74 & ~n1544 ) | ( n1478 & ~n1544 ) ;
  assign n1610 = x74 & n1478 ;
  assign n1611 = ( ~n1483 & n1609 ) | ( ~n1483 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1612 = ( n1483 & n1609 ) | ( n1483 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1613 = ( n1483 & n1611 ) | ( n1483 & ~n1612 ) | ( n1611 & ~n1612 ) ;
  assign n1614 = ( x75 & n1608 ) | ( x75 & ~n1613 ) | ( n1608 & ~n1613 ) ;
  assign n1615 = ( x75 & n1484 ) | ( x75 & ~n1544 ) | ( n1484 & ~n1544 ) ;
  assign n1616 = x75 & n1484 ;
  assign n1617 = ( ~n1489 & n1615 ) | ( ~n1489 & n1616 ) | ( n1615 & n1616 ) ;
  assign n1618 = ( n1489 & n1615 ) | ( n1489 & n1616 ) | ( n1615 & n1616 ) ;
  assign n1619 = ( n1489 & n1617 ) | ( n1489 & ~n1618 ) | ( n1617 & ~n1618 ) ;
  assign n1620 = ( x76 & n1614 ) | ( x76 & ~n1619 ) | ( n1614 & ~n1619 ) ;
  assign n1621 = ( x76 & n1490 ) | ( x76 & ~n1544 ) | ( n1490 & ~n1544 ) ;
  assign n1622 = x76 & n1490 ;
  assign n1623 = ( ~n1495 & n1621 ) | ( ~n1495 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = ( n1495 & n1621 ) | ( n1495 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1625 = ( n1495 & n1623 ) | ( n1495 & ~n1624 ) | ( n1623 & ~n1624 ) ;
  assign n1626 = ( x77 & n1620 ) | ( x77 & ~n1625 ) | ( n1620 & ~n1625 ) ;
  assign n1627 = ( x77 & n1496 ) | ( x77 & ~n1544 ) | ( n1496 & ~n1544 ) ;
  assign n1628 = x77 & n1496 ;
  assign n1629 = ( ~n1501 & n1627 ) | ( ~n1501 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1630 = ( n1501 & n1627 ) | ( n1501 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1631 = ( n1501 & n1629 ) | ( n1501 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1632 = ( x78 & n1626 ) | ( x78 & ~n1631 ) | ( n1626 & ~n1631 ) ;
  assign n1633 = ( x78 & n1502 ) | ( x78 & ~n1544 ) | ( n1502 & ~n1544 ) ;
  assign n1634 = x78 & n1502 ;
  assign n1635 = ( ~n1507 & n1633 ) | ( ~n1507 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = ( n1507 & n1633 ) | ( n1507 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1637 = ( n1507 & n1635 ) | ( n1507 & ~n1636 ) | ( n1635 & ~n1636 ) ;
  assign n1638 = ( x79 & n1632 ) | ( x79 & ~n1637 ) | ( n1632 & ~n1637 ) ;
  assign n1639 = ( x79 & n1508 ) | ( x79 & ~n1544 ) | ( n1508 & ~n1544 ) ;
  assign n1640 = x79 & n1508 ;
  assign n1641 = ( ~n1513 & n1639 ) | ( ~n1513 & n1640 ) | ( n1639 & n1640 ) ;
  assign n1642 = ( n1513 & n1639 ) | ( n1513 & n1640 ) | ( n1639 & n1640 ) ;
  assign n1643 = ( n1513 & n1641 ) | ( n1513 & ~n1642 ) | ( n1641 & ~n1642 ) ;
  assign n1644 = ( x80 & n1638 ) | ( x80 & ~n1643 ) | ( n1638 & ~n1643 ) ;
  assign n1645 = ( x80 & n1514 ) | ( x80 & ~n1544 ) | ( n1514 & ~n1544 ) ;
  assign n1646 = x80 & n1514 ;
  assign n1647 = ( ~n1519 & n1645 ) | ( ~n1519 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = ( n1519 & n1645 ) | ( n1519 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1649 = ( n1519 & n1647 ) | ( n1519 & ~n1648 ) | ( n1647 & ~n1648 ) ;
  assign n1650 = ( x81 & n1644 ) | ( x81 & ~n1649 ) | ( n1644 & ~n1649 ) ;
  assign n1651 = ( x81 & n1520 ) | ( x81 & ~n1544 ) | ( n1520 & ~n1544 ) ;
  assign n1652 = x81 & n1520 ;
  assign n1653 = ( ~n1525 & n1651 ) | ( ~n1525 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1654 = ( n1525 & n1651 ) | ( n1525 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1655 = ( n1525 & n1653 ) | ( n1525 & ~n1654 ) | ( n1653 & ~n1654 ) ;
  assign n1656 = ( x82 & n1650 ) | ( x82 & ~n1655 ) | ( n1650 & ~n1655 ) ;
  assign n1657 = ( x82 & n1526 ) | ( x82 & ~n1544 ) | ( n1526 & ~n1544 ) ;
  assign n1658 = x82 & n1526 ;
  assign n1659 = ( ~n1531 & n1657 ) | ( ~n1531 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = ( n1531 & n1657 ) | ( n1531 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1661 = ( n1531 & n1659 ) | ( n1531 & ~n1660 ) | ( n1659 & ~n1660 ) ;
  assign n1662 = ( x83 & n1656 ) | ( x83 & ~n1661 ) | ( n1656 & ~n1661 ) ;
  assign n1663 = ( x83 & n1532 ) | ( x83 & ~n1544 ) | ( n1532 & ~n1544 ) ;
  assign n1664 = x83 & n1532 ;
  assign n1665 = ( ~n1537 & n1663 ) | ( ~n1537 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1666 = ( n1537 & n1663 ) | ( n1537 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1667 = ( n1537 & n1665 ) | ( n1537 & ~n1666 ) | ( n1665 & ~n1666 ) ;
  assign n1668 = ( x84 & n1662 ) | ( x84 & ~n1667 ) | ( n1662 & ~n1667 ) ;
  assign n1669 = ( x85 & n171 ) | ( x85 & n1542 ) | ( n171 & n1542 ) ;
  assign n1670 = x85 | n1542 ;
  assign n1671 = ( n1541 & n1669 ) | ( n1541 & ~n1670 ) | ( n1669 & ~n1670 ) ;
  assign n1672 = ( x85 & ~n1549 ) | ( x85 & n1668 ) | ( ~n1549 & n1668 ) ;
  assign n1673 = ( x86 & ~n1671 ) | ( x86 & n1672 ) | ( ~n1671 & n1672 ) ;
  assign n1674 = n170 | n1673 ;
  assign n1675 = ( x85 & n1668 ) | ( x85 & n1674 ) | ( n1668 & n1674 ) ;
  assign n1676 = x85 | n1668 ;
  assign n1677 = ( ~n1549 & n1675 ) | ( ~n1549 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1678 = ( n1549 & n1675 ) | ( n1549 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1679 = ( n1549 & n1677 ) | ( n1549 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n1680 = ~x40 & x64 ;
  assign n1681 = ~x41 & n1674 ;
  assign n1682 = ( x41 & ~x64 ) | ( x41 & n1674 ) | ( ~x64 & n1674 ) ;
  assign n1683 = ( n1550 & ~n1681 ) | ( n1550 & n1682 ) | ( ~n1681 & n1682 ) ;
  assign n1684 = ( x65 & n1680 ) | ( x65 & ~n1683 ) | ( n1680 & ~n1683 ) ;
  assign n1685 = ( x65 & n1550 ) | ( x65 & n1674 ) | ( n1550 & n1674 ) ;
  assign n1686 = x65 | n1550 ;
  assign n1687 = ( ~n1553 & n1685 ) | ( ~n1553 & n1686 ) | ( n1685 & n1686 ) ;
  assign n1688 = ( n1553 & n1685 ) | ( n1553 & n1686 ) | ( n1685 & n1686 ) ;
  assign n1689 = ( n1553 & n1687 ) | ( n1553 & ~n1688 ) | ( n1687 & ~n1688 ) ;
  assign n1690 = ( x66 & n1684 ) | ( x66 & ~n1689 ) | ( n1684 & ~n1689 ) ;
  assign n1691 = ( x66 & n1554 ) | ( x66 & n1674 ) | ( n1554 & n1674 ) ;
  assign n1692 = x66 | n1554 ;
  assign n1693 = ( ~n1559 & n1691 ) | ( ~n1559 & n1692 ) | ( n1691 & n1692 ) ;
  assign n1694 = ( n1559 & n1691 ) | ( n1559 & n1692 ) | ( n1691 & n1692 ) ;
  assign n1695 = ( n1559 & n1693 ) | ( n1559 & ~n1694 ) | ( n1693 & ~n1694 ) ;
  assign n1696 = ( x67 & n1690 ) | ( x67 & ~n1695 ) | ( n1690 & ~n1695 ) ;
  assign n1697 = ( x67 & n1560 ) | ( x67 & ~n1674 ) | ( n1560 & ~n1674 ) ;
  assign n1698 = x67 & n1560 ;
  assign n1699 = ( ~n1565 & n1697 ) | ( ~n1565 & n1698 ) | ( n1697 & n1698 ) ;
  assign n1700 = ( n1565 & n1697 ) | ( n1565 & n1698 ) | ( n1697 & n1698 ) ;
  assign n1701 = ( n1565 & n1699 ) | ( n1565 & ~n1700 ) | ( n1699 & ~n1700 ) ;
  assign n1702 = ( x68 & n1696 ) | ( x68 & ~n1701 ) | ( n1696 & ~n1701 ) ;
  assign n1703 = ( x68 & n1566 ) | ( x68 & ~n1674 ) | ( n1566 & ~n1674 ) ;
  assign n1704 = x68 & n1566 ;
  assign n1705 = ( ~n1571 & n1703 ) | ( ~n1571 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ( n1571 & n1703 ) | ( n1571 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1707 = ( n1571 & n1705 ) | ( n1571 & ~n1706 ) | ( n1705 & ~n1706 ) ;
  assign n1708 = ( x69 & n1702 ) | ( x69 & ~n1707 ) | ( n1702 & ~n1707 ) ;
  assign n1709 = ( x69 & n1572 ) | ( x69 & ~n1674 ) | ( n1572 & ~n1674 ) ;
  assign n1710 = x69 & n1572 ;
  assign n1711 = ( ~n1577 & n1709 ) | ( ~n1577 & n1710 ) | ( n1709 & n1710 ) ;
  assign n1712 = ( n1577 & n1709 ) | ( n1577 & n1710 ) | ( n1709 & n1710 ) ;
  assign n1713 = ( n1577 & n1711 ) | ( n1577 & ~n1712 ) | ( n1711 & ~n1712 ) ;
  assign n1714 = ( x70 & n1708 ) | ( x70 & ~n1713 ) | ( n1708 & ~n1713 ) ;
  assign n1715 = ( x70 & n1578 ) | ( x70 & ~n1674 ) | ( n1578 & ~n1674 ) ;
  assign n1716 = x70 & n1578 ;
  assign n1717 = ( ~n1583 & n1715 ) | ( ~n1583 & n1716 ) | ( n1715 & n1716 ) ;
  assign n1718 = ( n1583 & n1715 ) | ( n1583 & n1716 ) | ( n1715 & n1716 ) ;
  assign n1719 = ( n1583 & n1717 ) | ( n1583 & ~n1718 ) | ( n1717 & ~n1718 ) ;
  assign n1720 = ( x71 & n1714 ) | ( x71 & ~n1719 ) | ( n1714 & ~n1719 ) ;
  assign n1721 = ( x71 & n1584 ) | ( x71 & ~n1674 ) | ( n1584 & ~n1674 ) ;
  assign n1722 = x71 & n1584 ;
  assign n1723 = ( ~n1589 & n1721 ) | ( ~n1589 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1724 = ( n1589 & n1721 ) | ( n1589 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1725 = ( n1589 & n1723 ) | ( n1589 & ~n1724 ) | ( n1723 & ~n1724 ) ;
  assign n1726 = ( x72 & n1720 ) | ( x72 & ~n1725 ) | ( n1720 & ~n1725 ) ;
  assign n1727 = ( x72 & n1590 ) | ( x72 & ~n1674 ) | ( n1590 & ~n1674 ) ;
  assign n1728 = x72 & n1590 ;
  assign n1729 = ( ~n1595 & n1727 ) | ( ~n1595 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = ( n1595 & n1727 ) | ( n1595 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1731 = ( n1595 & n1729 ) | ( n1595 & ~n1730 ) | ( n1729 & ~n1730 ) ;
  assign n1732 = ( x73 & n1726 ) | ( x73 & ~n1731 ) | ( n1726 & ~n1731 ) ;
  assign n1733 = ( x73 & n1596 ) | ( x73 & ~n1674 ) | ( n1596 & ~n1674 ) ;
  assign n1734 = x73 & n1596 ;
  assign n1735 = ( ~n1601 & n1733 ) | ( ~n1601 & n1734 ) | ( n1733 & n1734 ) ;
  assign n1736 = ( n1601 & n1733 ) | ( n1601 & n1734 ) | ( n1733 & n1734 ) ;
  assign n1737 = ( n1601 & n1735 ) | ( n1601 & ~n1736 ) | ( n1735 & ~n1736 ) ;
  assign n1738 = ( x74 & n1732 ) | ( x74 & ~n1737 ) | ( n1732 & ~n1737 ) ;
  assign n1739 = ( x74 & n1602 ) | ( x74 & ~n1674 ) | ( n1602 & ~n1674 ) ;
  assign n1740 = x74 & n1602 ;
  assign n1741 = ( ~n1607 & n1739 ) | ( ~n1607 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1742 = ( n1607 & n1739 ) | ( n1607 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1743 = ( n1607 & n1741 ) | ( n1607 & ~n1742 ) | ( n1741 & ~n1742 ) ;
  assign n1744 = ( x75 & n1738 ) | ( x75 & ~n1743 ) | ( n1738 & ~n1743 ) ;
  assign n1745 = ( x75 & n1608 ) | ( x75 & ~n1674 ) | ( n1608 & ~n1674 ) ;
  assign n1746 = x75 & n1608 ;
  assign n1747 = ( ~n1613 & n1745 ) | ( ~n1613 & n1746 ) | ( n1745 & n1746 ) ;
  assign n1748 = ( n1613 & n1745 ) | ( n1613 & n1746 ) | ( n1745 & n1746 ) ;
  assign n1749 = ( n1613 & n1747 ) | ( n1613 & ~n1748 ) | ( n1747 & ~n1748 ) ;
  assign n1750 = ( x76 & n1744 ) | ( x76 & ~n1749 ) | ( n1744 & ~n1749 ) ;
  assign n1751 = ( x76 & n1614 ) | ( x76 & ~n1674 ) | ( n1614 & ~n1674 ) ;
  assign n1752 = x76 & n1614 ;
  assign n1753 = ( ~n1619 & n1751 ) | ( ~n1619 & n1752 ) | ( n1751 & n1752 ) ;
  assign n1754 = ( n1619 & n1751 ) | ( n1619 & n1752 ) | ( n1751 & n1752 ) ;
  assign n1755 = ( n1619 & n1753 ) | ( n1619 & ~n1754 ) | ( n1753 & ~n1754 ) ;
  assign n1756 = ( x77 & n1750 ) | ( x77 & ~n1755 ) | ( n1750 & ~n1755 ) ;
  assign n1757 = ( x77 & n1620 ) | ( x77 & ~n1674 ) | ( n1620 & ~n1674 ) ;
  assign n1758 = x77 & n1620 ;
  assign n1759 = ( ~n1625 & n1757 ) | ( ~n1625 & n1758 ) | ( n1757 & n1758 ) ;
  assign n1760 = ( n1625 & n1757 ) | ( n1625 & n1758 ) | ( n1757 & n1758 ) ;
  assign n1761 = ( n1625 & n1759 ) | ( n1625 & ~n1760 ) | ( n1759 & ~n1760 ) ;
  assign n1762 = ( x78 & n1756 ) | ( x78 & ~n1761 ) | ( n1756 & ~n1761 ) ;
  assign n1763 = ( x78 & n1626 ) | ( x78 & ~n1674 ) | ( n1626 & ~n1674 ) ;
  assign n1764 = x78 & n1626 ;
  assign n1765 = ( ~n1631 & n1763 ) | ( ~n1631 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1766 = ( n1631 & n1763 ) | ( n1631 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1767 = ( n1631 & n1765 ) | ( n1631 & ~n1766 ) | ( n1765 & ~n1766 ) ;
  assign n1768 = ( x79 & n1762 ) | ( x79 & ~n1767 ) | ( n1762 & ~n1767 ) ;
  assign n1769 = ( x79 & n1632 ) | ( x79 & ~n1674 ) | ( n1632 & ~n1674 ) ;
  assign n1770 = x79 & n1632 ;
  assign n1771 = ( ~n1637 & n1769 ) | ( ~n1637 & n1770 ) | ( n1769 & n1770 ) ;
  assign n1772 = ( n1637 & n1769 ) | ( n1637 & n1770 ) | ( n1769 & n1770 ) ;
  assign n1773 = ( n1637 & n1771 ) | ( n1637 & ~n1772 ) | ( n1771 & ~n1772 ) ;
  assign n1774 = ( x80 & n1768 ) | ( x80 & ~n1773 ) | ( n1768 & ~n1773 ) ;
  assign n1775 = ( x80 & n1638 ) | ( x80 & ~n1674 ) | ( n1638 & ~n1674 ) ;
  assign n1776 = x80 & n1638 ;
  assign n1777 = ( ~n1643 & n1775 ) | ( ~n1643 & n1776 ) | ( n1775 & n1776 ) ;
  assign n1778 = ( n1643 & n1775 ) | ( n1643 & n1776 ) | ( n1775 & n1776 ) ;
  assign n1779 = ( n1643 & n1777 ) | ( n1643 & ~n1778 ) | ( n1777 & ~n1778 ) ;
  assign n1780 = ( x81 & n1774 ) | ( x81 & ~n1779 ) | ( n1774 & ~n1779 ) ;
  assign n1781 = ( x81 & n1644 ) | ( x81 & ~n1674 ) | ( n1644 & ~n1674 ) ;
  assign n1782 = x81 & n1644 ;
  assign n1783 = ( ~n1649 & n1781 ) | ( ~n1649 & n1782 ) | ( n1781 & n1782 ) ;
  assign n1784 = ( n1649 & n1781 ) | ( n1649 & n1782 ) | ( n1781 & n1782 ) ;
  assign n1785 = ( n1649 & n1783 ) | ( n1649 & ~n1784 ) | ( n1783 & ~n1784 ) ;
  assign n1786 = ( x82 & n1780 ) | ( x82 & ~n1785 ) | ( n1780 & ~n1785 ) ;
  assign n1787 = ( x82 & n1650 ) | ( x82 & ~n1674 ) | ( n1650 & ~n1674 ) ;
  assign n1788 = x82 & n1650 ;
  assign n1789 = ( ~n1655 & n1787 ) | ( ~n1655 & n1788 ) | ( n1787 & n1788 ) ;
  assign n1790 = ( n1655 & n1787 ) | ( n1655 & n1788 ) | ( n1787 & n1788 ) ;
  assign n1791 = ( n1655 & n1789 ) | ( n1655 & ~n1790 ) | ( n1789 & ~n1790 ) ;
  assign n1792 = ( x83 & n1786 ) | ( x83 & ~n1791 ) | ( n1786 & ~n1791 ) ;
  assign n1793 = ( x83 & n1656 ) | ( x83 & ~n1674 ) | ( n1656 & ~n1674 ) ;
  assign n1794 = x83 & n1656 ;
  assign n1795 = ( ~n1661 & n1793 ) | ( ~n1661 & n1794 ) | ( n1793 & n1794 ) ;
  assign n1796 = ( n1661 & n1793 ) | ( n1661 & n1794 ) | ( n1793 & n1794 ) ;
  assign n1797 = ( n1661 & n1795 ) | ( n1661 & ~n1796 ) | ( n1795 & ~n1796 ) ;
  assign n1798 = ( x84 & n1792 ) | ( x84 & ~n1797 ) | ( n1792 & ~n1797 ) ;
  assign n1799 = ( x84 & n1662 ) | ( x84 & ~n1674 ) | ( n1662 & ~n1674 ) ;
  assign n1800 = x84 & n1662 ;
  assign n1801 = ( ~n1667 & n1799 ) | ( ~n1667 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1802 = ( n1667 & n1799 ) | ( n1667 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1803 = ( n1667 & n1801 ) | ( n1667 & ~n1802 ) | ( n1801 & ~n1802 ) ;
  assign n1804 = ( x85 & n1798 ) | ( x85 & ~n1803 ) | ( n1798 & ~n1803 ) ;
  assign n1805 = ( x86 & ~n1679 ) | ( x86 & n1804 ) | ( ~n1679 & n1804 ) ;
  assign n1806 = n169 | n1805 ;
  assign n1807 = x87 & ~n1671 ;
  assign n1808 = x86 & ~n170 ;
  assign n1809 = n1540 & n1808 ;
  assign n1810 = n1672 & n1809 ;
  assign n1811 = ~n1807 & n1810 ;
  assign n1812 = ( n1806 & n1807 ) | ( n1806 & ~n1811 ) | ( n1807 & ~n1811 ) ;
  assign n1813 = ( x86 & n1804 ) | ( x86 & n1812 ) | ( n1804 & n1812 ) ;
  assign n1814 = x86 | n1804 ;
  assign n1815 = ( ~n1679 & n1813 ) | ( ~n1679 & n1814 ) | ( n1813 & n1814 ) ;
  assign n1816 = ( n1679 & n1813 ) | ( n1679 & n1814 ) | ( n1813 & n1814 ) ;
  assign n1817 = ( n1679 & n1815 ) | ( n1679 & ~n1816 ) | ( n1815 & ~n1816 ) ;
  assign n1818 = ~x39 & x64 ;
  assign n1819 = ~x40 & n1812 ;
  assign n1820 = ( x40 & ~x64 ) | ( x40 & n1812 ) | ( ~x64 & n1812 ) ;
  assign n1821 = ( n1680 & ~n1819 ) | ( n1680 & n1820 ) | ( ~n1819 & n1820 ) ;
  assign n1822 = ( x65 & n1818 ) | ( x65 & ~n1821 ) | ( n1818 & ~n1821 ) ;
  assign n1823 = ( x65 & n1680 ) | ( x65 & n1812 ) | ( n1680 & n1812 ) ;
  assign n1824 = x65 | n1680 ;
  assign n1825 = ( ~n1683 & n1823 ) | ( ~n1683 & n1824 ) | ( n1823 & n1824 ) ;
  assign n1826 = ( n1683 & n1823 ) | ( n1683 & n1824 ) | ( n1823 & n1824 ) ;
  assign n1827 = ( n1683 & n1825 ) | ( n1683 & ~n1826 ) | ( n1825 & ~n1826 ) ;
  assign n1828 = ( x66 & n1822 ) | ( x66 & ~n1827 ) | ( n1822 & ~n1827 ) ;
  assign n1829 = ( x66 & n1684 ) | ( x66 & n1812 ) | ( n1684 & n1812 ) ;
  assign n1830 = x66 | n1684 ;
  assign n1831 = ( ~n1689 & n1829 ) | ( ~n1689 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1832 = ( n1689 & n1829 ) | ( n1689 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1833 = ( n1689 & n1831 ) | ( n1689 & ~n1832 ) | ( n1831 & ~n1832 ) ;
  assign n1834 = ( x67 & n1828 ) | ( x67 & ~n1833 ) | ( n1828 & ~n1833 ) ;
  assign n1835 = ( x67 & n1690 ) | ( x67 & ~n1812 ) | ( n1690 & ~n1812 ) ;
  assign n1836 = x67 & n1690 ;
  assign n1837 = ( ~n1695 & n1835 ) | ( ~n1695 & n1836 ) | ( n1835 & n1836 ) ;
  assign n1838 = ( n1695 & n1835 ) | ( n1695 & n1836 ) | ( n1835 & n1836 ) ;
  assign n1839 = ( n1695 & n1837 ) | ( n1695 & ~n1838 ) | ( n1837 & ~n1838 ) ;
  assign n1840 = ( x68 & n1834 ) | ( x68 & ~n1839 ) | ( n1834 & ~n1839 ) ;
  assign n1841 = ( x68 & n1696 ) | ( x68 & ~n1812 ) | ( n1696 & ~n1812 ) ;
  assign n1842 = x68 & n1696 ;
  assign n1843 = ( ~n1701 & n1841 ) | ( ~n1701 & n1842 ) | ( n1841 & n1842 ) ;
  assign n1844 = ( n1701 & n1841 ) | ( n1701 & n1842 ) | ( n1841 & n1842 ) ;
  assign n1845 = ( n1701 & n1843 ) | ( n1701 & ~n1844 ) | ( n1843 & ~n1844 ) ;
  assign n1846 = ( x69 & n1840 ) | ( x69 & ~n1845 ) | ( n1840 & ~n1845 ) ;
  assign n1847 = ( x69 & n1702 ) | ( x69 & ~n1812 ) | ( n1702 & ~n1812 ) ;
  assign n1848 = x69 & n1702 ;
  assign n1849 = ( ~n1707 & n1847 ) | ( ~n1707 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1850 = ( n1707 & n1847 ) | ( n1707 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1851 = ( n1707 & n1849 ) | ( n1707 & ~n1850 ) | ( n1849 & ~n1850 ) ;
  assign n1852 = ( x70 & n1846 ) | ( x70 & ~n1851 ) | ( n1846 & ~n1851 ) ;
  assign n1853 = ( x70 & n1708 ) | ( x70 & ~n1812 ) | ( n1708 & ~n1812 ) ;
  assign n1854 = x70 & n1708 ;
  assign n1855 = ( ~n1713 & n1853 ) | ( ~n1713 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1856 = ( n1713 & n1853 ) | ( n1713 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1857 = ( n1713 & n1855 ) | ( n1713 & ~n1856 ) | ( n1855 & ~n1856 ) ;
  assign n1858 = ( x71 & n1852 ) | ( x71 & ~n1857 ) | ( n1852 & ~n1857 ) ;
  assign n1859 = ( x71 & n1714 ) | ( x71 & ~n1812 ) | ( n1714 & ~n1812 ) ;
  assign n1860 = x71 & n1714 ;
  assign n1861 = ( ~n1719 & n1859 ) | ( ~n1719 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1862 = ( n1719 & n1859 ) | ( n1719 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1863 = ( n1719 & n1861 ) | ( n1719 & ~n1862 ) | ( n1861 & ~n1862 ) ;
  assign n1864 = ( x72 & n1858 ) | ( x72 & ~n1863 ) | ( n1858 & ~n1863 ) ;
  assign n1865 = ( x72 & n1720 ) | ( x72 & ~n1812 ) | ( n1720 & ~n1812 ) ;
  assign n1866 = x72 & n1720 ;
  assign n1867 = ( ~n1725 & n1865 ) | ( ~n1725 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1868 = ( n1725 & n1865 ) | ( n1725 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1869 = ( n1725 & n1867 ) | ( n1725 & ~n1868 ) | ( n1867 & ~n1868 ) ;
  assign n1870 = ( x73 & n1864 ) | ( x73 & ~n1869 ) | ( n1864 & ~n1869 ) ;
  assign n1871 = ( x73 & n1726 ) | ( x73 & ~n1812 ) | ( n1726 & ~n1812 ) ;
  assign n1872 = x73 & n1726 ;
  assign n1873 = ( ~n1731 & n1871 ) | ( ~n1731 & n1872 ) | ( n1871 & n1872 ) ;
  assign n1874 = ( n1731 & n1871 ) | ( n1731 & n1872 ) | ( n1871 & n1872 ) ;
  assign n1875 = ( n1731 & n1873 ) | ( n1731 & ~n1874 ) | ( n1873 & ~n1874 ) ;
  assign n1876 = ( x74 & n1870 ) | ( x74 & ~n1875 ) | ( n1870 & ~n1875 ) ;
  assign n1877 = ( x74 & n1732 ) | ( x74 & ~n1812 ) | ( n1732 & ~n1812 ) ;
  assign n1878 = x74 & n1732 ;
  assign n1879 = ( ~n1737 & n1877 ) | ( ~n1737 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1880 = ( n1737 & n1877 ) | ( n1737 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1881 = ( n1737 & n1879 ) | ( n1737 & ~n1880 ) | ( n1879 & ~n1880 ) ;
  assign n1882 = ( x75 & n1876 ) | ( x75 & ~n1881 ) | ( n1876 & ~n1881 ) ;
  assign n1883 = ( x75 & n1738 ) | ( x75 & ~n1812 ) | ( n1738 & ~n1812 ) ;
  assign n1884 = x75 & n1738 ;
  assign n1885 = ( ~n1743 & n1883 ) | ( ~n1743 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1886 = ( n1743 & n1883 ) | ( n1743 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1887 = ( n1743 & n1885 ) | ( n1743 & ~n1886 ) | ( n1885 & ~n1886 ) ;
  assign n1888 = ( x76 & n1882 ) | ( x76 & ~n1887 ) | ( n1882 & ~n1887 ) ;
  assign n1889 = ( x76 & n1744 ) | ( x76 & ~n1812 ) | ( n1744 & ~n1812 ) ;
  assign n1890 = x76 & n1744 ;
  assign n1891 = ( ~n1749 & n1889 ) | ( ~n1749 & n1890 ) | ( n1889 & n1890 ) ;
  assign n1892 = ( n1749 & n1889 ) | ( n1749 & n1890 ) | ( n1889 & n1890 ) ;
  assign n1893 = ( n1749 & n1891 ) | ( n1749 & ~n1892 ) | ( n1891 & ~n1892 ) ;
  assign n1894 = ( x77 & n1888 ) | ( x77 & ~n1893 ) | ( n1888 & ~n1893 ) ;
  assign n1895 = ( x77 & n1750 ) | ( x77 & ~n1812 ) | ( n1750 & ~n1812 ) ;
  assign n1896 = x77 & n1750 ;
  assign n1897 = ( ~n1755 & n1895 ) | ( ~n1755 & n1896 ) | ( n1895 & n1896 ) ;
  assign n1898 = ( n1755 & n1895 ) | ( n1755 & n1896 ) | ( n1895 & n1896 ) ;
  assign n1899 = ( n1755 & n1897 ) | ( n1755 & ~n1898 ) | ( n1897 & ~n1898 ) ;
  assign n1900 = ( x78 & n1894 ) | ( x78 & ~n1899 ) | ( n1894 & ~n1899 ) ;
  assign n1901 = ( x78 & n1756 ) | ( x78 & ~n1812 ) | ( n1756 & ~n1812 ) ;
  assign n1902 = x78 & n1756 ;
  assign n1903 = ( ~n1761 & n1901 ) | ( ~n1761 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = ( n1761 & n1901 ) | ( n1761 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1905 = ( n1761 & n1903 ) | ( n1761 & ~n1904 ) | ( n1903 & ~n1904 ) ;
  assign n1906 = ( x79 & n1900 ) | ( x79 & ~n1905 ) | ( n1900 & ~n1905 ) ;
  assign n1907 = ( x79 & n1762 ) | ( x79 & ~n1812 ) | ( n1762 & ~n1812 ) ;
  assign n1908 = x79 & n1762 ;
  assign n1909 = ( ~n1767 & n1907 ) | ( ~n1767 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1910 = ( n1767 & n1907 ) | ( n1767 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1911 = ( n1767 & n1909 ) | ( n1767 & ~n1910 ) | ( n1909 & ~n1910 ) ;
  assign n1912 = ( x80 & n1906 ) | ( x80 & ~n1911 ) | ( n1906 & ~n1911 ) ;
  assign n1913 = ( x80 & n1768 ) | ( x80 & ~n1812 ) | ( n1768 & ~n1812 ) ;
  assign n1914 = x80 & n1768 ;
  assign n1915 = ( ~n1773 & n1913 ) | ( ~n1773 & n1914 ) | ( n1913 & n1914 ) ;
  assign n1916 = ( n1773 & n1913 ) | ( n1773 & n1914 ) | ( n1913 & n1914 ) ;
  assign n1917 = ( n1773 & n1915 ) | ( n1773 & ~n1916 ) | ( n1915 & ~n1916 ) ;
  assign n1918 = ( x81 & n1912 ) | ( x81 & ~n1917 ) | ( n1912 & ~n1917 ) ;
  assign n1919 = ( x81 & n1774 ) | ( x81 & ~n1812 ) | ( n1774 & ~n1812 ) ;
  assign n1920 = x81 & n1774 ;
  assign n1921 = ( ~n1779 & n1919 ) | ( ~n1779 & n1920 ) | ( n1919 & n1920 ) ;
  assign n1922 = ( n1779 & n1919 ) | ( n1779 & n1920 ) | ( n1919 & n1920 ) ;
  assign n1923 = ( n1779 & n1921 ) | ( n1779 & ~n1922 ) | ( n1921 & ~n1922 ) ;
  assign n1924 = ( x82 & n1918 ) | ( x82 & ~n1923 ) | ( n1918 & ~n1923 ) ;
  assign n1925 = ( x82 & n1780 ) | ( x82 & ~n1812 ) | ( n1780 & ~n1812 ) ;
  assign n1926 = x82 & n1780 ;
  assign n1927 = ( ~n1785 & n1925 ) | ( ~n1785 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1928 = ( n1785 & n1925 ) | ( n1785 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1929 = ( n1785 & n1927 ) | ( n1785 & ~n1928 ) | ( n1927 & ~n1928 ) ;
  assign n1930 = ( x83 & n1924 ) | ( x83 & ~n1929 ) | ( n1924 & ~n1929 ) ;
  assign n1931 = ( x83 & n1786 ) | ( x83 & ~n1812 ) | ( n1786 & ~n1812 ) ;
  assign n1932 = x83 & n1786 ;
  assign n1933 = ( ~n1791 & n1931 ) | ( ~n1791 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1934 = ( n1791 & n1931 ) | ( n1791 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1935 = ( n1791 & n1933 ) | ( n1791 & ~n1934 ) | ( n1933 & ~n1934 ) ;
  assign n1936 = ( x84 & n1930 ) | ( x84 & ~n1935 ) | ( n1930 & ~n1935 ) ;
  assign n1937 = ( x84 & n1792 ) | ( x84 & ~n1812 ) | ( n1792 & ~n1812 ) ;
  assign n1938 = x84 & n1792 ;
  assign n1939 = ( ~n1797 & n1937 ) | ( ~n1797 & n1938 ) | ( n1937 & n1938 ) ;
  assign n1940 = ( n1797 & n1937 ) | ( n1797 & n1938 ) | ( n1937 & n1938 ) ;
  assign n1941 = ( n1797 & n1939 ) | ( n1797 & ~n1940 ) | ( n1939 & ~n1940 ) ;
  assign n1942 = ( x85 & n1936 ) | ( x85 & ~n1941 ) | ( n1936 & ~n1941 ) ;
  assign n1943 = ( x85 & n1798 ) | ( x85 & ~n1812 ) | ( n1798 & ~n1812 ) ;
  assign n1944 = x85 & n1798 ;
  assign n1945 = ( ~n1803 & n1943 ) | ( ~n1803 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1946 = ( n1803 & n1943 ) | ( n1803 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1947 = ( n1803 & n1945 ) | ( n1803 & ~n1946 ) | ( n1945 & ~n1946 ) ;
  assign n1948 = ( x86 & n1942 ) | ( x86 & ~n1947 ) | ( n1942 & ~n1947 ) ;
  assign n1949 = ( x87 & ~n1817 ) | ( x87 & n1948 ) | ( ~n1817 & n1948 ) ;
  assign n1950 = ( n170 & n389 ) | ( n170 & n1541 ) | ( n389 & n1541 ) ;
  assign n1951 = ( n389 & n1806 ) | ( n389 & n1950 ) | ( n1806 & n1950 ) ;
  assign n1952 = ( x88 & n1949 ) | ( x88 & ~n1951 ) | ( n1949 & ~n1951 ) ;
  assign n1953 = n168 | n1952 ;
  assign n1954 = ( x87 & n1948 ) | ( x87 & n1953 ) | ( n1948 & n1953 ) ;
  assign n1955 = x87 | n1948 ;
  assign n1956 = ( ~n1817 & n1954 ) | ( ~n1817 & n1955 ) | ( n1954 & n1955 ) ;
  assign n1957 = ( n1817 & n1954 ) | ( n1817 & n1955 ) | ( n1954 & n1955 ) ;
  assign n1958 = ( n1817 & n1956 ) | ( n1817 & ~n1957 ) | ( n1956 & ~n1957 ) ;
  assign n1959 = ~x38 & x64 ;
  assign n1960 = ~x39 & n1953 ;
  assign n1961 = ( x39 & ~x64 ) | ( x39 & n1953 ) | ( ~x64 & n1953 ) ;
  assign n1962 = ( n1818 & ~n1960 ) | ( n1818 & n1961 ) | ( ~n1960 & n1961 ) ;
  assign n1963 = ( x65 & n1959 ) | ( x65 & ~n1962 ) | ( n1959 & ~n1962 ) ;
  assign n1964 = ( x65 & n1818 ) | ( x65 & n1953 ) | ( n1818 & n1953 ) ;
  assign n1965 = x65 | n1818 ;
  assign n1966 = ( ~n1821 & n1964 ) | ( ~n1821 & n1965 ) | ( n1964 & n1965 ) ;
  assign n1967 = ( n1821 & n1964 ) | ( n1821 & n1965 ) | ( n1964 & n1965 ) ;
  assign n1968 = ( n1821 & n1966 ) | ( n1821 & ~n1967 ) | ( n1966 & ~n1967 ) ;
  assign n1969 = ( x66 & n1963 ) | ( x66 & ~n1968 ) | ( n1963 & ~n1968 ) ;
  assign n1970 = ( x66 & n1822 ) | ( x66 & n1953 ) | ( n1822 & n1953 ) ;
  assign n1971 = x66 | n1822 ;
  assign n1972 = ( ~n1827 & n1970 ) | ( ~n1827 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1973 = ( n1827 & n1970 ) | ( n1827 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1974 = ( n1827 & n1972 ) | ( n1827 & ~n1973 ) | ( n1972 & ~n1973 ) ;
  assign n1975 = ( x67 & n1969 ) | ( x67 & ~n1974 ) | ( n1969 & ~n1974 ) ;
  assign n1976 = ( x67 & n1828 ) | ( x67 & ~n1953 ) | ( n1828 & ~n1953 ) ;
  assign n1977 = x67 & n1828 ;
  assign n1978 = ( ~n1833 & n1976 ) | ( ~n1833 & n1977 ) | ( n1976 & n1977 ) ;
  assign n1979 = ( n1833 & n1976 ) | ( n1833 & n1977 ) | ( n1976 & n1977 ) ;
  assign n1980 = ( n1833 & n1978 ) | ( n1833 & ~n1979 ) | ( n1978 & ~n1979 ) ;
  assign n1981 = ( x68 & n1975 ) | ( x68 & ~n1980 ) | ( n1975 & ~n1980 ) ;
  assign n1982 = ( x68 & n1834 ) | ( x68 & ~n1953 ) | ( n1834 & ~n1953 ) ;
  assign n1983 = x68 & n1834 ;
  assign n1984 = ( ~n1839 & n1982 ) | ( ~n1839 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1985 = ( n1839 & n1982 ) | ( n1839 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1986 = ( n1839 & n1984 ) | ( n1839 & ~n1985 ) | ( n1984 & ~n1985 ) ;
  assign n1987 = ( x69 & n1981 ) | ( x69 & ~n1986 ) | ( n1981 & ~n1986 ) ;
  assign n1988 = ( x69 & n1840 ) | ( x69 & ~n1953 ) | ( n1840 & ~n1953 ) ;
  assign n1989 = x69 & n1840 ;
  assign n1990 = ( ~n1845 & n1988 ) | ( ~n1845 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1991 = ( n1845 & n1988 ) | ( n1845 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1992 = ( n1845 & n1990 ) | ( n1845 & ~n1991 ) | ( n1990 & ~n1991 ) ;
  assign n1993 = ( x70 & n1987 ) | ( x70 & ~n1992 ) | ( n1987 & ~n1992 ) ;
  assign n1994 = ( x70 & n1846 ) | ( x70 & ~n1953 ) | ( n1846 & ~n1953 ) ;
  assign n1995 = x70 & n1846 ;
  assign n1996 = ( ~n1851 & n1994 ) | ( ~n1851 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1997 = ( n1851 & n1994 ) | ( n1851 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1998 = ( n1851 & n1996 ) | ( n1851 & ~n1997 ) | ( n1996 & ~n1997 ) ;
  assign n1999 = ( x71 & n1993 ) | ( x71 & ~n1998 ) | ( n1993 & ~n1998 ) ;
  assign n2000 = ( x71 & n1852 ) | ( x71 & ~n1953 ) | ( n1852 & ~n1953 ) ;
  assign n2001 = x71 & n1852 ;
  assign n2002 = ( ~n1857 & n2000 ) | ( ~n1857 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2003 = ( n1857 & n2000 ) | ( n1857 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2004 = ( n1857 & n2002 ) | ( n1857 & ~n2003 ) | ( n2002 & ~n2003 ) ;
  assign n2005 = ( x72 & n1999 ) | ( x72 & ~n2004 ) | ( n1999 & ~n2004 ) ;
  assign n2006 = ( x72 & n1858 ) | ( x72 & ~n1953 ) | ( n1858 & ~n1953 ) ;
  assign n2007 = x72 & n1858 ;
  assign n2008 = ( ~n1863 & n2006 ) | ( ~n1863 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = ( n1863 & n2006 ) | ( n1863 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2010 = ( n1863 & n2008 ) | ( n1863 & ~n2009 ) | ( n2008 & ~n2009 ) ;
  assign n2011 = ( x73 & n2005 ) | ( x73 & ~n2010 ) | ( n2005 & ~n2010 ) ;
  assign n2012 = ( x73 & n1864 ) | ( x73 & ~n1953 ) | ( n1864 & ~n1953 ) ;
  assign n2013 = x73 & n1864 ;
  assign n2014 = ( ~n1869 & n2012 ) | ( ~n1869 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2015 = ( n1869 & n2012 ) | ( n1869 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2016 = ( n1869 & n2014 ) | ( n1869 & ~n2015 ) | ( n2014 & ~n2015 ) ;
  assign n2017 = ( x74 & n2011 ) | ( x74 & ~n2016 ) | ( n2011 & ~n2016 ) ;
  assign n2018 = ( x74 & n1870 ) | ( x74 & ~n1953 ) | ( n1870 & ~n1953 ) ;
  assign n2019 = x74 & n1870 ;
  assign n2020 = ( ~n1875 & n2018 ) | ( ~n1875 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2021 = ( n1875 & n2018 ) | ( n1875 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2022 = ( n1875 & n2020 ) | ( n1875 & ~n2021 ) | ( n2020 & ~n2021 ) ;
  assign n2023 = ( x75 & n2017 ) | ( x75 & ~n2022 ) | ( n2017 & ~n2022 ) ;
  assign n2024 = ( x75 & n1876 ) | ( x75 & ~n1953 ) | ( n1876 & ~n1953 ) ;
  assign n2025 = x75 & n1876 ;
  assign n2026 = ( ~n1881 & n2024 ) | ( ~n1881 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2027 = ( n1881 & n2024 ) | ( n1881 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2028 = ( n1881 & n2026 ) | ( n1881 & ~n2027 ) | ( n2026 & ~n2027 ) ;
  assign n2029 = ( x76 & n2023 ) | ( x76 & ~n2028 ) | ( n2023 & ~n2028 ) ;
  assign n2030 = ( x76 & n1882 ) | ( x76 & ~n1953 ) | ( n1882 & ~n1953 ) ;
  assign n2031 = x76 & n1882 ;
  assign n2032 = ( ~n1887 & n2030 ) | ( ~n1887 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = ( n1887 & n2030 ) | ( n1887 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2034 = ( n1887 & n2032 ) | ( n1887 & ~n2033 ) | ( n2032 & ~n2033 ) ;
  assign n2035 = ( x77 & n2029 ) | ( x77 & ~n2034 ) | ( n2029 & ~n2034 ) ;
  assign n2036 = ( x77 & n1888 ) | ( x77 & ~n1953 ) | ( n1888 & ~n1953 ) ;
  assign n2037 = x77 & n1888 ;
  assign n2038 = ( ~n1893 & n2036 ) | ( ~n1893 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2039 = ( n1893 & n2036 ) | ( n1893 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2040 = ( n1893 & n2038 ) | ( n1893 & ~n2039 ) | ( n2038 & ~n2039 ) ;
  assign n2041 = ( x78 & n2035 ) | ( x78 & ~n2040 ) | ( n2035 & ~n2040 ) ;
  assign n2042 = ( x78 & n1894 ) | ( x78 & ~n1953 ) | ( n1894 & ~n1953 ) ;
  assign n2043 = x78 & n1894 ;
  assign n2044 = ( ~n1899 & n2042 ) | ( ~n1899 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2045 = ( n1899 & n2042 ) | ( n1899 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2046 = ( n1899 & n2044 ) | ( n1899 & ~n2045 ) | ( n2044 & ~n2045 ) ;
  assign n2047 = ( x79 & n2041 ) | ( x79 & ~n2046 ) | ( n2041 & ~n2046 ) ;
  assign n2048 = ( x79 & n1900 ) | ( x79 & ~n1953 ) | ( n1900 & ~n1953 ) ;
  assign n2049 = x79 & n1900 ;
  assign n2050 = ( ~n1905 & n2048 ) | ( ~n1905 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = ( n1905 & n2048 ) | ( n1905 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2052 = ( n1905 & n2050 ) | ( n1905 & ~n2051 ) | ( n2050 & ~n2051 ) ;
  assign n2053 = ( x80 & n2047 ) | ( x80 & ~n2052 ) | ( n2047 & ~n2052 ) ;
  assign n2054 = ( x80 & n1906 ) | ( x80 & ~n1953 ) | ( n1906 & ~n1953 ) ;
  assign n2055 = x80 & n1906 ;
  assign n2056 = ( ~n1911 & n2054 ) | ( ~n1911 & n2055 ) | ( n2054 & n2055 ) ;
  assign n2057 = ( n1911 & n2054 ) | ( n1911 & n2055 ) | ( n2054 & n2055 ) ;
  assign n2058 = ( n1911 & n2056 ) | ( n1911 & ~n2057 ) | ( n2056 & ~n2057 ) ;
  assign n2059 = ( x81 & n2053 ) | ( x81 & ~n2058 ) | ( n2053 & ~n2058 ) ;
  assign n2060 = ( x81 & n1912 ) | ( x81 & ~n1953 ) | ( n1912 & ~n1953 ) ;
  assign n2061 = x81 & n1912 ;
  assign n2062 = ( ~n1917 & n2060 ) | ( ~n1917 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2063 = ( n1917 & n2060 ) | ( n1917 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2064 = ( n1917 & n2062 ) | ( n1917 & ~n2063 ) | ( n2062 & ~n2063 ) ;
  assign n2065 = ( x82 & n2059 ) | ( x82 & ~n2064 ) | ( n2059 & ~n2064 ) ;
  assign n2066 = ( x82 & n1918 ) | ( x82 & ~n1953 ) | ( n1918 & ~n1953 ) ;
  assign n2067 = x82 & n1918 ;
  assign n2068 = ( ~n1923 & n2066 ) | ( ~n1923 & n2067 ) | ( n2066 & n2067 ) ;
  assign n2069 = ( n1923 & n2066 ) | ( n1923 & n2067 ) | ( n2066 & n2067 ) ;
  assign n2070 = ( n1923 & n2068 ) | ( n1923 & ~n2069 ) | ( n2068 & ~n2069 ) ;
  assign n2071 = ( x83 & n2065 ) | ( x83 & ~n2070 ) | ( n2065 & ~n2070 ) ;
  assign n2072 = ( x83 & n1924 ) | ( x83 & ~n1953 ) | ( n1924 & ~n1953 ) ;
  assign n2073 = x83 & n1924 ;
  assign n2074 = ( ~n1929 & n2072 ) | ( ~n1929 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2075 = ( n1929 & n2072 ) | ( n1929 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2076 = ( n1929 & n2074 ) | ( n1929 & ~n2075 ) | ( n2074 & ~n2075 ) ;
  assign n2077 = ( x84 & n2071 ) | ( x84 & ~n2076 ) | ( n2071 & ~n2076 ) ;
  assign n2078 = ( x84 & n1930 ) | ( x84 & ~n1953 ) | ( n1930 & ~n1953 ) ;
  assign n2079 = x84 & n1930 ;
  assign n2080 = ( ~n1935 & n2078 ) | ( ~n1935 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2081 = ( n1935 & n2078 ) | ( n1935 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2082 = ( n1935 & n2080 ) | ( n1935 & ~n2081 ) | ( n2080 & ~n2081 ) ;
  assign n2083 = ( x85 & n2077 ) | ( x85 & ~n2082 ) | ( n2077 & ~n2082 ) ;
  assign n2084 = ( x85 & n1936 ) | ( x85 & ~n1953 ) | ( n1936 & ~n1953 ) ;
  assign n2085 = x85 & n1936 ;
  assign n2086 = ( ~n1941 & n2084 ) | ( ~n1941 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2087 = ( n1941 & n2084 ) | ( n1941 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2088 = ( n1941 & n2086 ) | ( n1941 & ~n2087 ) | ( n2086 & ~n2087 ) ;
  assign n2089 = ( x86 & n2083 ) | ( x86 & ~n2088 ) | ( n2083 & ~n2088 ) ;
  assign n2090 = ( x86 & n1942 ) | ( x86 & ~n1953 ) | ( n1942 & ~n1953 ) ;
  assign n2091 = x86 & n1942 ;
  assign n2092 = ( ~n1947 & n2090 ) | ( ~n1947 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = ( n1947 & n2090 ) | ( n1947 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2094 = ( n1947 & n2092 ) | ( n1947 & ~n2093 ) | ( n2092 & ~n2093 ) ;
  assign n2095 = ( x87 & n2089 ) | ( x87 & ~n2094 ) | ( n2089 & ~n2094 ) ;
  assign n2096 = ( x88 & n168 ) | ( x88 & n1949 ) | ( n168 & n1949 ) ;
  assign n2097 = x88 | n1949 ;
  assign n2098 = ( n1951 & n2096 ) | ( n1951 & ~n2097 ) | ( n2096 & ~n2097 ) ;
  assign n2099 = ( x88 & ~n1958 ) | ( x88 & n2095 ) | ( ~n1958 & n2095 ) ;
  assign n2100 = ( x89 & ~n2098 ) | ( x89 & n2099 ) | ( ~n2098 & n2099 ) ;
  assign n2101 = n167 | n2100 ;
  assign n2102 = ( x88 & n2095 ) | ( x88 & n2101 ) | ( n2095 & n2101 ) ;
  assign n2103 = x88 | n2095 ;
  assign n2104 = ( ~n1958 & n2102 ) | ( ~n1958 & n2103 ) | ( n2102 & n2103 ) ;
  assign n2105 = ( n1958 & n2102 ) | ( n1958 & n2103 ) | ( n2102 & n2103 ) ;
  assign n2106 = ( n1958 & n2104 ) | ( n1958 & ~n2105 ) | ( n2104 & ~n2105 ) ;
  assign n2107 = ~x37 & x64 ;
  assign n2108 = ~x38 & n2101 ;
  assign n2109 = ( x38 & ~x64 ) | ( x38 & n2101 ) | ( ~x64 & n2101 ) ;
  assign n2110 = ( n1959 & ~n2108 ) | ( n1959 & n2109 ) | ( ~n2108 & n2109 ) ;
  assign n2111 = ( x65 & n2107 ) | ( x65 & ~n2110 ) | ( n2107 & ~n2110 ) ;
  assign n2112 = ( x65 & n1959 ) | ( x65 & n2101 ) | ( n1959 & n2101 ) ;
  assign n2113 = x65 | n1959 ;
  assign n2114 = ( ~n1962 & n2112 ) | ( ~n1962 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2115 = ( n1962 & n2112 ) | ( n1962 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2116 = ( n1962 & n2114 ) | ( n1962 & ~n2115 ) | ( n2114 & ~n2115 ) ;
  assign n2117 = ( x66 & n2111 ) | ( x66 & ~n2116 ) | ( n2111 & ~n2116 ) ;
  assign n2118 = ( x66 & n1963 ) | ( x66 & n2101 ) | ( n1963 & n2101 ) ;
  assign n2119 = x66 | n1963 ;
  assign n2120 = ( ~n1968 & n2118 ) | ( ~n1968 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2121 = ( n1968 & n2118 ) | ( n1968 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2122 = ( n1968 & n2120 ) | ( n1968 & ~n2121 ) | ( n2120 & ~n2121 ) ;
  assign n2123 = ( x67 & n2117 ) | ( x67 & ~n2122 ) | ( n2117 & ~n2122 ) ;
  assign n2124 = ( x67 & n1969 ) | ( x67 & ~n2101 ) | ( n1969 & ~n2101 ) ;
  assign n2125 = x67 & n1969 ;
  assign n2126 = ( ~n1974 & n2124 ) | ( ~n1974 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( n1974 & n2124 ) | ( n1974 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2128 = ( n1974 & n2126 ) | ( n1974 & ~n2127 ) | ( n2126 & ~n2127 ) ;
  assign n2129 = ( x68 & n2123 ) | ( x68 & ~n2128 ) | ( n2123 & ~n2128 ) ;
  assign n2130 = ( x68 & n1975 ) | ( x68 & ~n2101 ) | ( n1975 & ~n2101 ) ;
  assign n2131 = x68 & n1975 ;
  assign n2132 = ( ~n1980 & n2130 ) | ( ~n1980 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2133 = ( n1980 & n2130 ) | ( n1980 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2134 = ( n1980 & n2132 ) | ( n1980 & ~n2133 ) | ( n2132 & ~n2133 ) ;
  assign n2135 = ( x69 & n2129 ) | ( x69 & ~n2134 ) | ( n2129 & ~n2134 ) ;
  assign n2136 = ( x69 & n1981 ) | ( x69 & ~n2101 ) | ( n1981 & ~n2101 ) ;
  assign n2137 = x69 & n1981 ;
  assign n2138 = ( ~n1986 & n2136 ) | ( ~n1986 & n2137 ) | ( n2136 & n2137 ) ;
  assign n2139 = ( n1986 & n2136 ) | ( n1986 & n2137 ) | ( n2136 & n2137 ) ;
  assign n2140 = ( n1986 & n2138 ) | ( n1986 & ~n2139 ) | ( n2138 & ~n2139 ) ;
  assign n2141 = ( x70 & n2135 ) | ( x70 & ~n2140 ) | ( n2135 & ~n2140 ) ;
  assign n2142 = ( x70 & n1987 ) | ( x70 & ~n2101 ) | ( n1987 & ~n2101 ) ;
  assign n2143 = x70 & n1987 ;
  assign n2144 = ( ~n1992 & n2142 ) | ( ~n1992 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2145 = ( n1992 & n2142 ) | ( n1992 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2146 = ( n1992 & n2144 ) | ( n1992 & ~n2145 ) | ( n2144 & ~n2145 ) ;
  assign n2147 = ( x71 & n2141 ) | ( x71 & ~n2146 ) | ( n2141 & ~n2146 ) ;
  assign n2148 = ( x71 & n1993 ) | ( x71 & ~n2101 ) | ( n1993 & ~n2101 ) ;
  assign n2149 = x71 & n1993 ;
  assign n2150 = ( ~n1998 & n2148 ) | ( ~n1998 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = ( n1998 & n2148 ) | ( n1998 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2152 = ( n1998 & n2150 ) | ( n1998 & ~n2151 ) | ( n2150 & ~n2151 ) ;
  assign n2153 = ( x72 & n2147 ) | ( x72 & ~n2152 ) | ( n2147 & ~n2152 ) ;
  assign n2154 = ( x72 & n1999 ) | ( x72 & ~n2101 ) | ( n1999 & ~n2101 ) ;
  assign n2155 = x72 & n1999 ;
  assign n2156 = ( ~n2004 & n2154 ) | ( ~n2004 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ( n2004 & n2154 ) | ( n2004 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2158 = ( n2004 & n2156 ) | ( n2004 & ~n2157 ) | ( n2156 & ~n2157 ) ;
  assign n2159 = ( x73 & n2153 ) | ( x73 & ~n2158 ) | ( n2153 & ~n2158 ) ;
  assign n2160 = ( x73 & n2005 ) | ( x73 & ~n2101 ) | ( n2005 & ~n2101 ) ;
  assign n2161 = x73 & n2005 ;
  assign n2162 = ( ~n2010 & n2160 ) | ( ~n2010 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = ( n2010 & n2160 ) | ( n2010 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2164 = ( n2010 & n2162 ) | ( n2010 & ~n2163 ) | ( n2162 & ~n2163 ) ;
  assign n2165 = ( x74 & n2159 ) | ( x74 & ~n2164 ) | ( n2159 & ~n2164 ) ;
  assign n2166 = ( x74 & n2011 ) | ( x74 & ~n2101 ) | ( n2011 & ~n2101 ) ;
  assign n2167 = x74 & n2011 ;
  assign n2168 = ( ~n2016 & n2166 ) | ( ~n2016 & n2167 ) | ( n2166 & n2167 ) ;
  assign n2169 = ( n2016 & n2166 ) | ( n2016 & n2167 ) | ( n2166 & n2167 ) ;
  assign n2170 = ( n2016 & n2168 ) | ( n2016 & ~n2169 ) | ( n2168 & ~n2169 ) ;
  assign n2171 = ( x75 & n2165 ) | ( x75 & ~n2170 ) | ( n2165 & ~n2170 ) ;
  assign n2172 = ( x75 & n2017 ) | ( x75 & ~n2101 ) | ( n2017 & ~n2101 ) ;
  assign n2173 = x75 & n2017 ;
  assign n2174 = ( ~n2022 & n2172 ) | ( ~n2022 & n2173 ) | ( n2172 & n2173 ) ;
  assign n2175 = ( n2022 & n2172 ) | ( n2022 & n2173 ) | ( n2172 & n2173 ) ;
  assign n2176 = ( n2022 & n2174 ) | ( n2022 & ~n2175 ) | ( n2174 & ~n2175 ) ;
  assign n2177 = ( x76 & n2171 ) | ( x76 & ~n2176 ) | ( n2171 & ~n2176 ) ;
  assign n2178 = ( x76 & n2023 ) | ( x76 & ~n2101 ) | ( n2023 & ~n2101 ) ;
  assign n2179 = x76 & n2023 ;
  assign n2180 = ( ~n2028 & n2178 ) | ( ~n2028 & n2179 ) | ( n2178 & n2179 ) ;
  assign n2181 = ( n2028 & n2178 ) | ( n2028 & n2179 ) | ( n2178 & n2179 ) ;
  assign n2182 = ( n2028 & n2180 ) | ( n2028 & ~n2181 ) | ( n2180 & ~n2181 ) ;
  assign n2183 = ( x77 & n2177 ) | ( x77 & ~n2182 ) | ( n2177 & ~n2182 ) ;
  assign n2184 = ( x77 & n2029 ) | ( x77 & ~n2101 ) | ( n2029 & ~n2101 ) ;
  assign n2185 = x77 & n2029 ;
  assign n2186 = ( ~n2034 & n2184 ) | ( ~n2034 & n2185 ) | ( n2184 & n2185 ) ;
  assign n2187 = ( n2034 & n2184 ) | ( n2034 & n2185 ) | ( n2184 & n2185 ) ;
  assign n2188 = ( n2034 & n2186 ) | ( n2034 & ~n2187 ) | ( n2186 & ~n2187 ) ;
  assign n2189 = ( x78 & n2183 ) | ( x78 & ~n2188 ) | ( n2183 & ~n2188 ) ;
  assign n2190 = ( x78 & n2035 ) | ( x78 & ~n2101 ) | ( n2035 & ~n2101 ) ;
  assign n2191 = x78 & n2035 ;
  assign n2192 = ( ~n2040 & n2190 ) | ( ~n2040 & n2191 ) | ( n2190 & n2191 ) ;
  assign n2193 = ( n2040 & n2190 ) | ( n2040 & n2191 ) | ( n2190 & n2191 ) ;
  assign n2194 = ( n2040 & n2192 ) | ( n2040 & ~n2193 ) | ( n2192 & ~n2193 ) ;
  assign n2195 = ( x79 & n2189 ) | ( x79 & ~n2194 ) | ( n2189 & ~n2194 ) ;
  assign n2196 = ( x79 & n2041 ) | ( x79 & ~n2101 ) | ( n2041 & ~n2101 ) ;
  assign n2197 = x79 & n2041 ;
  assign n2198 = ( ~n2046 & n2196 ) | ( ~n2046 & n2197 ) | ( n2196 & n2197 ) ;
  assign n2199 = ( n2046 & n2196 ) | ( n2046 & n2197 ) | ( n2196 & n2197 ) ;
  assign n2200 = ( n2046 & n2198 ) | ( n2046 & ~n2199 ) | ( n2198 & ~n2199 ) ;
  assign n2201 = ( x80 & n2195 ) | ( x80 & ~n2200 ) | ( n2195 & ~n2200 ) ;
  assign n2202 = ( x80 & n2047 ) | ( x80 & ~n2101 ) | ( n2047 & ~n2101 ) ;
  assign n2203 = x80 & n2047 ;
  assign n2204 = ( ~n2052 & n2202 ) | ( ~n2052 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2205 = ( n2052 & n2202 ) | ( n2052 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2206 = ( n2052 & n2204 ) | ( n2052 & ~n2205 ) | ( n2204 & ~n2205 ) ;
  assign n2207 = ( x81 & n2201 ) | ( x81 & ~n2206 ) | ( n2201 & ~n2206 ) ;
  assign n2208 = ( x81 & n2053 ) | ( x81 & ~n2101 ) | ( n2053 & ~n2101 ) ;
  assign n2209 = x81 & n2053 ;
  assign n2210 = ( ~n2058 & n2208 ) | ( ~n2058 & n2209 ) | ( n2208 & n2209 ) ;
  assign n2211 = ( n2058 & n2208 ) | ( n2058 & n2209 ) | ( n2208 & n2209 ) ;
  assign n2212 = ( n2058 & n2210 ) | ( n2058 & ~n2211 ) | ( n2210 & ~n2211 ) ;
  assign n2213 = ( x82 & n2207 ) | ( x82 & ~n2212 ) | ( n2207 & ~n2212 ) ;
  assign n2214 = ( x82 & n2059 ) | ( x82 & ~n2101 ) | ( n2059 & ~n2101 ) ;
  assign n2215 = x82 & n2059 ;
  assign n2216 = ( ~n2064 & n2214 ) | ( ~n2064 & n2215 ) | ( n2214 & n2215 ) ;
  assign n2217 = ( n2064 & n2214 ) | ( n2064 & n2215 ) | ( n2214 & n2215 ) ;
  assign n2218 = ( n2064 & n2216 ) | ( n2064 & ~n2217 ) | ( n2216 & ~n2217 ) ;
  assign n2219 = ( x83 & n2213 ) | ( x83 & ~n2218 ) | ( n2213 & ~n2218 ) ;
  assign n2220 = ( x83 & n2065 ) | ( x83 & ~n2101 ) | ( n2065 & ~n2101 ) ;
  assign n2221 = x83 & n2065 ;
  assign n2222 = ( ~n2070 & n2220 ) | ( ~n2070 & n2221 ) | ( n2220 & n2221 ) ;
  assign n2223 = ( n2070 & n2220 ) | ( n2070 & n2221 ) | ( n2220 & n2221 ) ;
  assign n2224 = ( n2070 & n2222 ) | ( n2070 & ~n2223 ) | ( n2222 & ~n2223 ) ;
  assign n2225 = ( x84 & n2219 ) | ( x84 & ~n2224 ) | ( n2219 & ~n2224 ) ;
  assign n2226 = ( x84 & n2071 ) | ( x84 & ~n2101 ) | ( n2071 & ~n2101 ) ;
  assign n2227 = x84 & n2071 ;
  assign n2228 = ( ~n2076 & n2226 ) | ( ~n2076 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2229 = ( n2076 & n2226 ) | ( n2076 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2230 = ( n2076 & n2228 ) | ( n2076 & ~n2229 ) | ( n2228 & ~n2229 ) ;
  assign n2231 = ( x85 & n2225 ) | ( x85 & ~n2230 ) | ( n2225 & ~n2230 ) ;
  assign n2232 = ( x85 & n2077 ) | ( x85 & ~n2101 ) | ( n2077 & ~n2101 ) ;
  assign n2233 = x85 & n2077 ;
  assign n2234 = ( ~n2082 & n2232 ) | ( ~n2082 & n2233 ) | ( n2232 & n2233 ) ;
  assign n2235 = ( n2082 & n2232 ) | ( n2082 & n2233 ) | ( n2232 & n2233 ) ;
  assign n2236 = ( n2082 & n2234 ) | ( n2082 & ~n2235 ) | ( n2234 & ~n2235 ) ;
  assign n2237 = ( x86 & n2231 ) | ( x86 & ~n2236 ) | ( n2231 & ~n2236 ) ;
  assign n2238 = ( x86 & n2083 ) | ( x86 & ~n2101 ) | ( n2083 & ~n2101 ) ;
  assign n2239 = x86 & n2083 ;
  assign n2240 = ( ~n2088 & n2238 ) | ( ~n2088 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2241 = ( n2088 & n2238 ) | ( n2088 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2242 = ( n2088 & n2240 ) | ( n2088 & ~n2241 ) | ( n2240 & ~n2241 ) ;
  assign n2243 = ( x87 & n2237 ) | ( x87 & ~n2242 ) | ( n2237 & ~n2242 ) ;
  assign n2244 = ( x87 & n2089 ) | ( x87 & ~n2101 ) | ( n2089 & ~n2101 ) ;
  assign n2245 = x87 & n2089 ;
  assign n2246 = ( ~n2094 & n2244 ) | ( ~n2094 & n2245 ) | ( n2244 & n2245 ) ;
  assign n2247 = ( n2094 & n2244 ) | ( n2094 & n2245 ) | ( n2244 & n2245 ) ;
  assign n2248 = ( n2094 & n2246 ) | ( n2094 & ~n2247 ) | ( n2246 & ~n2247 ) ;
  assign n2249 = ( x88 & n2243 ) | ( x88 & ~n2248 ) | ( n2243 & ~n2248 ) ;
  assign n2250 = ( x89 & ~n2106 ) | ( x89 & n2249 ) | ( ~n2106 & n2249 ) ;
  assign n2251 = ~n166 & n2098 ;
  assign n2252 = n167 & ~n2251 ;
  assign n2253 = ( x89 & x90 ) | ( x89 & ~n2099 ) | ( x90 & ~n2099 ) ;
  assign n2254 = ( ~x89 & x90 ) | ( ~x89 & n2099 ) | ( x90 & n2099 ) ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = n2251 & ~n2255 ;
  assign n2257 = ( n2250 & n2252 ) | ( n2250 & ~n2256 ) | ( n2252 & ~n2256 ) ;
  assign n2258 = ( x89 & n2249 ) | ( x89 & n2257 ) | ( n2249 & n2257 ) ;
  assign n2259 = x89 | n2249 ;
  assign n2260 = ( ~n2106 & n2258 ) | ( ~n2106 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2261 = ( n2106 & n2258 ) | ( n2106 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2262 = ( n2106 & n2260 ) | ( n2106 & ~n2261 ) | ( n2260 & ~n2261 ) ;
  assign n2263 = ~x36 & x64 ;
  assign n2264 = ~x37 & n2257 ;
  assign n2265 = ( x37 & ~x64 ) | ( x37 & n2257 ) | ( ~x64 & n2257 ) ;
  assign n2266 = ( n2107 & ~n2264 ) | ( n2107 & n2265 ) | ( ~n2264 & n2265 ) ;
  assign n2267 = ( x65 & n2263 ) | ( x65 & ~n2266 ) | ( n2263 & ~n2266 ) ;
  assign n2268 = ( x65 & n2107 ) | ( x65 & n2257 ) | ( n2107 & n2257 ) ;
  assign n2269 = x65 | n2107 ;
  assign n2270 = ( ~n2110 & n2268 ) | ( ~n2110 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2271 = ( n2110 & n2268 ) | ( n2110 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2272 = ( n2110 & n2270 ) | ( n2110 & ~n2271 ) | ( n2270 & ~n2271 ) ;
  assign n2273 = ( x66 & n2267 ) | ( x66 & ~n2272 ) | ( n2267 & ~n2272 ) ;
  assign n2274 = ( x66 & n2111 ) | ( x66 & n2257 ) | ( n2111 & n2257 ) ;
  assign n2275 = x66 | n2111 ;
  assign n2276 = ( ~n2116 & n2274 ) | ( ~n2116 & n2275 ) | ( n2274 & n2275 ) ;
  assign n2277 = ( n2116 & n2274 ) | ( n2116 & n2275 ) | ( n2274 & n2275 ) ;
  assign n2278 = ( n2116 & n2276 ) | ( n2116 & ~n2277 ) | ( n2276 & ~n2277 ) ;
  assign n2279 = ( x67 & n2273 ) | ( x67 & ~n2278 ) | ( n2273 & ~n2278 ) ;
  assign n2280 = ( x67 & n2117 ) | ( x67 & ~n2257 ) | ( n2117 & ~n2257 ) ;
  assign n2281 = x67 & n2117 ;
  assign n2282 = ( ~n2122 & n2280 ) | ( ~n2122 & n2281 ) | ( n2280 & n2281 ) ;
  assign n2283 = ( n2122 & n2280 ) | ( n2122 & n2281 ) | ( n2280 & n2281 ) ;
  assign n2284 = ( n2122 & n2282 ) | ( n2122 & ~n2283 ) | ( n2282 & ~n2283 ) ;
  assign n2285 = ( x68 & n2279 ) | ( x68 & ~n2284 ) | ( n2279 & ~n2284 ) ;
  assign n2286 = ( x68 & n2123 ) | ( x68 & ~n2257 ) | ( n2123 & ~n2257 ) ;
  assign n2287 = x68 & n2123 ;
  assign n2288 = ( ~n2128 & n2286 ) | ( ~n2128 & n2287 ) | ( n2286 & n2287 ) ;
  assign n2289 = ( n2128 & n2286 ) | ( n2128 & n2287 ) | ( n2286 & n2287 ) ;
  assign n2290 = ( n2128 & n2288 ) | ( n2128 & ~n2289 ) | ( n2288 & ~n2289 ) ;
  assign n2291 = ( x69 & n2285 ) | ( x69 & ~n2290 ) | ( n2285 & ~n2290 ) ;
  assign n2292 = ( x69 & n2129 ) | ( x69 & ~n2257 ) | ( n2129 & ~n2257 ) ;
  assign n2293 = x69 & n2129 ;
  assign n2294 = ( ~n2134 & n2292 ) | ( ~n2134 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2295 = ( n2134 & n2292 ) | ( n2134 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2296 = ( n2134 & n2294 ) | ( n2134 & ~n2295 ) | ( n2294 & ~n2295 ) ;
  assign n2297 = ( x70 & n2291 ) | ( x70 & ~n2296 ) | ( n2291 & ~n2296 ) ;
  assign n2298 = ( x70 & n2135 ) | ( x70 & ~n2257 ) | ( n2135 & ~n2257 ) ;
  assign n2299 = x70 & n2135 ;
  assign n2300 = ( ~n2140 & n2298 ) | ( ~n2140 & n2299 ) | ( n2298 & n2299 ) ;
  assign n2301 = ( n2140 & n2298 ) | ( n2140 & n2299 ) | ( n2298 & n2299 ) ;
  assign n2302 = ( n2140 & n2300 ) | ( n2140 & ~n2301 ) | ( n2300 & ~n2301 ) ;
  assign n2303 = ( x71 & n2297 ) | ( x71 & ~n2302 ) | ( n2297 & ~n2302 ) ;
  assign n2304 = ( x71 & n2141 ) | ( x71 & ~n2257 ) | ( n2141 & ~n2257 ) ;
  assign n2305 = x71 & n2141 ;
  assign n2306 = ( ~n2146 & n2304 ) | ( ~n2146 & n2305 ) | ( n2304 & n2305 ) ;
  assign n2307 = ( n2146 & n2304 ) | ( n2146 & n2305 ) | ( n2304 & n2305 ) ;
  assign n2308 = ( n2146 & n2306 ) | ( n2146 & ~n2307 ) | ( n2306 & ~n2307 ) ;
  assign n2309 = ( x72 & n2303 ) | ( x72 & ~n2308 ) | ( n2303 & ~n2308 ) ;
  assign n2310 = ( x72 & n2147 ) | ( x72 & ~n2257 ) | ( n2147 & ~n2257 ) ;
  assign n2311 = x72 & n2147 ;
  assign n2312 = ( ~n2152 & n2310 ) | ( ~n2152 & n2311 ) | ( n2310 & n2311 ) ;
  assign n2313 = ( n2152 & n2310 ) | ( n2152 & n2311 ) | ( n2310 & n2311 ) ;
  assign n2314 = ( n2152 & n2312 ) | ( n2152 & ~n2313 ) | ( n2312 & ~n2313 ) ;
  assign n2315 = ( x73 & n2309 ) | ( x73 & ~n2314 ) | ( n2309 & ~n2314 ) ;
  assign n2316 = ( x73 & n2153 ) | ( x73 & ~n2257 ) | ( n2153 & ~n2257 ) ;
  assign n2317 = x73 & n2153 ;
  assign n2318 = ( ~n2158 & n2316 ) | ( ~n2158 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2319 = ( n2158 & n2316 ) | ( n2158 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2320 = ( n2158 & n2318 ) | ( n2158 & ~n2319 ) | ( n2318 & ~n2319 ) ;
  assign n2321 = ( x74 & n2315 ) | ( x74 & ~n2320 ) | ( n2315 & ~n2320 ) ;
  assign n2322 = ( x74 & n2159 ) | ( x74 & ~n2257 ) | ( n2159 & ~n2257 ) ;
  assign n2323 = x74 & n2159 ;
  assign n2324 = ( ~n2164 & n2322 ) | ( ~n2164 & n2323 ) | ( n2322 & n2323 ) ;
  assign n2325 = ( n2164 & n2322 ) | ( n2164 & n2323 ) | ( n2322 & n2323 ) ;
  assign n2326 = ( n2164 & n2324 ) | ( n2164 & ~n2325 ) | ( n2324 & ~n2325 ) ;
  assign n2327 = ( x75 & n2321 ) | ( x75 & ~n2326 ) | ( n2321 & ~n2326 ) ;
  assign n2328 = ( x75 & n2165 ) | ( x75 & ~n2257 ) | ( n2165 & ~n2257 ) ;
  assign n2329 = x75 & n2165 ;
  assign n2330 = ( ~n2170 & n2328 ) | ( ~n2170 & n2329 ) | ( n2328 & n2329 ) ;
  assign n2331 = ( n2170 & n2328 ) | ( n2170 & n2329 ) | ( n2328 & n2329 ) ;
  assign n2332 = ( n2170 & n2330 ) | ( n2170 & ~n2331 ) | ( n2330 & ~n2331 ) ;
  assign n2333 = ( x76 & n2327 ) | ( x76 & ~n2332 ) | ( n2327 & ~n2332 ) ;
  assign n2334 = ( x76 & n2171 ) | ( x76 & ~n2257 ) | ( n2171 & ~n2257 ) ;
  assign n2335 = x76 & n2171 ;
  assign n2336 = ( ~n2176 & n2334 ) | ( ~n2176 & n2335 ) | ( n2334 & n2335 ) ;
  assign n2337 = ( n2176 & n2334 ) | ( n2176 & n2335 ) | ( n2334 & n2335 ) ;
  assign n2338 = ( n2176 & n2336 ) | ( n2176 & ~n2337 ) | ( n2336 & ~n2337 ) ;
  assign n2339 = ( x77 & n2333 ) | ( x77 & ~n2338 ) | ( n2333 & ~n2338 ) ;
  assign n2340 = ( x77 & n2177 ) | ( x77 & ~n2257 ) | ( n2177 & ~n2257 ) ;
  assign n2341 = x77 & n2177 ;
  assign n2342 = ( ~n2182 & n2340 ) | ( ~n2182 & n2341 ) | ( n2340 & n2341 ) ;
  assign n2343 = ( n2182 & n2340 ) | ( n2182 & n2341 ) | ( n2340 & n2341 ) ;
  assign n2344 = ( n2182 & n2342 ) | ( n2182 & ~n2343 ) | ( n2342 & ~n2343 ) ;
  assign n2345 = ( x78 & n2339 ) | ( x78 & ~n2344 ) | ( n2339 & ~n2344 ) ;
  assign n2346 = ( x78 & n2183 ) | ( x78 & ~n2257 ) | ( n2183 & ~n2257 ) ;
  assign n2347 = x78 & n2183 ;
  assign n2348 = ( ~n2188 & n2346 ) | ( ~n2188 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2349 = ( n2188 & n2346 ) | ( n2188 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2350 = ( n2188 & n2348 ) | ( n2188 & ~n2349 ) | ( n2348 & ~n2349 ) ;
  assign n2351 = ( x79 & n2345 ) | ( x79 & ~n2350 ) | ( n2345 & ~n2350 ) ;
  assign n2352 = ( x79 & n2189 ) | ( x79 & ~n2257 ) | ( n2189 & ~n2257 ) ;
  assign n2353 = x79 & n2189 ;
  assign n2354 = ( ~n2194 & n2352 ) | ( ~n2194 & n2353 ) | ( n2352 & n2353 ) ;
  assign n2355 = ( n2194 & n2352 ) | ( n2194 & n2353 ) | ( n2352 & n2353 ) ;
  assign n2356 = ( n2194 & n2354 ) | ( n2194 & ~n2355 ) | ( n2354 & ~n2355 ) ;
  assign n2357 = ( x80 & n2351 ) | ( x80 & ~n2356 ) | ( n2351 & ~n2356 ) ;
  assign n2358 = ( x80 & n2195 ) | ( x80 & ~n2257 ) | ( n2195 & ~n2257 ) ;
  assign n2359 = x80 & n2195 ;
  assign n2360 = ( ~n2200 & n2358 ) | ( ~n2200 & n2359 ) | ( n2358 & n2359 ) ;
  assign n2361 = ( n2200 & n2358 ) | ( n2200 & n2359 ) | ( n2358 & n2359 ) ;
  assign n2362 = ( n2200 & n2360 ) | ( n2200 & ~n2361 ) | ( n2360 & ~n2361 ) ;
  assign n2363 = ( x81 & n2357 ) | ( x81 & ~n2362 ) | ( n2357 & ~n2362 ) ;
  assign n2364 = ( x81 & n2201 ) | ( x81 & ~n2257 ) | ( n2201 & ~n2257 ) ;
  assign n2365 = x81 & n2201 ;
  assign n2366 = ( ~n2206 & n2364 ) | ( ~n2206 & n2365 ) | ( n2364 & n2365 ) ;
  assign n2367 = ( n2206 & n2364 ) | ( n2206 & n2365 ) | ( n2364 & n2365 ) ;
  assign n2368 = ( n2206 & n2366 ) | ( n2206 & ~n2367 ) | ( n2366 & ~n2367 ) ;
  assign n2369 = ( x82 & n2363 ) | ( x82 & ~n2368 ) | ( n2363 & ~n2368 ) ;
  assign n2370 = ( x82 & n2207 ) | ( x82 & ~n2257 ) | ( n2207 & ~n2257 ) ;
  assign n2371 = x82 & n2207 ;
  assign n2372 = ( ~n2212 & n2370 ) | ( ~n2212 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = ( n2212 & n2370 ) | ( n2212 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2374 = ( n2212 & n2372 ) | ( n2212 & ~n2373 ) | ( n2372 & ~n2373 ) ;
  assign n2375 = ( x83 & n2369 ) | ( x83 & ~n2374 ) | ( n2369 & ~n2374 ) ;
  assign n2376 = ( x83 & n2213 ) | ( x83 & ~n2257 ) | ( n2213 & ~n2257 ) ;
  assign n2377 = x83 & n2213 ;
  assign n2378 = ( ~n2218 & n2376 ) | ( ~n2218 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2379 = ( n2218 & n2376 ) | ( n2218 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2380 = ( n2218 & n2378 ) | ( n2218 & ~n2379 ) | ( n2378 & ~n2379 ) ;
  assign n2381 = ( x84 & n2375 ) | ( x84 & ~n2380 ) | ( n2375 & ~n2380 ) ;
  assign n2382 = ( x84 & n2219 ) | ( x84 & ~n2257 ) | ( n2219 & ~n2257 ) ;
  assign n2383 = x84 & n2219 ;
  assign n2384 = ( ~n2224 & n2382 ) | ( ~n2224 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2385 = ( n2224 & n2382 ) | ( n2224 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2386 = ( n2224 & n2384 ) | ( n2224 & ~n2385 ) | ( n2384 & ~n2385 ) ;
  assign n2387 = ( x85 & n2381 ) | ( x85 & ~n2386 ) | ( n2381 & ~n2386 ) ;
  assign n2388 = ( x85 & n2225 ) | ( x85 & ~n2257 ) | ( n2225 & ~n2257 ) ;
  assign n2389 = x85 & n2225 ;
  assign n2390 = ( ~n2230 & n2388 ) | ( ~n2230 & n2389 ) | ( n2388 & n2389 ) ;
  assign n2391 = ( n2230 & n2388 ) | ( n2230 & n2389 ) | ( n2388 & n2389 ) ;
  assign n2392 = ( n2230 & n2390 ) | ( n2230 & ~n2391 ) | ( n2390 & ~n2391 ) ;
  assign n2393 = ( x86 & n2387 ) | ( x86 & ~n2392 ) | ( n2387 & ~n2392 ) ;
  assign n2394 = ( x86 & n2231 ) | ( x86 & ~n2257 ) | ( n2231 & ~n2257 ) ;
  assign n2395 = x86 & n2231 ;
  assign n2396 = ( ~n2236 & n2394 ) | ( ~n2236 & n2395 ) | ( n2394 & n2395 ) ;
  assign n2397 = ( n2236 & n2394 ) | ( n2236 & n2395 ) | ( n2394 & n2395 ) ;
  assign n2398 = ( n2236 & n2396 ) | ( n2236 & ~n2397 ) | ( n2396 & ~n2397 ) ;
  assign n2399 = ( x87 & n2393 ) | ( x87 & ~n2398 ) | ( n2393 & ~n2398 ) ;
  assign n2400 = ( x87 & n2237 ) | ( x87 & ~n2257 ) | ( n2237 & ~n2257 ) ;
  assign n2401 = x87 & n2237 ;
  assign n2402 = ( ~n2242 & n2400 ) | ( ~n2242 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2403 = ( n2242 & n2400 ) | ( n2242 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2404 = ( n2242 & n2402 ) | ( n2242 & ~n2403 ) | ( n2402 & ~n2403 ) ;
  assign n2405 = ( x88 & n2399 ) | ( x88 & ~n2404 ) | ( n2399 & ~n2404 ) ;
  assign n2406 = ( x88 & n2243 ) | ( x88 & ~n2257 ) | ( n2243 & ~n2257 ) ;
  assign n2407 = x88 & n2243 ;
  assign n2408 = ( ~n2248 & n2406 ) | ( ~n2248 & n2407 ) | ( n2406 & n2407 ) ;
  assign n2409 = ( n2248 & n2406 ) | ( n2248 & n2407 ) | ( n2406 & n2407 ) ;
  assign n2410 = ( n2248 & n2408 ) | ( n2248 & ~n2409 ) | ( n2408 & ~n2409 ) ;
  assign n2411 = ( x89 & n2405 ) | ( x89 & ~n2410 ) | ( n2405 & ~n2410 ) ;
  assign n2412 = ( x90 & ~n2262 ) | ( x90 & n2411 ) | ( ~n2262 & n2411 ) ;
  assign n2413 = n167 & n2250 ;
  assign n2414 = ~n166 & n2255 ;
  assign n2415 = n2250 | n2414 ;
  assign n2416 = ( n2098 & n2413 ) | ( n2098 & ~n2415 ) | ( n2413 & ~n2415 ) ;
  assign n2417 = ( x91 & n2412 ) | ( x91 & ~n2416 ) | ( n2412 & ~n2416 ) ;
  assign n2418 = n165 | n2417 ;
  assign n2419 = ( x90 & n2411 ) | ( x90 & n2418 ) | ( n2411 & n2418 ) ;
  assign n2420 = x90 | n2411 ;
  assign n2421 = ( ~n2262 & n2419 ) | ( ~n2262 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2422 = ( n2262 & n2419 ) | ( n2262 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2423 = ( n2262 & n2421 ) | ( n2262 & ~n2422 ) | ( n2421 & ~n2422 ) ;
  assign n2424 = ~x35 & x64 ;
  assign n2425 = ~x36 & n2418 ;
  assign n2426 = ( x36 & ~x64 ) | ( x36 & n2418 ) | ( ~x64 & n2418 ) ;
  assign n2427 = ( n2263 & ~n2425 ) | ( n2263 & n2426 ) | ( ~n2425 & n2426 ) ;
  assign n2428 = ( x65 & n2424 ) | ( x65 & ~n2427 ) | ( n2424 & ~n2427 ) ;
  assign n2429 = ( x65 & n2263 ) | ( x65 & n2418 ) | ( n2263 & n2418 ) ;
  assign n2430 = x65 | n2263 ;
  assign n2431 = ( ~n2266 & n2429 ) | ( ~n2266 & n2430 ) | ( n2429 & n2430 ) ;
  assign n2432 = ( n2266 & n2429 ) | ( n2266 & n2430 ) | ( n2429 & n2430 ) ;
  assign n2433 = ( n2266 & n2431 ) | ( n2266 & ~n2432 ) | ( n2431 & ~n2432 ) ;
  assign n2434 = ( x66 & n2428 ) | ( x66 & ~n2433 ) | ( n2428 & ~n2433 ) ;
  assign n2435 = ( x66 & n2267 ) | ( x66 & n2418 ) | ( n2267 & n2418 ) ;
  assign n2436 = x66 | n2267 ;
  assign n2437 = ( ~n2272 & n2435 ) | ( ~n2272 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2438 = ( n2272 & n2435 ) | ( n2272 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2439 = ( n2272 & n2437 ) | ( n2272 & ~n2438 ) | ( n2437 & ~n2438 ) ;
  assign n2440 = ( x67 & n2434 ) | ( x67 & ~n2439 ) | ( n2434 & ~n2439 ) ;
  assign n2441 = ( x67 & n2273 ) | ( x67 & ~n2418 ) | ( n2273 & ~n2418 ) ;
  assign n2442 = x67 & n2273 ;
  assign n2443 = ( ~n2278 & n2441 ) | ( ~n2278 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2444 = ( n2278 & n2441 ) | ( n2278 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2445 = ( n2278 & n2443 ) | ( n2278 & ~n2444 ) | ( n2443 & ~n2444 ) ;
  assign n2446 = ( x68 & n2440 ) | ( x68 & ~n2445 ) | ( n2440 & ~n2445 ) ;
  assign n2447 = ( x68 & n2279 ) | ( x68 & ~n2418 ) | ( n2279 & ~n2418 ) ;
  assign n2448 = x68 & n2279 ;
  assign n2449 = ( ~n2284 & n2447 ) | ( ~n2284 & n2448 ) | ( n2447 & n2448 ) ;
  assign n2450 = ( n2284 & n2447 ) | ( n2284 & n2448 ) | ( n2447 & n2448 ) ;
  assign n2451 = ( n2284 & n2449 ) | ( n2284 & ~n2450 ) | ( n2449 & ~n2450 ) ;
  assign n2452 = ( x69 & n2446 ) | ( x69 & ~n2451 ) | ( n2446 & ~n2451 ) ;
  assign n2453 = ( x69 & n2285 ) | ( x69 & ~n2418 ) | ( n2285 & ~n2418 ) ;
  assign n2454 = x69 & n2285 ;
  assign n2455 = ( ~n2290 & n2453 ) | ( ~n2290 & n2454 ) | ( n2453 & n2454 ) ;
  assign n2456 = ( n2290 & n2453 ) | ( n2290 & n2454 ) | ( n2453 & n2454 ) ;
  assign n2457 = ( n2290 & n2455 ) | ( n2290 & ~n2456 ) | ( n2455 & ~n2456 ) ;
  assign n2458 = ( x70 & n2452 ) | ( x70 & ~n2457 ) | ( n2452 & ~n2457 ) ;
  assign n2459 = ( x70 & n2291 ) | ( x70 & ~n2418 ) | ( n2291 & ~n2418 ) ;
  assign n2460 = x70 & n2291 ;
  assign n2461 = ( ~n2296 & n2459 ) | ( ~n2296 & n2460 ) | ( n2459 & n2460 ) ;
  assign n2462 = ( n2296 & n2459 ) | ( n2296 & n2460 ) | ( n2459 & n2460 ) ;
  assign n2463 = ( n2296 & n2461 ) | ( n2296 & ~n2462 ) | ( n2461 & ~n2462 ) ;
  assign n2464 = ( x71 & n2458 ) | ( x71 & ~n2463 ) | ( n2458 & ~n2463 ) ;
  assign n2465 = ( x71 & n2297 ) | ( x71 & ~n2418 ) | ( n2297 & ~n2418 ) ;
  assign n2466 = x71 & n2297 ;
  assign n2467 = ( ~n2302 & n2465 ) | ( ~n2302 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = ( n2302 & n2465 ) | ( n2302 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2469 = ( n2302 & n2467 ) | ( n2302 & ~n2468 ) | ( n2467 & ~n2468 ) ;
  assign n2470 = ( x72 & n2464 ) | ( x72 & ~n2469 ) | ( n2464 & ~n2469 ) ;
  assign n2471 = ( x72 & n2303 ) | ( x72 & ~n2418 ) | ( n2303 & ~n2418 ) ;
  assign n2472 = x72 & n2303 ;
  assign n2473 = ( ~n2308 & n2471 ) | ( ~n2308 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2474 = ( n2308 & n2471 ) | ( n2308 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2475 = ( n2308 & n2473 ) | ( n2308 & ~n2474 ) | ( n2473 & ~n2474 ) ;
  assign n2476 = ( x73 & n2470 ) | ( x73 & ~n2475 ) | ( n2470 & ~n2475 ) ;
  assign n2477 = ( x73 & n2309 ) | ( x73 & ~n2418 ) | ( n2309 & ~n2418 ) ;
  assign n2478 = x73 & n2309 ;
  assign n2479 = ( ~n2314 & n2477 ) | ( ~n2314 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2480 = ( n2314 & n2477 ) | ( n2314 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2481 = ( n2314 & n2479 ) | ( n2314 & ~n2480 ) | ( n2479 & ~n2480 ) ;
  assign n2482 = ( x74 & n2476 ) | ( x74 & ~n2481 ) | ( n2476 & ~n2481 ) ;
  assign n2483 = ( x74 & n2315 ) | ( x74 & ~n2418 ) | ( n2315 & ~n2418 ) ;
  assign n2484 = x74 & n2315 ;
  assign n2485 = ( ~n2320 & n2483 ) | ( ~n2320 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2486 = ( n2320 & n2483 ) | ( n2320 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2487 = ( n2320 & n2485 ) | ( n2320 & ~n2486 ) | ( n2485 & ~n2486 ) ;
  assign n2488 = ( x75 & n2482 ) | ( x75 & ~n2487 ) | ( n2482 & ~n2487 ) ;
  assign n2489 = ( x75 & n2321 ) | ( x75 & ~n2418 ) | ( n2321 & ~n2418 ) ;
  assign n2490 = x75 & n2321 ;
  assign n2491 = ( ~n2326 & n2489 ) | ( ~n2326 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = ( n2326 & n2489 ) | ( n2326 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2493 = ( n2326 & n2491 ) | ( n2326 & ~n2492 ) | ( n2491 & ~n2492 ) ;
  assign n2494 = ( x76 & n2488 ) | ( x76 & ~n2493 ) | ( n2488 & ~n2493 ) ;
  assign n2495 = ( x76 & n2327 ) | ( x76 & ~n2418 ) | ( n2327 & ~n2418 ) ;
  assign n2496 = x76 & n2327 ;
  assign n2497 = ( ~n2332 & n2495 ) | ( ~n2332 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2498 = ( n2332 & n2495 ) | ( n2332 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2499 = ( n2332 & n2497 ) | ( n2332 & ~n2498 ) | ( n2497 & ~n2498 ) ;
  assign n2500 = ( x77 & n2494 ) | ( x77 & ~n2499 ) | ( n2494 & ~n2499 ) ;
  assign n2501 = ( x77 & n2333 ) | ( x77 & ~n2418 ) | ( n2333 & ~n2418 ) ;
  assign n2502 = x77 & n2333 ;
  assign n2503 = ( ~n2338 & n2501 ) | ( ~n2338 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2504 = ( n2338 & n2501 ) | ( n2338 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2505 = ( n2338 & n2503 ) | ( n2338 & ~n2504 ) | ( n2503 & ~n2504 ) ;
  assign n2506 = ( x78 & n2500 ) | ( x78 & ~n2505 ) | ( n2500 & ~n2505 ) ;
  assign n2507 = ( x78 & n2339 ) | ( x78 & ~n2418 ) | ( n2339 & ~n2418 ) ;
  assign n2508 = x78 & n2339 ;
  assign n2509 = ( ~n2344 & n2507 ) | ( ~n2344 & n2508 ) | ( n2507 & n2508 ) ;
  assign n2510 = ( n2344 & n2507 ) | ( n2344 & n2508 ) | ( n2507 & n2508 ) ;
  assign n2511 = ( n2344 & n2509 ) | ( n2344 & ~n2510 ) | ( n2509 & ~n2510 ) ;
  assign n2512 = ( x79 & n2506 ) | ( x79 & ~n2511 ) | ( n2506 & ~n2511 ) ;
  assign n2513 = ( x79 & n2345 ) | ( x79 & ~n2418 ) | ( n2345 & ~n2418 ) ;
  assign n2514 = x79 & n2345 ;
  assign n2515 = ( ~n2350 & n2513 ) | ( ~n2350 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2516 = ( n2350 & n2513 ) | ( n2350 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2517 = ( n2350 & n2515 ) | ( n2350 & ~n2516 ) | ( n2515 & ~n2516 ) ;
  assign n2518 = ( x80 & n2512 ) | ( x80 & ~n2517 ) | ( n2512 & ~n2517 ) ;
  assign n2519 = ( x80 & n2351 ) | ( x80 & ~n2418 ) | ( n2351 & ~n2418 ) ;
  assign n2520 = x80 & n2351 ;
  assign n2521 = ( ~n2356 & n2519 ) | ( ~n2356 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2522 = ( n2356 & n2519 ) | ( n2356 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2523 = ( n2356 & n2521 ) | ( n2356 & ~n2522 ) | ( n2521 & ~n2522 ) ;
  assign n2524 = ( x81 & n2518 ) | ( x81 & ~n2523 ) | ( n2518 & ~n2523 ) ;
  assign n2525 = ( x81 & n2357 ) | ( x81 & ~n2418 ) | ( n2357 & ~n2418 ) ;
  assign n2526 = x81 & n2357 ;
  assign n2527 = ( ~n2362 & n2525 ) | ( ~n2362 & n2526 ) | ( n2525 & n2526 ) ;
  assign n2528 = ( n2362 & n2525 ) | ( n2362 & n2526 ) | ( n2525 & n2526 ) ;
  assign n2529 = ( n2362 & n2527 ) | ( n2362 & ~n2528 ) | ( n2527 & ~n2528 ) ;
  assign n2530 = ( x82 & n2524 ) | ( x82 & ~n2529 ) | ( n2524 & ~n2529 ) ;
  assign n2531 = ( x82 & n2363 ) | ( x82 & ~n2418 ) | ( n2363 & ~n2418 ) ;
  assign n2532 = x82 & n2363 ;
  assign n2533 = ( ~n2368 & n2531 ) | ( ~n2368 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2534 = ( n2368 & n2531 ) | ( n2368 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2535 = ( n2368 & n2533 ) | ( n2368 & ~n2534 ) | ( n2533 & ~n2534 ) ;
  assign n2536 = ( x83 & n2530 ) | ( x83 & ~n2535 ) | ( n2530 & ~n2535 ) ;
  assign n2537 = ( x83 & n2369 ) | ( x83 & ~n2418 ) | ( n2369 & ~n2418 ) ;
  assign n2538 = x83 & n2369 ;
  assign n2539 = ( ~n2374 & n2537 ) | ( ~n2374 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2540 = ( n2374 & n2537 ) | ( n2374 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2541 = ( n2374 & n2539 ) | ( n2374 & ~n2540 ) | ( n2539 & ~n2540 ) ;
  assign n2542 = ( x84 & n2536 ) | ( x84 & ~n2541 ) | ( n2536 & ~n2541 ) ;
  assign n2543 = ( x84 & n2375 ) | ( x84 & ~n2418 ) | ( n2375 & ~n2418 ) ;
  assign n2544 = x84 & n2375 ;
  assign n2545 = ( ~n2380 & n2543 ) | ( ~n2380 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2546 = ( n2380 & n2543 ) | ( n2380 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2547 = ( n2380 & n2545 ) | ( n2380 & ~n2546 ) | ( n2545 & ~n2546 ) ;
  assign n2548 = ( x85 & n2542 ) | ( x85 & ~n2547 ) | ( n2542 & ~n2547 ) ;
  assign n2549 = ( x85 & n2381 ) | ( x85 & ~n2418 ) | ( n2381 & ~n2418 ) ;
  assign n2550 = x85 & n2381 ;
  assign n2551 = ( ~n2386 & n2549 ) | ( ~n2386 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2552 = ( n2386 & n2549 ) | ( n2386 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2553 = ( n2386 & n2551 ) | ( n2386 & ~n2552 ) | ( n2551 & ~n2552 ) ;
  assign n2554 = ( x86 & n2548 ) | ( x86 & ~n2553 ) | ( n2548 & ~n2553 ) ;
  assign n2555 = ( x86 & n2387 ) | ( x86 & ~n2418 ) | ( n2387 & ~n2418 ) ;
  assign n2556 = x86 & n2387 ;
  assign n2557 = ( ~n2392 & n2555 ) | ( ~n2392 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2558 = ( n2392 & n2555 ) | ( n2392 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2559 = ( n2392 & n2557 ) | ( n2392 & ~n2558 ) | ( n2557 & ~n2558 ) ;
  assign n2560 = ( x87 & n2554 ) | ( x87 & ~n2559 ) | ( n2554 & ~n2559 ) ;
  assign n2561 = ( x87 & n2393 ) | ( x87 & ~n2418 ) | ( n2393 & ~n2418 ) ;
  assign n2562 = x87 & n2393 ;
  assign n2563 = ( ~n2398 & n2561 ) | ( ~n2398 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2564 = ( n2398 & n2561 ) | ( n2398 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2565 = ( n2398 & n2563 ) | ( n2398 & ~n2564 ) | ( n2563 & ~n2564 ) ;
  assign n2566 = ( x88 & n2560 ) | ( x88 & ~n2565 ) | ( n2560 & ~n2565 ) ;
  assign n2567 = ( x88 & n2399 ) | ( x88 & ~n2418 ) | ( n2399 & ~n2418 ) ;
  assign n2568 = x88 & n2399 ;
  assign n2569 = ( ~n2404 & n2567 ) | ( ~n2404 & n2568 ) | ( n2567 & n2568 ) ;
  assign n2570 = ( n2404 & n2567 ) | ( n2404 & n2568 ) | ( n2567 & n2568 ) ;
  assign n2571 = ( n2404 & n2569 ) | ( n2404 & ~n2570 ) | ( n2569 & ~n2570 ) ;
  assign n2572 = ( x89 & n2566 ) | ( x89 & ~n2571 ) | ( n2566 & ~n2571 ) ;
  assign n2573 = ( x89 & n2405 ) | ( x89 & ~n2418 ) | ( n2405 & ~n2418 ) ;
  assign n2574 = x89 & n2405 ;
  assign n2575 = ( ~n2410 & n2573 ) | ( ~n2410 & n2574 ) | ( n2573 & n2574 ) ;
  assign n2576 = ( n2410 & n2573 ) | ( n2410 & n2574 ) | ( n2573 & n2574 ) ;
  assign n2577 = ( n2410 & n2575 ) | ( n2410 & ~n2576 ) | ( n2575 & ~n2576 ) ;
  assign n2578 = ( x90 & n2572 ) | ( x90 & ~n2577 ) | ( n2572 & ~n2577 ) ;
  assign n2579 = ( x91 & ~n165 ) | ( x91 & n2412 ) | ( ~n165 & n2412 ) ;
  assign n2580 = x91 & n2412 ;
  assign n2581 = ( n2416 & ~n2579 ) | ( n2416 & n2580 ) | ( ~n2579 & n2580 ) ;
  assign n2582 = ( x91 & ~n2423 ) | ( x91 & n2578 ) | ( ~n2423 & n2578 ) ;
  assign n2583 = ( x92 & ~n2581 ) | ( x92 & n2582 ) | ( ~n2581 & n2582 ) ;
  assign n2584 = n164 | n2583 ;
  assign n2585 = ( x91 & n2578 ) | ( x91 & n2584 ) | ( n2578 & n2584 ) ;
  assign n2586 = x91 | n2578 ;
  assign n2587 = ( ~n2423 & n2585 ) | ( ~n2423 & n2586 ) | ( n2585 & n2586 ) ;
  assign n2588 = ( n2423 & n2585 ) | ( n2423 & n2586 ) | ( n2585 & n2586 ) ;
  assign n2589 = ( n2423 & n2587 ) | ( n2423 & ~n2588 ) | ( n2587 & ~n2588 ) ;
  assign n2590 = ~x34 & x64 ;
  assign n2591 = ~x35 & n2584 ;
  assign n2592 = ( x35 & ~x64 ) | ( x35 & n2584 ) | ( ~x64 & n2584 ) ;
  assign n2593 = ( n2424 & ~n2591 ) | ( n2424 & n2592 ) | ( ~n2591 & n2592 ) ;
  assign n2594 = ( x65 & n2590 ) | ( x65 & ~n2593 ) | ( n2590 & ~n2593 ) ;
  assign n2595 = ( x65 & n2424 ) | ( x65 & n2584 ) | ( n2424 & n2584 ) ;
  assign n2596 = x65 | n2424 ;
  assign n2597 = ( ~n2427 & n2595 ) | ( ~n2427 & n2596 ) | ( n2595 & n2596 ) ;
  assign n2598 = ( n2427 & n2595 ) | ( n2427 & n2596 ) | ( n2595 & n2596 ) ;
  assign n2599 = ( n2427 & n2597 ) | ( n2427 & ~n2598 ) | ( n2597 & ~n2598 ) ;
  assign n2600 = ( x66 & n2594 ) | ( x66 & ~n2599 ) | ( n2594 & ~n2599 ) ;
  assign n2601 = ( x66 & n2428 ) | ( x66 & n2584 ) | ( n2428 & n2584 ) ;
  assign n2602 = x66 | n2428 ;
  assign n2603 = ( ~n2433 & n2601 ) | ( ~n2433 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = ( n2433 & n2601 ) | ( n2433 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2605 = ( n2433 & n2603 ) | ( n2433 & ~n2604 ) | ( n2603 & ~n2604 ) ;
  assign n2606 = ( x67 & n2600 ) | ( x67 & ~n2605 ) | ( n2600 & ~n2605 ) ;
  assign n2607 = ( x67 & n2434 ) | ( x67 & ~n2584 ) | ( n2434 & ~n2584 ) ;
  assign n2608 = x67 & n2434 ;
  assign n2609 = ( ~n2439 & n2607 ) | ( ~n2439 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2610 = ( n2439 & n2607 ) | ( n2439 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2611 = ( n2439 & n2609 ) | ( n2439 & ~n2610 ) | ( n2609 & ~n2610 ) ;
  assign n2612 = ( x68 & n2606 ) | ( x68 & ~n2611 ) | ( n2606 & ~n2611 ) ;
  assign n2613 = ( x68 & n2440 ) | ( x68 & ~n2584 ) | ( n2440 & ~n2584 ) ;
  assign n2614 = x68 & n2440 ;
  assign n2615 = ( ~n2445 & n2613 ) | ( ~n2445 & n2614 ) | ( n2613 & n2614 ) ;
  assign n2616 = ( n2445 & n2613 ) | ( n2445 & n2614 ) | ( n2613 & n2614 ) ;
  assign n2617 = ( n2445 & n2615 ) | ( n2445 & ~n2616 ) | ( n2615 & ~n2616 ) ;
  assign n2618 = ( x69 & n2612 ) | ( x69 & ~n2617 ) | ( n2612 & ~n2617 ) ;
  assign n2619 = ( x69 & n2446 ) | ( x69 & ~n2584 ) | ( n2446 & ~n2584 ) ;
  assign n2620 = x69 & n2446 ;
  assign n2621 = ( ~n2451 & n2619 ) | ( ~n2451 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2622 = ( n2451 & n2619 ) | ( n2451 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2623 = ( n2451 & n2621 ) | ( n2451 & ~n2622 ) | ( n2621 & ~n2622 ) ;
  assign n2624 = ( x70 & n2618 ) | ( x70 & ~n2623 ) | ( n2618 & ~n2623 ) ;
  assign n2625 = ( x70 & n2452 ) | ( x70 & ~n2584 ) | ( n2452 & ~n2584 ) ;
  assign n2626 = x70 & n2452 ;
  assign n2627 = ( ~n2457 & n2625 ) | ( ~n2457 & n2626 ) | ( n2625 & n2626 ) ;
  assign n2628 = ( n2457 & n2625 ) | ( n2457 & n2626 ) | ( n2625 & n2626 ) ;
  assign n2629 = ( n2457 & n2627 ) | ( n2457 & ~n2628 ) | ( n2627 & ~n2628 ) ;
  assign n2630 = ( x71 & n2624 ) | ( x71 & ~n2629 ) | ( n2624 & ~n2629 ) ;
  assign n2631 = ( x71 & n2458 ) | ( x71 & ~n2584 ) | ( n2458 & ~n2584 ) ;
  assign n2632 = x71 & n2458 ;
  assign n2633 = ( ~n2463 & n2631 ) | ( ~n2463 & n2632 ) | ( n2631 & n2632 ) ;
  assign n2634 = ( n2463 & n2631 ) | ( n2463 & n2632 ) | ( n2631 & n2632 ) ;
  assign n2635 = ( n2463 & n2633 ) | ( n2463 & ~n2634 ) | ( n2633 & ~n2634 ) ;
  assign n2636 = ( x72 & n2630 ) | ( x72 & ~n2635 ) | ( n2630 & ~n2635 ) ;
  assign n2637 = ( x72 & n2464 ) | ( x72 & ~n2584 ) | ( n2464 & ~n2584 ) ;
  assign n2638 = x72 & n2464 ;
  assign n2639 = ( ~n2469 & n2637 ) | ( ~n2469 & n2638 ) | ( n2637 & n2638 ) ;
  assign n2640 = ( n2469 & n2637 ) | ( n2469 & n2638 ) | ( n2637 & n2638 ) ;
  assign n2641 = ( n2469 & n2639 ) | ( n2469 & ~n2640 ) | ( n2639 & ~n2640 ) ;
  assign n2642 = ( x73 & n2636 ) | ( x73 & ~n2641 ) | ( n2636 & ~n2641 ) ;
  assign n2643 = ( x73 & n2470 ) | ( x73 & ~n2584 ) | ( n2470 & ~n2584 ) ;
  assign n2644 = x73 & n2470 ;
  assign n2645 = ( ~n2475 & n2643 ) | ( ~n2475 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2646 = ( n2475 & n2643 ) | ( n2475 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2647 = ( n2475 & n2645 ) | ( n2475 & ~n2646 ) | ( n2645 & ~n2646 ) ;
  assign n2648 = ( x74 & n2642 ) | ( x74 & ~n2647 ) | ( n2642 & ~n2647 ) ;
  assign n2649 = ( x74 & n2476 ) | ( x74 & ~n2584 ) | ( n2476 & ~n2584 ) ;
  assign n2650 = x74 & n2476 ;
  assign n2651 = ( ~n2481 & n2649 ) | ( ~n2481 & n2650 ) | ( n2649 & n2650 ) ;
  assign n2652 = ( n2481 & n2649 ) | ( n2481 & n2650 ) | ( n2649 & n2650 ) ;
  assign n2653 = ( n2481 & n2651 ) | ( n2481 & ~n2652 ) | ( n2651 & ~n2652 ) ;
  assign n2654 = ( x75 & n2648 ) | ( x75 & ~n2653 ) | ( n2648 & ~n2653 ) ;
  assign n2655 = ( x75 & n2482 ) | ( x75 & ~n2584 ) | ( n2482 & ~n2584 ) ;
  assign n2656 = x75 & n2482 ;
  assign n2657 = ( ~n2487 & n2655 ) | ( ~n2487 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = ( n2487 & n2655 ) | ( n2487 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2659 = ( n2487 & n2657 ) | ( n2487 & ~n2658 ) | ( n2657 & ~n2658 ) ;
  assign n2660 = ( x76 & n2654 ) | ( x76 & ~n2659 ) | ( n2654 & ~n2659 ) ;
  assign n2661 = ( x76 & n2488 ) | ( x76 & ~n2584 ) | ( n2488 & ~n2584 ) ;
  assign n2662 = x76 & n2488 ;
  assign n2663 = ( ~n2493 & n2661 ) | ( ~n2493 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2664 = ( n2493 & n2661 ) | ( n2493 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2665 = ( n2493 & n2663 ) | ( n2493 & ~n2664 ) | ( n2663 & ~n2664 ) ;
  assign n2666 = ( x77 & n2660 ) | ( x77 & ~n2665 ) | ( n2660 & ~n2665 ) ;
  assign n2667 = ( x77 & n2494 ) | ( x77 & ~n2584 ) | ( n2494 & ~n2584 ) ;
  assign n2668 = x77 & n2494 ;
  assign n2669 = ( ~n2499 & n2667 ) | ( ~n2499 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = ( n2499 & n2667 ) | ( n2499 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2671 = ( n2499 & n2669 ) | ( n2499 & ~n2670 ) | ( n2669 & ~n2670 ) ;
  assign n2672 = ( x78 & n2666 ) | ( x78 & ~n2671 ) | ( n2666 & ~n2671 ) ;
  assign n2673 = ( x78 & n2500 ) | ( x78 & ~n2584 ) | ( n2500 & ~n2584 ) ;
  assign n2674 = x78 & n2500 ;
  assign n2675 = ( ~n2505 & n2673 ) | ( ~n2505 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = ( n2505 & n2673 ) | ( n2505 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2677 = ( n2505 & n2675 ) | ( n2505 & ~n2676 ) | ( n2675 & ~n2676 ) ;
  assign n2678 = ( x79 & n2672 ) | ( x79 & ~n2677 ) | ( n2672 & ~n2677 ) ;
  assign n2679 = ( x79 & n2506 ) | ( x79 & ~n2584 ) | ( n2506 & ~n2584 ) ;
  assign n2680 = x79 & n2506 ;
  assign n2681 = ( ~n2511 & n2679 ) | ( ~n2511 & n2680 ) | ( n2679 & n2680 ) ;
  assign n2682 = ( n2511 & n2679 ) | ( n2511 & n2680 ) | ( n2679 & n2680 ) ;
  assign n2683 = ( n2511 & n2681 ) | ( n2511 & ~n2682 ) | ( n2681 & ~n2682 ) ;
  assign n2684 = ( x80 & n2678 ) | ( x80 & ~n2683 ) | ( n2678 & ~n2683 ) ;
  assign n2685 = ( x80 & n2512 ) | ( x80 & ~n2584 ) | ( n2512 & ~n2584 ) ;
  assign n2686 = x80 & n2512 ;
  assign n2687 = ( ~n2517 & n2685 ) | ( ~n2517 & n2686 ) | ( n2685 & n2686 ) ;
  assign n2688 = ( n2517 & n2685 ) | ( n2517 & n2686 ) | ( n2685 & n2686 ) ;
  assign n2689 = ( n2517 & n2687 ) | ( n2517 & ~n2688 ) | ( n2687 & ~n2688 ) ;
  assign n2690 = ( x81 & n2684 ) | ( x81 & ~n2689 ) | ( n2684 & ~n2689 ) ;
  assign n2691 = ( x81 & n2518 ) | ( x81 & ~n2584 ) | ( n2518 & ~n2584 ) ;
  assign n2692 = x81 & n2518 ;
  assign n2693 = ( ~n2523 & n2691 ) | ( ~n2523 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2694 = ( n2523 & n2691 ) | ( n2523 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2695 = ( n2523 & n2693 ) | ( n2523 & ~n2694 ) | ( n2693 & ~n2694 ) ;
  assign n2696 = ( x82 & n2690 ) | ( x82 & ~n2695 ) | ( n2690 & ~n2695 ) ;
  assign n2697 = ( x82 & n2524 ) | ( x82 & ~n2584 ) | ( n2524 & ~n2584 ) ;
  assign n2698 = x82 & n2524 ;
  assign n2699 = ( ~n2529 & n2697 ) | ( ~n2529 & n2698 ) | ( n2697 & n2698 ) ;
  assign n2700 = ( n2529 & n2697 ) | ( n2529 & n2698 ) | ( n2697 & n2698 ) ;
  assign n2701 = ( n2529 & n2699 ) | ( n2529 & ~n2700 ) | ( n2699 & ~n2700 ) ;
  assign n2702 = ( x83 & n2696 ) | ( x83 & ~n2701 ) | ( n2696 & ~n2701 ) ;
  assign n2703 = ( x83 & n2530 ) | ( x83 & ~n2584 ) | ( n2530 & ~n2584 ) ;
  assign n2704 = x83 & n2530 ;
  assign n2705 = ( ~n2535 & n2703 ) | ( ~n2535 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2706 = ( n2535 & n2703 ) | ( n2535 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2707 = ( n2535 & n2705 ) | ( n2535 & ~n2706 ) | ( n2705 & ~n2706 ) ;
  assign n2708 = ( x84 & n2702 ) | ( x84 & ~n2707 ) | ( n2702 & ~n2707 ) ;
  assign n2709 = ( x84 & n2536 ) | ( x84 & ~n2584 ) | ( n2536 & ~n2584 ) ;
  assign n2710 = x84 & n2536 ;
  assign n2711 = ( ~n2541 & n2709 ) | ( ~n2541 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2712 = ( n2541 & n2709 ) | ( n2541 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2713 = ( n2541 & n2711 ) | ( n2541 & ~n2712 ) | ( n2711 & ~n2712 ) ;
  assign n2714 = ( x85 & n2708 ) | ( x85 & ~n2713 ) | ( n2708 & ~n2713 ) ;
  assign n2715 = ( x85 & n2542 ) | ( x85 & ~n2584 ) | ( n2542 & ~n2584 ) ;
  assign n2716 = x85 & n2542 ;
  assign n2717 = ( ~n2547 & n2715 ) | ( ~n2547 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2718 = ( n2547 & n2715 ) | ( n2547 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2719 = ( n2547 & n2717 ) | ( n2547 & ~n2718 ) | ( n2717 & ~n2718 ) ;
  assign n2720 = ( x86 & n2714 ) | ( x86 & ~n2719 ) | ( n2714 & ~n2719 ) ;
  assign n2721 = ( x86 & n2548 ) | ( x86 & ~n2584 ) | ( n2548 & ~n2584 ) ;
  assign n2722 = x86 & n2548 ;
  assign n2723 = ( ~n2553 & n2721 ) | ( ~n2553 & n2722 ) | ( n2721 & n2722 ) ;
  assign n2724 = ( n2553 & n2721 ) | ( n2553 & n2722 ) | ( n2721 & n2722 ) ;
  assign n2725 = ( n2553 & n2723 ) | ( n2553 & ~n2724 ) | ( n2723 & ~n2724 ) ;
  assign n2726 = ( x87 & n2720 ) | ( x87 & ~n2725 ) | ( n2720 & ~n2725 ) ;
  assign n2727 = ( x87 & n2554 ) | ( x87 & ~n2584 ) | ( n2554 & ~n2584 ) ;
  assign n2728 = x87 & n2554 ;
  assign n2729 = ( ~n2559 & n2727 ) | ( ~n2559 & n2728 ) | ( n2727 & n2728 ) ;
  assign n2730 = ( n2559 & n2727 ) | ( n2559 & n2728 ) | ( n2727 & n2728 ) ;
  assign n2731 = ( n2559 & n2729 ) | ( n2559 & ~n2730 ) | ( n2729 & ~n2730 ) ;
  assign n2732 = ( x88 & n2726 ) | ( x88 & ~n2731 ) | ( n2726 & ~n2731 ) ;
  assign n2733 = ( x88 & n2560 ) | ( x88 & ~n2584 ) | ( n2560 & ~n2584 ) ;
  assign n2734 = x88 & n2560 ;
  assign n2735 = ( ~n2565 & n2733 ) | ( ~n2565 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2736 = ( n2565 & n2733 ) | ( n2565 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2737 = ( n2565 & n2735 ) | ( n2565 & ~n2736 ) | ( n2735 & ~n2736 ) ;
  assign n2738 = ( x89 & n2732 ) | ( x89 & ~n2737 ) | ( n2732 & ~n2737 ) ;
  assign n2739 = ( x89 & n2566 ) | ( x89 & ~n2584 ) | ( n2566 & ~n2584 ) ;
  assign n2740 = x89 & n2566 ;
  assign n2741 = ( ~n2571 & n2739 ) | ( ~n2571 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2742 = ( n2571 & n2739 ) | ( n2571 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2743 = ( n2571 & n2741 ) | ( n2571 & ~n2742 ) | ( n2741 & ~n2742 ) ;
  assign n2744 = ( x90 & n2738 ) | ( x90 & ~n2743 ) | ( n2738 & ~n2743 ) ;
  assign n2745 = ( x90 & n2572 ) | ( x90 & ~n2584 ) | ( n2572 & ~n2584 ) ;
  assign n2746 = x90 & n2572 ;
  assign n2747 = ( ~n2577 & n2745 ) | ( ~n2577 & n2746 ) | ( n2745 & n2746 ) ;
  assign n2748 = ( n2577 & n2745 ) | ( n2577 & n2746 ) | ( n2745 & n2746 ) ;
  assign n2749 = ( n2577 & n2747 ) | ( n2577 & ~n2748 ) | ( n2747 & ~n2748 ) ;
  assign n2750 = ( x91 & n2744 ) | ( x91 & ~n2749 ) | ( n2744 & ~n2749 ) ;
  assign n2751 = ( n163 & n164 ) | ( n163 & ~n2581 ) | ( n164 & ~n2581 ) ;
  assign n2752 = ( ~x92 & x93 ) | ( ~x92 & n2582 ) | ( x93 & n2582 ) ;
  assign n2753 = ( ~x92 & n2581 ) | ( ~x92 & n2582 ) | ( n2581 & n2582 ) ;
  assign n2754 = ~n2752 & n2753 ;
  assign n2755 = ( x92 & ~n2589 ) | ( x92 & n2750 ) | ( ~n2589 & n2750 ) ;
  assign n2756 = ~n2754 & n2755 ;
  assign n2757 = n2751 | n2756 ;
  assign n2758 = ( x92 & n2750 ) | ( x92 & n2757 ) | ( n2750 & n2757 ) ;
  assign n2759 = x92 | n2750 ;
  assign n2760 = ( ~n2589 & n2758 ) | ( ~n2589 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = ( n2589 & n2758 ) | ( n2589 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2762 = ( n2589 & n2760 ) | ( n2589 & ~n2761 ) | ( n2760 & ~n2761 ) ;
  assign n2763 = ~x33 & x64 ;
  assign n2764 = ~x34 & n2757 ;
  assign n2765 = ( x34 & ~x64 ) | ( x34 & n2757 ) | ( ~x64 & n2757 ) ;
  assign n2766 = ( n2590 & ~n2764 ) | ( n2590 & n2765 ) | ( ~n2764 & n2765 ) ;
  assign n2767 = ( x65 & n2763 ) | ( x65 & ~n2766 ) | ( n2763 & ~n2766 ) ;
  assign n2768 = ( x65 & n2590 ) | ( x65 & n2757 ) | ( n2590 & n2757 ) ;
  assign n2769 = x65 | n2590 ;
  assign n2770 = ( ~n2593 & n2768 ) | ( ~n2593 & n2769 ) | ( n2768 & n2769 ) ;
  assign n2771 = ( n2593 & n2768 ) | ( n2593 & n2769 ) | ( n2768 & n2769 ) ;
  assign n2772 = ( n2593 & n2770 ) | ( n2593 & ~n2771 ) | ( n2770 & ~n2771 ) ;
  assign n2773 = ( x66 & n2767 ) | ( x66 & ~n2772 ) | ( n2767 & ~n2772 ) ;
  assign n2774 = ( x66 & n2594 ) | ( x66 & n2757 ) | ( n2594 & n2757 ) ;
  assign n2775 = x66 | n2594 ;
  assign n2776 = ( ~n2599 & n2774 ) | ( ~n2599 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2777 = ( n2599 & n2774 ) | ( n2599 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2778 = ( n2599 & n2776 ) | ( n2599 & ~n2777 ) | ( n2776 & ~n2777 ) ;
  assign n2779 = ( x67 & n2773 ) | ( x67 & ~n2778 ) | ( n2773 & ~n2778 ) ;
  assign n2780 = ( x67 & n2600 ) | ( x67 & ~n2757 ) | ( n2600 & ~n2757 ) ;
  assign n2781 = x67 & n2600 ;
  assign n2782 = ( ~n2605 & n2780 ) | ( ~n2605 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2783 = ( n2605 & n2780 ) | ( n2605 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2784 = ( n2605 & n2782 ) | ( n2605 & ~n2783 ) | ( n2782 & ~n2783 ) ;
  assign n2785 = ( x68 & n2779 ) | ( x68 & ~n2784 ) | ( n2779 & ~n2784 ) ;
  assign n2786 = ( x68 & n2606 ) | ( x68 & ~n2757 ) | ( n2606 & ~n2757 ) ;
  assign n2787 = x68 & n2606 ;
  assign n2788 = ( ~n2611 & n2786 ) | ( ~n2611 & n2787 ) | ( n2786 & n2787 ) ;
  assign n2789 = ( n2611 & n2786 ) | ( n2611 & n2787 ) | ( n2786 & n2787 ) ;
  assign n2790 = ( n2611 & n2788 ) | ( n2611 & ~n2789 ) | ( n2788 & ~n2789 ) ;
  assign n2791 = ( x69 & n2785 ) | ( x69 & ~n2790 ) | ( n2785 & ~n2790 ) ;
  assign n2792 = ( x69 & n2612 ) | ( x69 & ~n2757 ) | ( n2612 & ~n2757 ) ;
  assign n2793 = x69 & n2612 ;
  assign n2794 = ( ~n2617 & n2792 ) | ( ~n2617 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2795 = ( n2617 & n2792 ) | ( n2617 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2796 = ( n2617 & n2794 ) | ( n2617 & ~n2795 ) | ( n2794 & ~n2795 ) ;
  assign n2797 = ( x70 & n2791 ) | ( x70 & ~n2796 ) | ( n2791 & ~n2796 ) ;
  assign n2798 = ( x70 & n2618 ) | ( x70 & ~n2757 ) | ( n2618 & ~n2757 ) ;
  assign n2799 = x70 & n2618 ;
  assign n2800 = ( ~n2623 & n2798 ) | ( ~n2623 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = ( n2623 & n2798 ) | ( n2623 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2802 = ( n2623 & n2800 ) | ( n2623 & ~n2801 ) | ( n2800 & ~n2801 ) ;
  assign n2803 = ( x71 & n2797 ) | ( x71 & ~n2802 ) | ( n2797 & ~n2802 ) ;
  assign n2804 = ( x71 & n2624 ) | ( x71 & ~n2757 ) | ( n2624 & ~n2757 ) ;
  assign n2805 = x71 & n2624 ;
  assign n2806 = ( ~n2629 & n2804 ) | ( ~n2629 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2807 = ( n2629 & n2804 ) | ( n2629 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2808 = ( n2629 & n2806 ) | ( n2629 & ~n2807 ) | ( n2806 & ~n2807 ) ;
  assign n2809 = ( x72 & n2803 ) | ( x72 & ~n2808 ) | ( n2803 & ~n2808 ) ;
  assign n2810 = ( x72 & n2630 ) | ( x72 & ~n2757 ) | ( n2630 & ~n2757 ) ;
  assign n2811 = x72 & n2630 ;
  assign n2812 = ( ~n2635 & n2810 ) | ( ~n2635 & n2811 ) | ( n2810 & n2811 ) ;
  assign n2813 = ( n2635 & n2810 ) | ( n2635 & n2811 ) | ( n2810 & n2811 ) ;
  assign n2814 = ( n2635 & n2812 ) | ( n2635 & ~n2813 ) | ( n2812 & ~n2813 ) ;
  assign n2815 = ( x73 & n2809 ) | ( x73 & ~n2814 ) | ( n2809 & ~n2814 ) ;
  assign n2816 = ( x73 & n2636 ) | ( x73 & ~n2757 ) | ( n2636 & ~n2757 ) ;
  assign n2817 = x73 & n2636 ;
  assign n2818 = ( ~n2641 & n2816 ) | ( ~n2641 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2819 = ( n2641 & n2816 ) | ( n2641 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2820 = ( n2641 & n2818 ) | ( n2641 & ~n2819 ) | ( n2818 & ~n2819 ) ;
  assign n2821 = ( x74 & n2815 ) | ( x74 & ~n2820 ) | ( n2815 & ~n2820 ) ;
  assign n2822 = ( x74 & n2642 ) | ( x74 & ~n2757 ) | ( n2642 & ~n2757 ) ;
  assign n2823 = x74 & n2642 ;
  assign n2824 = ( ~n2647 & n2822 ) | ( ~n2647 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = ( n2647 & n2822 ) | ( n2647 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2826 = ( n2647 & n2824 ) | ( n2647 & ~n2825 ) | ( n2824 & ~n2825 ) ;
  assign n2827 = ( x75 & n2821 ) | ( x75 & ~n2826 ) | ( n2821 & ~n2826 ) ;
  assign n2828 = ( x75 & n2648 ) | ( x75 & ~n2757 ) | ( n2648 & ~n2757 ) ;
  assign n2829 = x75 & n2648 ;
  assign n2830 = ( ~n2653 & n2828 ) | ( ~n2653 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( n2653 & n2828 ) | ( n2653 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2832 = ( n2653 & n2830 ) | ( n2653 & ~n2831 ) | ( n2830 & ~n2831 ) ;
  assign n2833 = ( x76 & n2827 ) | ( x76 & ~n2832 ) | ( n2827 & ~n2832 ) ;
  assign n2834 = ( x76 & n2654 ) | ( x76 & ~n2757 ) | ( n2654 & ~n2757 ) ;
  assign n2835 = x76 & n2654 ;
  assign n2836 = ( ~n2659 & n2834 ) | ( ~n2659 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2837 = ( n2659 & n2834 ) | ( n2659 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2838 = ( n2659 & n2836 ) | ( n2659 & ~n2837 ) | ( n2836 & ~n2837 ) ;
  assign n2839 = ( x77 & n2833 ) | ( x77 & ~n2838 ) | ( n2833 & ~n2838 ) ;
  assign n2840 = ( x77 & n2660 ) | ( x77 & ~n2757 ) | ( n2660 & ~n2757 ) ;
  assign n2841 = x77 & n2660 ;
  assign n2842 = ( ~n2665 & n2840 ) | ( ~n2665 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2843 = ( n2665 & n2840 ) | ( n2665 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2844 = ( n2665 & n2842 ) | ( n2665 & ~n2843 ) | ( n2842 & ~n2843 ) ;
  assign n2845 = ( x78 & n2839 ) | ( x78 & ~n2844 ) | ( n2839 & ~n2844 ) ;
  assign n2846 = ( x78 & n2666 ) | ( x78 & ~n2757 ) | ( n2666 & ~n2757 ) ;
  assign n2847 = x78 & n2666 ;
  assign n2848 = ( ~n2671 & n2846 ) | ( ~n2671 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = ( n2671 & n2846 ) | ( n2671 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2850 = ( n2671 & n2848 ) | ( n2671 & ~n2849 ) | ( n2848 & ~n2849 ) ;
  assign n2851 = ( x79 & n2845 ) | ( x79 & ~n2850 ) | ( n2845 & ~n2850 ) ;
  assign n2852 = ( x79 & n2672 ) | ( x79 & ~n2757 ) | ( n2672 & ~n2757 ) ;
  assign n2853 = x79 & n2672 ;
  assign n2854 = ( ~n2677 & n2852 ) | ( ~n2677 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = ( n2677 & n2852 ) | ( n2677 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2856 = ( n2677 & n2854 ) | ( n2677 & ~n2855 ) | ( n2854 & ~n2855 ) ;
  assign n2857 = ( x80 & n2851 ) | ( x80 & ~n2856 ) | ( n2851 & ~n2856 ) ;
  assign n2858 = ( x80 & n2678 ) | ( x80 & ~n2757 ) | ( n2678 & ~n2757 ) ;
  assign n2859 = x80 & n2678 ;
  assign n2860 = ( ~n2683 & n2858 ) | ( ~n2683 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2861 = ( n2683 & n2858 ) | ( n2683 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2862 = ( n2683 & n2860 ) | ( n2683 & ~n2861 ) | ( n2860 & ~n2861 ) ;
  assign n2863 = ( x81 & n2857 ) | ( x81 & ~n2862 ) | ( n2857 & ~n2862 ) ;
  assign n2864 = ( x81 & n2684 ) | ( x81 & ~n2757 ) | ( n2684 & ~n2757 ) ;
  assign n2865 = x81 & n2684 ;
  assign n2866 = ( ~n2689 & n2864 ) | ( ~n2689 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2867 = ( n2689 & n2864 ) | ( n2689 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2868 = ( n2689 & n2866 ) | ( n2689 & ~n2867 ) | ( n2866 & ~n2867 ) ;
  assign n2869 = ( x82 & n2863 ) | ( x82 & ~n2868 ) | ( n2863 & ~n2868 ) ;
  assign n2870 = ( x82 & n2690 ) | ( x82 & ~n2757 ) | ( n2690 & ~n2757 ) ;
  assign n2871 = x82 & n2690 ;
  assign n2872 = ( ~n2695 & n2870 ) | ( ~n2695 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2873 = ( n2695 & n2870 ) | ( n2695 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2874 = ( n2695 & n2872 ) | ( n2695 & ~n2873 ) | ( n2872 & ~n2873 ) ;
  assign n2875 = ( x83 & n2869 ) | ( x83 & ~n2874 ) | ( n2869 & ~n2874 ) ;
  assign n2876 = ( x83 & n2696 ) | ( x83 & ~n2757 ) | ( n2696 & ~n2757 ) ;
  assign n2877 = x83 & n2696 ;
  assign n2878 = ( ~n2701 & n2876 ) | ( ~n2701 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2879 = ( n2701 & n2876 ) | ( n2701 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2880 = ( n2701 & n2878 ) | ( n2701 & ~n2879 ) | ( n2878 & ~n2879 ) ;
  assign n2881 = ( x84 & n2875 ) | ( x84 & ~n2880 ) | ( n2875 & ~n2880 ) ;
  assign n2882 = ( x84 & n2702 ) | ( x84 & ~n2757 ) | ( n2702 & ~n2757 ) ;
  assign n2883 = x84 & n2702 ;
  assign n2884 = ( ~n2707 & n2882 ) | ( ~n2707 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = ( n2707 & n2882 ) | ( n2707 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2886 = ( n2707 & n2884 ) | ( n2707 & ~n2885 ) | ( n2884 & ~n2885 ) ;
  assign n2887 = ( x85 & n2881 ) | ( x85 & ~n2886 ) | ( n2881 & ~n2886 ) ;
  assign n2888 = ( x85 & n2708 ) | ( x85 & ~n2757 ) | ( n2708 & ~n2757 ) ;
  assign n2889 = x85 & n2708 ;
  assign n2890 = ( ~n2713 & n2888 ) | ( ~n2713 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2891 = ( n2713 & n2888 ) | ( n2713 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2892 = ( n2713 & n2890 ) | ( n2713 & ~n2891 ) | ( n2890 & ~n2891 ) ;
  assign n2893 = ( x86 & n2887 ) | ( x86 & ~n2892 ) | ( n2887 & ~n2892 ) ;
  assign n2894 = ( x86 & n2714 ) | ( x86 & ~n2757 ) | ( n2714 & ~n2757 ) ;
  assign n2895 = x86 & n2714 ;
  assign n2896 = ( ~n2719 & n2894 ) | ( ~n2719 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2897 = ( n2719 & n2894 ) | ( n2719 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2898 = ( n2719 & n2896 ) | ( n2719 & ~n2897 ) | ( n2896 & ~n2897 ) ;
  assign n2899 = ( x87 & n2893 ) | ( x87 & ~n2898 ) | ( n2893 & ~n2898 ) ;
  assign n2900 = ( x87 & n2720 ) | ( x87 & ~n2757 ) | ( n2720 & ~n2757 ) ;
  assign n2901 = x87 & n2720 ;
  assign n2902 = ( ~n2725 & n2900 ) | ( ~n2725 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2903 = ( n2725 & n2900 ) | ( n2725 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2904 = ( n2725 & n2902 ) | ( n2725 & ~n2903 ) | ( n2902 & ~n2903 ) ;
  assign n2905 = ( x88 & n2899 ) | ( x88 & ~n2904 ) | ( n2899 & ~n2904 ) ;
  assign n2906 = ( x88 & n2726 ) | ( x88 & ~n2757 ) | ( n2726 & ~n2757 ) ;
  assign n2907 = x88 & n2726 ;
  assign n2908 = ( ~n2731 & n2906 ) | ( ~n2731 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ( n2731 & n2906 ) | ( n2731 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2910 = ( n2731 & n2908 ) | ( n2731 & ~n2909 ) | ( n2908 & ~n2909 ) ;
  assign n2911 = ( x89 & n2905 ) | ( x89 & ~n2910 ) | ( n2905 & ~n2910 ) ;
  assign n2912 = ( x89 & n2732 ) | ( x89 & ~n2757 ) | ( n2732 & ~n2757 ) ;
  assign n2913 = x89 & n2732 ;
  assign n2914 = ( ~n2737 & n2912 ) | ( ~n2737 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = ( n2737 & n2912 ) | ( n2737 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2916 = ( n2737 & n2914 ) | ( n2737 & ~n2915 ) | ( n2914 & ~n2915 ) ;
  assign n2917 = ( x90 & n2911 ) | ( x90 & ~n2916 ) | ( n2911 & ~n2916 ) ;
  assign n2918 = ( x90 & n2738 ) | ( x90 & ~n2757 ) | ( n2738 & ~n2757 ) ;
  assign n2919 = x90 & n2738 ;
  assign n2920 = ( ~n2743 & n2918 ) | ( ~n2743 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2921 = ( n2743 & n2918 ) | ( n2743 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2922 = ( n2743 & n2920 ) | ( n2743 & ~n2921 ) | ( n2920 & ~n2921 ) ;
  assign n2923 = ( x91 & n2917 ) | ( x91 & ~n2922 ) | ( n2917 & ~n2922 ) ;
  assign n2924 = ( x91 & n2744 ) | ( x91 & ~n2757 ) | ( n2744 & ~n2757 ) ;
  assign n2925 = x91 & n2744 ;
  assign n2926 = ( ~n2749 & n2924 ) | ( ~n2749 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2927 = ( n2749 & n2924 ) | ( n2749 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2928 = ( n2749 & n2926 ) | ( n2749 & ~n2927 ) | ( n2926 & ~n2927 ) ;
  assign n2929 = ( x92 & n2923 ) | ( x92 & ~n2928 ) | ( n2923 & ~n2928 ) ;
  assign n2930 = ( x93 & ~n2762 ) | ( x93 & n2929 ) | ( ~n2762 & n2929 ) ;
  assign n2931 = ~n164 & n2755 ;
  assign n2932 = n163 & n2581 ;
  assign n2933 = ( n2581 & n2755 ) | ( n2581 & n2932 ) | ( n2755 & n2932 ) ;
  assign n2934 = n2754 | n2933 ;
  assign n2935 = ~n2931 & n2934 ;
  assign n2936 = ( x94 & n2930 ) | ( x94 & ~n2935 ) | ( n2930 & ~n2935 ) ;
  assign n2937 = n162 | n2936 ;
  assign n2938 = ( x93 & n2929 ) | ( x93 & n2937 ) | ( n2929 & n2937 ) ;
  assign n2939 = x93 | n2929 ;
  assign n2940 = ( ~n2762 & n2938 ) | ( ~n2762 & n2939 ) | ( n2938 & n2939 ) ;
  assign n2941 = ( n2762 & n2938 ) | ( n2762 & n2939 ) | ( n2938 & n2939 ) ;
  assign n2942 = ( n2762 & n2940 ) | ( n2762 & ~n2941 ) | ( n2940 & ~n2941 ) ;
  assign n2943 = ~x32 & x64 ;
  assign n2944 = ~x33 & n2937 ;
  assign n2945 = ( x33 & ~x64 ) | ( x33 & n2937 ) | ( ~x64 & n2937 ) ;
  assign n2946 = ( n2763 & ~n2944 ) | ( n2763 & n2945 ) | ( ~n2944 & n2945 ) ;
  assign n2947 = ( x65 & n2943 ) | ( x65 & ~n2946 ) | ( n2943 & ~n2946 ) ;
  assign n2948 = ( x65 & n2763 ) | ( x65 & n2937 ) | ( n2763 & n2937 ) ;
  assign n2949 = x65 | n2763 ;
  assign n2950 = ( ~n2766 & n2948 ) | ( ~n2766 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2951 = ( n2766 & n2948 ) | ( n2766 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2952 = ( n2766 & n2950 ) | ( n2766 & ~n2951 ) | ( n2950 & ~n2951 ) ;
  assign n2953 = ( x66 & n2947 ) | ( x66 & ~n2952 ) | ( n2947 & ~n2952 ) ;
  assign n2954 = ( x66 & n2767 ) | ( x66 & n2937 ) | ( n2767 & n2937 ) ;
  assign n2955 = x66 | n2767 ;
  assign n2956 = ( ~n2772 & n2954 ) | ( ~n2772 & n2955 ) | ( n2954 & n2955 ) ;
  assign n2957 = ( n2772 & n2954 ) | ( n2772 & n2955 ) | ( n2954 & n2955 ) ;
  assign n2958 = ( n2772 & n2956 ) | ( n2772 & ~n2957 ) | ( n2956 & ~n2957 ) ;
  assign n2959 = ( x67 & n2953 ) | ( x67 & ~n2958 ) | ( n2953 & ~n2958 ) ;
  assign n2960 = ( x67 & n2773 ) | ( x67 & ~n2937 ) | ( n2773 & ~n2937 ) ;
  assign n2961 = x67 & n2773 ;
  assign n2962 = ( ~n2778 & n2960 ) | ( ~n2778 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2963 = ( n2778 & n2960 ) | ( n2778 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2964 = ( n2778 & n2962 ) | ( n2778 & ~n2963 ) | ( n2962 & ~n2963 ) ;
  assign n2965 = ( x68 & n2959 ) | ( x68 & ~n2964 ) | ( n2959 & ~n2964 ) ;
  assign n2966 = ( x68 & n2779 ) | ( x68 & ~n2937 ) | ( n2779 & ~n2937 ) ;
  assign n2967 = x68 & n2779 ;
  assign n2968 = ( ~n2784 & n2966 ) | ( ~n2784 & n2967 ) | ( n2966 & n2967 ) ;
  assign n2969 = ( n2784 & n2966 ) | ( n2784 & n2967 ) | ( n2966 & n2967 ) ;
  assign n2970 = ( n2784 & n2968 ) | ( n2784 & ~n2969 ) | ( n2968 & ~n2969 ) ;
  assign n2971 = ( x69 & n2965 ) | ( x69 & ~n2970 ) | ( n2965 & ~n2970 ) ;
  assign n2972 = ( x69 & n2785 ) | ( x69 & ~n2937 ) | ( n2785 & ~n2937 ) ;
  assign n2973 = x69 & n2785 ;
  assign n2974 = ( ~n2790 & n2972 ) | ( ~n2790 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = ( n2790 & n2972 ) | ( n2790 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2976 = ( n2790 & n2974 ) | ( n2790 & ~n2975 ) | ( n2974 & ~n2975 ) ;
  assign n2977 = ( x70 & n2971 ) | ( x70 & ~n2976 ) | ( n2971 & ~n2976 ) ;
  assign n2978 = ( x70 & n2791 ) | ( x70 & ~n2937 ) | ( n2791 & ~n2937 ) ;
  assign n2979 = x70 & n2791 ;
  assign n2980 = ( ~n2796 & n2978 ) | ( ~n2796 & n2979 ) | ( n2978 & n2979 ) ;
  assign n2981 = ( n2796 & n2978 ) | ( n2796 & n2979 ) | ( n2978 & n2979 ) ;
  assign n2982 = ( n2796 & n2980 ) | ( n2796 & ~n2981 ) | ( n2980 & ~n2981 ) ;
  assign n2983 = ( x71 & n2977 ) | ( x71 & ~n2982 ) | ( n2977 & ~n2982 ) ;
  assign n2984 = ( x71 & n2797 ) | ( x71 & ~n2937 ) | ( n2797 & ~n2937 ) ;
  assign n2985 = x71 & n2797 ;
  assign n2986 = ( ~n2802 & n2984 ) | ( ~n2802 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = ( n2802 & n2984 ) | ( n2802 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2988 = ( n2802 & n2986 ) | ( n2802 & ~n2987 ) | ( n2986 & ~n2987 ) ;
  assign n2989 = ( x72 & n2983 ) | ( x72 & ~n2988 ) | ( n2983 & ~n2988 ) ;
  assign n2990 = ( x72 & n2803 ) | ( x72 & ~n2937 ) | ( n2803 & ~n2937 ) ;
  assign n2991 = x72 & n2803 ;
  assign n2992 = ( ~n2808 & n2990 ) | ( ~n2808 & n2991 ) | ( n2990 & n2991 ) ;
  assign n2993 = ( n2808 & n2990 ) | ( n2808 & n2991 ) | ( n2990 & n2991 ) ;
  assign n2994 = ( n2808 & n2992 ) | ( n2808 & ~n2993 ) | ( n2992 & ~n2993 ) ;
  assign n2995 = ( x73 & n2989 ) | ( x73 & ~n2994 ) | ( n2989 & ~n2994 ) ;
  assign n2996 = ( x73 & n2809 ) | ( x73 & ~n2937 ) | ( n2809 & ~n2937 ) ;
  assign n2997 = x73 & n2809 ;
  assign n2998 = ( ~n2814 & n2996 ) | ( ~n2814 & n2997 ) | ( n2996 & n2997 ) ;
  assign n2999 = ( n2814 & n2996 ) | ( n2814 & n2997 ) | ( n2996 & n2997 ) ;
  assign n3000 = ( n2814 & n2998 ) | ( n2814 & ~n2999 ) | ( n2998 & ~n2999 ) ;
  assign n3001 = ( x74 & n2995 ) | ( x74 & ~n3000 ) | ( n2995 & ~n3000 ) ;
  assign n3002 = ( x74 & n2815 ) | ( x74 & ~n2937 ) | ( n2815 & ~n2937 ) ;
  assign n3003 = x74 & n2815 ;
  assign n3004 = ( ~n2820 & n3002 ) | ( ~n2820 & n3003 ) | ( n3002 & n3003 ) ;
  assign n3005 = ( n2820 & n3002 ) | ( n2820 & n3003 ) | ( n3002 & n3003 ) ;
  assign n3006 = ( n2820 & n3004 ) | ( n2820 & ~n3005 ) | ( n3004 & ~n3005 ) ;
  assign n3007 = ( x75 & n3001 ) | ( x75 & ~n3006 ) | ( n3001 & ~n3006 ) ;
  assign n3008 = ( x75 & n2821 ) | ( x75 & ~n2937 ) | ( n2821 & ~n2937 ) ;
  assign n3009 = x75 & n2821 ;
  assign n3010 = ( ~n2826 & n3008 ) | ( ~n2826 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3011 = ( n2826 & n3008 ) | ( n2826 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3012 = ( n2826 & n3010 ) | ( n2826 & ~n3011 ) | ( n3010 & ~n3011 ) ;
  assign n3013 = ( x76 & n3007 ) | ( x76 & ~n3012 ) | ( n3007 & ~n3012 ) ;
  assign n3014 = ( x76 & n2827 ) | ( x76 & ~n2937 ) | ( n2827 & ~n2937 ) ;
  assign n3015 = x76 & n2827 ;
  assign n3016 = ( ~n2832 & n3014 ) | ( ~n2832 & n3015 ) | ( n3014 & n3015 ) ;
  assign n3017 = ( n2832 & n3014 ) | ( n2832 & n3015 ) | ( n3014 & n3015 ) ;
  assign n3018 = ( n2832 & n3016 ) | ( n2832 & ~n3017 ) | ( n3016 & ~n3017 ) ;
  assign n3019 = ( x77 & n3013 ) | ( x77 & ~n3018 ) | ( n3013 & ~n3018 ) ;
  assign n3020 = ( x77 & n2833 ) | ( x77 & ~n2937 ) | ( n2833 & ~n2937 ) ;
  assign n3021 = x77 & n2833 ;
  assign n3022 = ( ~n2838 & n3020 ) | ( ~n2838 & n3021 ) | ( n3020 & n3021 ) ;
  assign n3023 = ( n2838 & n3020 ) | ( n2838 & n3021 ) | ( n3020 & n3021 ) ;
  assign n3024 = ( n2838 & n3022 ) | ( n2838 & ~n3023 ) | ( n3022 & ~n3023 ) ;
  assign n3025 = ( x78 & n3019 ) | ( x78 & ~n3024 ) | ( n3019 & ~n3024 ) ;
  assign n3026 = ( x78 & n2839 ) | ( x78 & ~n2937 ) | ( n2839 & ~n2937 ) ;
  assign n3027 = x78 & n2839 ;
  assign n3028 = ( ~n2844 & n3026 ) | ( ~n2844 & n3027 ) | ( n3026 & n3027 ) ;
  assign n3029 = ( n2844 & n3026 ) | ( n2844 & n3027 ) | ( n3026 & n3027 ) ;
  assign n3030 = ( n2844 & n3028 ) | ( n2844 & ~n3029 ) | ( n3028 & ~n3029 ) ;
  assign n3031 = ( x79 & n3025 ) | ( x79 & ~n3030 ) | ( n3025 & ~n3030 ) ;
  assign n3032 = ( x79 & n2845 ) | ( x79 & ~n2937 ) | ( n2845 & ~n2937 ) ;
  assign n3033 = x79 & n2845 ;
  assign n3034 = ( ~n2850 & n3032 ) | ( ~n2850 & n3033 ) | ( n3032 & n3033 ) ;
  assign n3035 = ( n2850 & n3032 ) | ( n2850 & n3033 ) | ( n3032 & n3033 ) ;
  assign n3036 = ( n2850 & n3034 ) | ( n2850 & ~n3035 ) | ( n3034 & ~n3035 ) ;
  assign n3037 = ( x80 & n3031 ) | ( x80 & ~n3036 ) | ( n3031 & ~n3036 ) ;
  assign n3038 = ( x80 & n2851 ) | ( x80 & ~n2937 ) | ( n2851 & ~n2937 ) ;
  assign n3039 = x80 & n2851 ;
  assign n3040 = ( ~n2856 & n3038 ) | ( ~n2856 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3041 = ( n2856 & n3038 ) | ( n2856 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3042 = ( n2856 & n3040 ) | ( n2856 & ~n3041 ) | ( n3040 & ~n3041 ) ;
  assign n3043 = ( x81 & n3037 ) | ( x81 & ~n3042 ) | ( n3037 & ~n3042 ) ;
  assign n3044 = ( x81 & n2857 ) | ( x81 & ~n2937 ) | ( n2857 & ~n2937 ) ;
  assign n3045 = x81 & n2857 ;
  assign n3046 = ( ~n2862 & n3044 ) | ( ~n2862 & n3045 ) | ( n3044 & n3045 ) ;
  assign n3047 = ( n2862 & n3044 ) | ( n2862 & n3045 ) | ( n3044 & n3045 ) ;
  assign n3048 = ( n2862 & n3046 ) | ( n2862 & ~n3047 ) | ( n3046 & ~n3047 ) ;
  assign n3049 = ( x82 & n3043 ) | ( x82 & ~n3048 ) | ( n3043 & ~n3048 ) ;
  assign n3050 = ( x82 & n2863 ) | ( x82 & ~n2937 ) | ( n2863 & ~n2937 ) ;
  assign n3051 = x82 & n2863 ;
  assign n3052 = ( ~n2868 & n3050 ) | ( ~n2868 & n3051 ) | ( n3050 & n3051 ) ;
  assign n3053 = ( n2868 & n3050 ) | ( n2868 & n3051 ) | ( n3050 & n3051 ) ;
  assign n3054 = ( n2868 & n3052 ) | ( n2868 & ~n3053 ) | ( n3052 & ~n3053 ) ;
  assign n3055 = ( x83 & n3049 ) | ( x83 & ~n3054 ) | ( n3049 & ~n3054 ) ;
  assign n3056 = ( x83 & n2869 ) | ( x83 & ~n2937 ) | ( n2869 & ~n2937 ) ;
  assign n3057 = x83 & n2869 ;
  assign n3058 = ( ~n2874 & n3056 ) | ( ~n2874 & n3057 ) | ( n3056 & n3057 ) ;
  assign n3059 = ( n2874 & n3056 ) | ( n2874 & n3057 ) | ( n3056 & n3057 ) ;
  assign n3060 = ( n2874 & n3058 ) | ( n2874 & ~n3059 ) | ( n3058 & ~n3059 ) ;
  assign n3061 = ( x84 & n3055 ) | ( x84 & ~n3060 ) | ( n3055 & ~n3060 ) ;
  assign n3062 = ( x84 & n2875 ) | ( x84 & ~n2937 ) | ( n2875 & ~n2937 ) ;
  assign n3063 = x84 & n2875 ;
  assign n3064 = ( ~n2880 & n3062 ) | ( ~n2880 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3065 = ( n2880 & n3062 ) | ( n2880 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3066 = ( n2880 & n3064 ) | ( n2880 & ~n3065 ) | ( n3064 & ~n3065 ) ;
  assign n3067 = ( x85 & n3061 ) | ( x85 & ~n3066 ) | ( n3061 & ~n3066 ) ;
  assign n3068 = ( x85 & n2881 ) | ( x85 & ~n2937 ) | ( n2881 & ~n2937 ) ;
  assign n3069 = x85 & n2881 ;
  assign n3070 = ( ~n2886 & n3068 ) | ( ~n2886 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3071 = ( n2886 & n3068 ) | ( n2886 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3072 = ( n2886 & n3070 ) | ( n2886 & ~n3071 ) | ( n3070 & ~n3071 ) ;
  assign n3073 = ( x86 & n3067 ) | ( x86 & ~n3072 ) | ( n3067 & ~n3072 ) ;
  assign n3074 = ( x86 & n2887 ) | ( x86 & ~n2937 ) | ( n2887 & ~n2937 ) ;
  assign n3075 = x86 & n2887 ;
  assign n3076 = ( ~n2892 & n3074 ) | ( ~n2892 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = ( n2892 & n3074 ) | ( n2892 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3078 = ( n2892 & n3076 ) | ( n2892 & ~n3077 ) | ( n3076 & ~n3077 ) ;
  assign n3079 = ( x87 & n3073 ) | ( x87 & ~n3078 ) | ( n3073 & ~n3078 ) ;
  assign n3080 = ( x87 & n2893 ) | ( x87 & ~n2937 ) | ( n2893 & ~n2937 ) ;
  assign n3081 = x87 & n2893 ;
  assign n3082 = ( ~n2898 & n3080 ) | ( ~n2898 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3083 = ( n2898 & n3080 ) | ( n2898 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3084 = ( n2898 & n3082 ) | ( n2898 & ~n3083 ) | ( n3082 & ~n3083 ) ;
  assign n3085 = ( x88 & n3079 ) | ( x88 & ~n3084 ) | ( n3079 & ~n3084 ) ;
  assign n3086 = ( x88 & n2899 ) | ( x88 & ~n2937 ) | ( n2899 & ~n2937 ) ;
  assign n3087 = x88 & n2899 ;
  assign n3088 = ( ~n2904 & n3086 ) | ( ~n2904 & n3087 ) | ( n3086 & n3087 ) ;
  assign n3089 = ( n2904 & n3086 ) | ( n2904 & n3087 ) | ( n3086 & n3087 ) ;
  assign n3090 = ( n2904 & n3088 ) | ( n2904 & ~n3089 ) | ( n3088 & ~n3089 ) ;
  assign n3091 = ( x89 & n3085 ) | ( x89 & ~n3090 ) | ( n3085 & ~n3090 ) ;
  assign n3092 = ( x89 & n2905 ) | ( x89 & ~n2937 ) | ( n2905 & ~n2937 ) ;
  assign n3093 = x89 & n2905 ;
  assign n3094 = ( ~n2910 & n3092 ) | ( ~n2910 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3095 = ( n2910 & n3092 ) | ( n2910 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3096 = ( n2910 & n3094 ) | ( n2910 & ~n3095 ) | ( n3094 & ~n3095 ) ;
  assign n3097 = ( x90 & n3091 ) | ( x90 & ~n3096 ) | ( n3091 & ~n3096 ) ;
  assign n3098 = ( x90 & n2911 ) | ( x90 & ~n2937 ) | ( n2911 & ~n2937 ) ;
  assign n3099 = x90 & n2911 ;
  assign n3100 = ( ~n2916 & n3098 ) | ( ~n2916 & n3099 ) | ( n3098 & n3099 ) ;
  assign n3101 = ( n2916 & n3098 ) | ( n2916 & n3099 ) | ( n3098 & n3099 ) ;
  assign n3102 = ( n2916 & n3100 ) | ( n2916 & ~n3101 ) | ( n3100 & ~n3101 ) ;
  assign n3103 = ( x91 & n3097 ) | ( x91 & ~n3102 ) | ( n3097 & ~n3102 ) ;
  assign n3104 = ( x91 & n2917 ) | ( x91 & ~n2937 ) | ( n2917 & ~n2937 ) ;
  assign n3105 = x91 & n2917 ;
  assign n3106 = ( ~n2922 & n3104 ) | ( ~n2922 & n3105 ) | ( n3104 & n3105 ) ;
  assign n3107 = ( n2922 & n3104 ) | ( n2922 & n3105 ) | ( n3104 & n3105 ) ;
  assign n3108 = ( n2922 & n3106 ) | ( n2922 & ~n3107 ) | ( n3106 & ~n3107 ) ;
  assign n3109 = ( x92 & n3103 ) | ( x92 & ~n3108 ) | ( n3103 & ~n3108 ) ;
  assign n3110 = ( x92 & n2923 ) | ( x92 & ~n2937 ) | ( n2923 & ~n2937 ) ;
  assign n3111 = x92 & n2923 ;
  assign n3112 = ( ~n2928 & n3110 ) | ( ~n2928 & n3111 ) | ( n3110 & n3111 ) ;
  assign n3113 = ( n2928 & n3110 ) | ( n2928 & n3111 ) | ( n3110 & n3111 ) ;
  assign n3114 = ( n2928 & n3112 ) | ( n2928 & ~n3113 ) | ( n3112 & ~n3113 ) ;
  assign n3115 = ( x93 & n3109 ) | ( x93 & ~n3114 ) | ( n3109 & ~n3114 ) ;
  assign n3116 = ( x94 & ~n162 ) | ( x94 & n2930 ) | ( ~n162 & n2930 ) ;
  assign n3117 = x94 & n2930 ;
  assign n3118 = ( n2935 & ~n3116 ) | ( n2935 & n3117 ) | ( ~n3116 & n3117 ) ;
  assign n3119 = ( x94 & ~n2942 ) | ( x94 & n3115 ) | ( ~n2942 & n3115 ) ;
  assign n3120 = ( x95 & ~n3118 ) | ( x95 & n3119 ) | ( ~n3118 & n3119 ) ;
  assign n3121 = n161 | n3120 ;
  assign n3122 = ( x94 & n3115 ) | ( x94 & n3121 ) | ( n3115 & n3121 ) ;
  assign n3123 = x94 | n3115 ;
  assign n3124 = ( ~n2942 & n3122 ) | ( ~n2942 & n3123 ) | ( n3122 & n3123 ) ;
  assign n3125 = ( n2942 & n3122 ) | ( n2942 & n3123 ) | ( n3122 & n3123 ) ;
  assign n3126 = ( n2942 & n3124 ) | ( n2942 & ~n3125 ) | ( n3124 & ~n3125 ) ;
  assign n3127 = ~x31 & x64 ;
  assign n3128 = ~x32 & n3121 ;
  assign n3129 = ( x32 & ~x64 ) | ( x32 & n3121 ) | ( ~x64 & n3121 ) ;
  assign n3130 = ( n2943 & ~n3128 ) | ( n2943 & n3129 ) | ( ~n3128 & n3129 ) ;
  assign n3131 = ( x65 & n3127 ) | ( x65 & ~n3130 ) | ( n3127 & ~n3130 ) ;
  assign n3132 = ( x65 & n2943 ) | ( x65 & n3121 ) | ( n2943 & n3121 ) ;
  assign n3133 = x65 | n2943 ;
  assign n3134 = ( ~n2946 & n3132 ) | ( ~n2946 & n3133 ) | ( n3132 & n3133 ) ;
  assign n3135 = ( n2946 & n3132 ) | ( n2946 & n3133 ) | ( n3132 & n3133 ) ;
  assign n3136 = ( n2946 & n3134 ) | ( n2946 & ~n3135 ) | ( n3134 & ~n3135 ) ;
  assign n3137 = ( x66 & n3131 ) | ( x66 & ~n3136 ) | ( n3131 & ~n3136 ) ;
  assign n3138 = ( x66 & n2947 ) | ( x66 & n3121 ) | ( n2947 & n3121 ) ;
  assign n3139 = x66 | n2947 ;
  assign n3140 = ( ~n2952 & n3138 ) | ( ~n2952 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3141 = ( n2952 & n3138 ) | ( n2952 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3142 = ( n2952 & n3140 ) | ( n2952 & ~n3141 ) | ( n3140 & ~n3141 ) ;
  assign n3143 = ( x67 & n3137 ) | ( x67 & ~n3142 ) | ( n3137 & ~n3142 ) ;
  assign n3144 = ( x67 & n2953 ) | ( x67 & ~n3121 ) | ( n2953 & ~n3121 ) ;
  assign n3145 = x67 & n2953 ;
  assign n3146 = ( ~n2958 & n3144 ) | ( ~n2958 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3147 = ( n2958 & n3144 ) | ( n2958 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3148 = ( n2958 & n3146 ) | ( n2958 & ~n3147 ) | ( n3146 & ~n3147 ) ;
  assign n3149 = ( x68 & n3143 ) | ( x68 & ~n3148 ) | ( n3143 & ~n3148 ) ;
  assign n3150 = ( x68 & n2959 ) | ( x68 & ~n3121 ) | ( n2959 & ~n3121 ) ;
  assign n3151 = x68 & n2959 ;
  assign n3152 = ( ~n2964 & n3150 ) | ( ~n2964 & n3151 ) | ( n3150 & n3151 ) ;
  assign n3153 = ( n2964 & n3150 ) | ( n2964 & n3151 ) | ( n3150 & n3151 ) ;
  assign n3154 = ( n2964 & n3152 ) | ( n2964 & ~n3153 ) | ( n3152 & ~n3153 ) ;
  assign n3155 = ( x69 & n3149 ) | ( x69 & ~n3154 ) | ( n3149 & ~n3154 ) ;
  assign n3156 = ( x69 & n2965 ) | ( x69 & ~n3121 ) | ( n2965 & ~n3121 ) ;
  assign n3157 = x69 & n2965 ;
  assign n3158 = ( ~n2970 & n3156 ) | ( ~n2970 & n3157 ) | ( n3156 & n3157 ) ;
  assign n3159 = ( n2970 & n3156 ) | ( n2970 & n3157 ) | ( n3156 & n3157 ) ;
  assign n3160 = ( n2970 & n3158 ) | ( n2970 & ~n3159 ) | ( n3158 & ~n3159 ) ;
  assign n3161 = ( x70 & n3155 ) | ( x70 & ~n3160 ) | ( n3155 & ~n3160 ) ;
  assign n3162 = ( x70 & n2971 ) | ( x70 & ~n3121 ) | ( n2971 & ~n3121 ) ;
  assign n3163 = x70 & n2971 ;
  assign n3164 = ( ~n2976 & n3162 ) | ( ~n2976 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3165 = ( n2976 & n3162 ) | ( n2976 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3166 = ( n2976 & n3164 ) | ( n2976 & ~n3165 ) | ( n3164 & ~n3165 ) ;
  assign n3167 = ( x71 & n3161 ) | ( x71 & ~n3166 ) | ( n3161 & ~n3166 ) ;
  assign n3168 = ( x71 & n2977 ) | ( x71 & ~n3121 ) | ( n2977 & ~n3121 ) ;
  assign n3169 = x71 & n2977 ;
  assign n3170 = ( ~n2982 & n3168 ) | ( ~n2982 & n3169 ) | ( n3168 & n3169 ) ;
  assign n3171 = ( n2982 & n3168 ) | ( n2982 & n3169 ) | ( n3168 & n3169 ) ;
  assign n3172 = ( n2982 & n3170 ) | ( n2982 & ~n3171 ) | ( n3170 & ~n3171 ) ;
  assign n3173 = ( x72 & n3167 ) | ( x72 & ~n3172 ) | ( n3167 & ~n3172 ) ;
  assign n3174 = ( x72 & n2983 ) | ( x72 & ~n3121 ) | ( n2983 & ~n3121 ) ;
  assign n3175 = x72 & n2983 ;
  assign n3176 = ( ~n2988 & n3174 ) | ( ~n2988 & n3175 ) | ( n3174 & n3175 ) ;
  assign n3177 = ( n2988 & n3174 ) | ( n2988 & n3175 ) | ( n3174 & n3175 ) ;
  assign n3178 = ( n2988 & n3176 ) | ( n2988 & ~n3177 ) | ( n3176 & ~n3177 ) ;
  assign n3179 = ( x73 & n3173 ) | ( x73 & ~n3178 ) | ( n3173 & ~n3178 ) ;
  assign n3180 = ( x73 & n2989 ) | ( x73 & ~n3121 ) | ( n2989 & ~n3121 ) ;
  assign n3181 = x73 & n2989 ;
  assign n3182 = ( ~n2994 & n3180 ) | ( ~n2994 & n3181 ) | ( n3180 & n3181 ) ;
  assign n3183 = ( n2994 & n3180 ) | ( n2994 & n3181 ) | ( n3180 & n3181 ) ;
  assign n3184 = ( n2994 & n3182 ) | ( n2994 & ~n3183 ) | ( n3182 & ~n3183 ) ;
  assign n3185 = ( x74 & n3179 ) | ( x74 & ~n3184 ) | ( n3179 & ~n3184 ) ;
  assign n3186 = ( x74 & n2995 ) | ( x74 & ~n3121 ) | ( n2995 & ~n3121 ) ;
  assign n3187 = x74 & n2995 ;
  assign n3188 = ( ~n3000 & n3186 ) | ( ~n3000 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3189 = ( n3000 & n3186 ) | ( n3000 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3190 = ( n3000 & n3188 ) | ( n3000 & ~n3189 ) | ( n3188 & ~n3189 ) ;
  assign n3191 = ( x75 & n3185 ) | ( x75 & ~n3190 ) | ( n3185 & ~n3190 ) ;
  assign n3192 = ( x75 & n3001 ) | ( x75 & ~n3121 ) | ( n3001 & ~n3121 ) ;
  assign n3193 = x75 & n3001 ;
  assign n3194 = ( ~n3006 & n3192 ) | ( ~n3006 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3195 = ( n3006 & n3192 ) | ( n3006 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3196 = ( n3006 & n3194 ) | ( n3006 & ~n3195 ) | ( n3194 & ~n3195 ) ;
  assign n3197 = ( x76 & n3191 ) | ( x76 & ~n3196 ) | ( n3191 & ~n3196 ) ;
  assign n3198 = ( x76 & n3007 ) | ( x76 & ~n3121 ) | ( n3007 & ~n3121 ) ;
  assign n3199 = x76 & n3007 ;
  assign n3200 = ( ~n3012 & n3198 ) | ( ~n3012 & n3199 ) | ( n3198 & n3199 ) ;
  assign n3201 = ( n3012 & n3198 ) | ( n3012 & n3199 ) | ( n3198 & n3199 ) ;
  assign n3202 = ( n3012 & n3200 ) | ( n3012 & ~n3201 ) | ( n3200 & ~n3201 ) ;
  assign n3203 = ( x77 & n3197 ) | ( x77 & ~n3202 ) | ( n3197 & ~n3202 ) ;
  assign n3204 = ( x77 & n3013 ) | ( x77 & ~n3121 ) | ( n3013 & ~n3121 ) ;
  assign n3205 = x77 & n3013 ;
  assign n3206 = ( ~n3018 & n3204 ) | ( ~n3018 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3207 = ( n3018 & n3204 ) | ( n3018 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3208 = ( n3018 & n3206 ) | ( n3018 & ~n3207 ) | ( n3206 & ~n3207 ) ;
  assign n3209 = ( x78 & n3203 ) | ( x78 & ~n3208 ) | ( n3203 & ~n3208 ) ;
  assign n3210 = ( x78 & n3019 ) | ( x78 & ~n3121 ) | ( n3019 & ~n3121 ) ;
  assign n3211 = x78 & n3019 ;
  assign n3212 = ( ~n3024 & n3210 ) | ( ~n3024 & n3211 ) | ( n3210 & n3211 ) ;
  assign n3213 = ( n3024 & n3210 ) | ( n3024 & n3211 ) | ( n3210 & n3211 ) ;
  assign n3214 = ( n3024 & n3212 ) | ( n3024 & ~n3213 ) | ( n3212 & ~n3213 ) ;
  assign n3215 = ( x79 & n3209 ) | ( x79 & ~n3214 ) | ( n3209 & ~n3214 ) ;
  assign n3216 = ( x79 & n3025 ) | ( x79 & ~n3121 ) | ( n3025 & ~n3121 ) ;
  assign n3217 = x79 & n3025 ;
  assign n3218 = ( ~n3030 & n3216 ) | ( ~n3030 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3219 = ( n3030 & n3216 ) | ( n3030 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3220 = ( n3030 & n3218 ) | ( n3030 & ~n3219 ) | ( n3218 & ~n3219 ) ;
  assign n3221 = ( x80 & n3215 ) | ( x80 & ~n3220 ) | ( n3215 & ~n3220 ) ;
  assign n3222 = ( x80 & n3031 ) | ( x80 & ~n3121 ) | ( n3031 & ~n3121 ) ;
  assign n3223 = x80 & n3031 ;
  assign n3224 = ( ~n3036 & n3222 ) | ( ~n3036 & n3223 ) | ( n3222 & n3223 ) ;
  assign n3225 = ( n3036 & n3222 ) | ( n3036 & n3223 ) | ( n3222 & n3223 ) ;
  assign n3226 = ( n3036 & n3224 ) | ( n3036 & ~n3225 ) | ( n3224 & ~n3225 ) ;
  assign n3227 = ( x81 & n3221 ) | ( x81 & ~n3226 ) | ( n3221 & ~n3226 ) ;
  assign n3228 = ( x81 & n3037 ) | ( x81 & ~n3121 ) | ( n3037 & ~n3121 ) ;
  assign n3229 = x81 & n3037 ;
  assign n3230 = ( ~n3042 & n3228 ) | ( ~n3042 & n3229 ) | ( n3228 & n3229 ) ;
  assign n3231 = ( n3042 & n3228 ) | ( n3042 & n3229 ) | ( n3228 & n3229 ) ;
  assign n3232 = ( n3042 & n3230 ) | ( n3042 & ~n3231 ) | ( n3230 & ~n3231 ) ;
  assign n3233 = ( x82 & n3227 ) | ( x82 & ~n3232 ) | ( n3227 & ~n3232 ) ;
  assign n3234 = ( x82 & n3043 ) | ( x82 & ~n3121 ) | ( n3043 & ~n3121 ) ;
  assign n3235 = x82 & n3043 ;
  assign n3236 = ( ~n3048 & n3234 ) | ( ~n3048 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3237 = ( n3048 & n3234 ) | ( n3048 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3238 = ( n3048 & n3236 ) | ( n3048 & ~n3237 ) | ( n3236 & ~n3237 ) ;
  assign n3239 = ( x83 & n3233 ) | ( x83 & ~n3238 ) | ( n3233 & ~n3238 ) ;
  assign n3240 = ( x83 & n3049 ) | ( x83 & ~n3121 ) | ( n3049 & ~n3121 ) ;
  assign n3241 = x83 & n3049 ;
  assign n3242 = ( ~n3054 & n3240 ) | ( ~n3054 & n3241 ) | ( n3240 & n3241 ) ;
  assign n3243 = ( n3054 & n3240 ) | ( n3054 & n3241 ) | ( n3240 & n3241 ) ;
  assign n3244 = ( n3054 & n3242 ) | ( n3054 & ~n3243 ) | ( n3242 & ~n3243 ) ;
  assign n3245 = ( x84 & n3239 ) | ( x84 & ~n3244 ) | ( n3239 & ~n3244 ) ;
  assign n3246 = ( x84 & n3055 ) | ( x84 & ~n3121 ) | ( n3055 & ~n3121 ) ;
  assign n3247 = x84 & n3055 ;
  assign n3248 = ( ~n3060 & n3246 ) | ( ~n3060 & n3247 ) | ( n3246 & n3247 ) ;
  assign n3249 = ( n3060 & n3246 ) | ( n3060 & n3247 ) | ( n3246 & n3247 ) ;
  assign n3250 = ( n3060 & n3248 ) | ( n3060 & ~n3249 ) | ( n3248 & ~n3249 ) ;
  assign n3251 = ( x85 & n3245 ) | ( x85 & ~n3250 ) | ( n3245 & ~n3250 ) ;
  assign n3252 = ( x85 & n3061 ) | ( x85 & ~n3121 ) | ( n3061 & ~n3121 ) ;
  assign n3253 = x85 & n3061 ;
  assign n3254 = ( ~n3066 & n3252 ) | ( ~n3066 & n3253 ) | ( n3252 & n3253 ) ;
  assign n3255 = ( n3066 & n3252 ) | ( n3066 & n3253 ) | ( n3252 & n3253 ) ;
  assign n3256 = ( n3066 & n3254 ) | ( n3066 & ~n3255 ) | ( n3254 & ~n3255 ) ;
  assign n3257 = ( x86 & n3251 ) | ( x86 & ~n3256 ) | ( n3251 & ~n3256 ) ;
  assign n3258 = ( x86 & n3067 ) | ( x86 & ~n3121 ) | ( n3067 & ~n3121 ) ;
  assign n3259 = x86 & n3067 ;
  assign n3260 = ( ~n3072 & n3258 ) | ( ~n3072 & n3259 ) | ( n3258 & n3259 ) ;
  assign n3261 = ( n3072 & n3258 ) | ( n3072 & n3259 ) | ( n3258 & n3259 ) ;
  assign n3262 = ( n3072 & n3260 ) | ( n3072 & ~n3261 ) | ( n3260 & ~n3261 ) ;
  assign n3263 = ( x87 & n3257 ) | ( x87 & ~n3262 ) | ( n3257 & ~n3262 ) ;
  assign n3264 = ( x87 & n3073 ) | ( x87 & ~n3121 ) | ( n3073 & ~n3121 ) ;
  assign n3265 = x87 & n3073 ;
  assign n3266 = ( ~n3078 & n3264 ) | ( ~n3078 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3267 = ( n3078 & n3264 ) | ( n3078 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3268 = ( n3078 & n3266 ) | ( n3078 & ~n3267 ) | ( n3266 & ~n3267 ) ;
  assign n3269 = ( x88 & n3263 ) | ( x88 & ~n3268 ) | ( n3263 & ~n3268 ) ;
  assign n3270 = ( x88 & n3079 ) | ( x88 & ~n3121 ) | ( n3079 & ~n3121 ) ;
  assign n3271 = x88 & n3079 ;
  assign n3272 = ( ~n3084 & n3270 ) | ( ~n3084 & n3271 ) | ( n3270 & n3271 ) ;
  assign n3273 = ( n3084 & n3270 ) | ( n3084 & n3271 ) | ( n3270 & n3271 ) ;
  assign n3274 = ( n3084 & n3272 ) | ( n3084 & ~n3273 ) | ( n3272 & ~n3273 ) ;
  assign n3275 = ( x89 & n3269 ) | ( x89 & ~n3274 ) | ( n3269 & ~n3274 ) ;
  assign n3276 = ( x89 & n3085 ) | ( x89 & ~n3121 ) | ( n3085 & ~n3121 ) ;
  assign n3277 = x89 & n3085 ;
  assign n3278 = ( ~n3090 & n3276 ) | ( ~n3090 & n3277 ) | ( n3276 & n3277 ) ;
  assign n3279 = ( n3090 & n3276 ) | ( n3090 & n3277 ) | ( n3276 & n3277 ) ;
  assign n3280 = ( n3090 & n3278 ) | ( n3090 & ~n3279 ) | ( n3278 & ~n3279 ) ;
  assign n3281 = ( x90 & n3275 ) | ( x90 & ~n3280 ) | ( n3275 & ~n3280 ) ;
  assign n3282 = ( x90 & n3091 ) | ( x90 & ~n3121 ) | ( n3091 & ~n3121 ) ;
  assign n3283 = x90 & n3091 ;
  assign n3284 = ( ~n3096 & n3282 ) | ( ~n3096 & n3283 ) | ( n3282 & n3283 ) ;
  assign n3285 = ( n3096 & n3282 ) | ( n3096 & n3283 ) | ( n3282 & n3283 ) ;
  assign n3286 = ( n3096 & n3284 ) | ( n3096 & ~n3285 ) | ( n3284 & ~n3285 ) ;
  assign n3287 = ( x91 & n3281 ) | ( x91 & ~n3286 ) | ( n3281 & ~n3286 ) ;
  assign n3288 = ( x91 & n3097 ) | ( x91 & ~n3121 ) | ( n3097 & ~n3121 ) ;
  assign n3289 = x91 & n3097 ;
  assign n3290 = ( ~n3102 & n3288 ) | ( ~n3102 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = ( n3102 & n3288 ) | ( n3102 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3292 = ( n3102 & n3290 ) | ( n3102 & ~n3291 ) | ( n3290 & ~n3291 ) ;
  assign n3293 = ( x92 & n3287 ) | ( x92 & ~n3292 ) | ( n3287 & ~n3292 ) ;
  assign n3294 = ( x92 & n3103 ) | ( x92 & ~n3121 ) | ( n3103 & ~n3121 ) ;
  assign n3295 = x92 & n3103 ;
  assign n3296 = ( ~n3108 & n3294 ) | ( ~n3108 & n3295 ) | ( n3294 & n3295 ) ;
  assign n3297 = ( n3108 & n3294 ) | ( n3108 & n3295 ) | ( n3294 & n3295 ) ;
  assign n3298 = ( n3108 & n3296 ) | ( n3108 & ~n3297 ) | ( n3296 & ~n3297 ) ;
  assign n3299 = ( x93 & n3293 ) | ( x93 & ~n3298 ) | ( n3293 & ~n3298 ) ;
  assign n3300 = ( x93 & n3109 ) | ( x93 & ~n3121 ) | ( n3109 & ~n3121 ) ;
  assign n3301 = x93 & n3109 ;
  assign n3302 = ( ~n3114 & n3300 ) | ( ~n3114 & n3301 ) | ( n3300 & n3301 ) ;
  assign n3303 = ( n3114 & n3300 ) | ( n3114 & n3301 ) | ( n3300 & n3301 ) ;
  assign n3304 = ( n3114 & n3302 ) | ( n3114 & ~n3303 ) | ( n3302 & ~n3303 ) ;
  assign n3305 = ( x94 & n3299 ) | ( x94 & ~n3304 ) | ( n3299 & ~n3304 ) ;
  assign n3306 = ( n160 & n161 ) | ( n160 & ~n3118 ) | ( n161 & ~n3118 ) ;
  assign n3307 = ( x95 & ~n3126 ) | ( x95 & n3305 ) | ( ~n3126 & n3305 ) ;
  assign n3308 = n3306 | n3307 ;
  assign n3309 = ( ~x95 & n161 ) | ( ~x95 & n3119 ) | ( n161 & n3119 ) ;
  assign n3310 = ( ~x95 & n3118 ) | ( ~x95 & n3119 ) | ( n3118 & n3119 ) ;
  assign n3311 = ~n3309 & n3310 ;
  assign n3312 = n3308 & ~n3311 ;
  assign n3313 = ( x95 & n3305 ) | ( x95 & ~n3312 ) | ( n3305 & ~n3312 ) ;
  assign n3314 = x95 & n3305 ;
  assign n3315 = ( ~n3126 & n3313 ) | ( ~n3126 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3316 = ( n3126 & n3313 ) | ( n3126 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3317 = ( n3126 & n3315 ) | ( n3126 & ~n3316 ) | ( n3315 & ~n3316 ) ;
  assign n3318 = ~x30 & x64 ;
  assign n3319 = x31 & n3312 ;
  assign n3320 = ( x31 & x64 ) | ( x31 & ~n3312 ) | ( x64 & ~n3312 ) ;
  assign n3321 = x31 & x64 ;
  assign n3322 = ( n3319 & n3320 ) | ( n3319 & ~n3321 ) | ( n3320 & ~n3321 ) ;
  assign n3323 = ( x65 & n3318 ) | ( x65 & ~n3322 ) | ( n3318 & ~n3322 ) ;
  assign n3324 = ( x65 & n3127 ) | ( x65 & n3312 ) | ( n3127 & n3312 ) ;
  assign n3325 = x65 | n3127 ;
  assign n3326 = ( ~n3130 & n3324 ) | ( ~n3130 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3327 = ( n3130 & n3324 ) | ( n3130 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3328 = ( n3130 & n3326 ) | ( n3130 & ~n3327 ) | ( n3326 & ~n3327 ) ;
  assign n3329 = ( x66 & n3323 ) | ( x66 & ~n3328 ) | ( n3323 & ~n3328 ) ;
  assign n3330 = ( x66 & n3131 ) | ( x66 & n3312 ) | ( n3131 & n3312 ) ;
  assign n3331 = x66 | n3131 ;
  assign n3332 = ( ~n3136 & n3330 ) | ( ~n3136 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3333 = ( n3136 & n3330 ) | ( n3136 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3334 = ( n3136 & n3332 ) | ( n3136 & ~n3333 ) | ( n3332 & ~n3333 ) ;
  assign n3335 = ( x67 & n3329 ) | ( x67 & ~n3334 ) | ( n3329 & ~n3334 ) ;
  assign n3336 = ( x67 & n3137 ) | ( x67 & ~n3312 ) | ( n3137 & ~n3312 ) ;
  assign n3337 = x67 & n3137 ;
  assign n3338 = ( ~n3142 & n3336 ) | ( ~n3142 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3339 = ( n3142 & n3336 ) | ( n3142 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3340 = ( n3142 & n3338 ) | ( n3142 & ~n3339 ) | ( n3338 & ~n3339 ) ;
  assign n3341 = ( x68 & n3335 ) | ( x68 & ~n3340 ) | ( n3335 & ~n3340 ) ;
  assign n3342 = ( x68 & n3143 ) | ( x68 & ~n3312 ) | ( n3143 & ~n3312 ) ;
  assign n3343 = x68 & n3143 ;
  assign n3344 = ( ~n3148 & n3342 ) | ( ~n3148 & n3343 ) | ( n3342 & n3343 ) ;
  assign n3345 = ( n3148 & n3342 ) | ( n3148 & n3343 ) | ( n3342 & n3343 ) ;
  assign n3346 = ( n3148 & n3344 ) | ( n3148 & ~n3345 ) | ( n3344 & ~n3345 ) ;
  assign n3347 = ( x69 & n3341 ) | ( x69 & ~n3346 ) | ( n3341 & ~n3346 ) ;
  assign n3348 = ( x69 & n3149 ) | ( x69 & ~n3312 ) | ( n3149 & ~n3312 ) ;
  assign n3349 = x69 & n3149 ;
  assign n3350 = ( ~n3154 & n3348 ) | ( ~n3154 & n3349 ) | ( n3348 & n3349 ) ;
  assign n3351 = ( n3154 & n3348 ) | ( n3154 & n3349 ) | ( n3348 & n3349 ) ;
  assign n3352 = ( n3154 & n3350 ) | ( n3154 & ~n3351 ) | ( n3350 & ~n3351 ) ;
  assign n3353 = ( x70 & n3347 ) | ( x70 & ~n3352 ) | ( n3347 & ~n3352 ) ;
  assign n3354 = ( x70 & n3155 ) | ( x70 & ~n3312 ) | ( n3155 & ~n3312 ) ;
  assign n3355 = x70 & n3155 ;
  assign n3356 = ( ~n3160 & n3354 ) | ( ~n3160 & n3355 ) | ( n3354 & n3355 ) ;
  assign n3357 = ( n3160 & n3354 ) | ( n3160 & n3355 ) | ( n3354 & n3355 ) ;
  assign n3358 = ( n3160 & n3356 ) | ( n3160 & ~n3357 ) | ( n3356 & ~n3357 ) ;
  assign n3359 = ( x71 & n3353 ) | ( x71 & ~n3358 ) | ( n3353 & ~n3358 ) ;
  assign n3360 = ( x71 & n3161 ) | ( x71 & ~n3312 ) | ( n3161 & ~n3312 ) ;
  assign n3361 = x71 & n3161 ;
  assign n3362 = ( ~n3166 & n3360 ) | ( ~n3166 & n3361 ) | ( n3360 & n3361 ) ;
  assign n3363 = ( n3166 & n3360 ) | ( n3166 & n3361 ) | ( n3360 & n3361 ) ;
  assign n3364 = ( n3166 & n3362 ) | ( n3166 & ~n3363 ) | ( n3362 & ~n3363 ) ;
  assign n3365 = ( x72 & n3359 ) | ( x72 & ~n3364 ) | ( n3359 & ~n3364 ) ;
  assign n3366 = ( x72 & n3167 ) | ( x72 & ~n3312 ) | ( n3167 & ~n3312 ) ;
  assign n3367 = x72 & n3167 ;
  assign n3368 = ( ~n3172 & n3366 ) | ( ~n3172 & n3367 ) | ( n3366 & n3367 ) ;
  assign n3369 = ( n3172 & n3366 ) | ( n3172 & n3367 ) | ( n3366 & n3367 ) ;
  assign n3370 = ( n3172 & n3368 ) | ( n3172 & ~n3369 ) | ( n3368 & ~n3369 ) ;
  assign n3371 = ( x73 & n3365 ) | ( x73 & ~n3370 ) | ( n3365 & ~n3370 ) ;
  assign n3372 = ( x73 & n3173 ) | ( x73 & ~n3312 ) | ( n3173 & ~n3312 ) ;
  assign n3373 = x73 & n3173 ;
  assign n3374 = ( ~n3178 & n3372 ) | ( ~n3178 & n3373 ) | ( n3372 & n3373 ) ;
  assign n3375 = ( n3178 & n3372 ) | ( n3178 & n3373 ) | ( n3372 & n3373 ) ;
  assign n3376 = ( n3178 & n3374 ) | ( n3178 & ~n3375 ) | ( n3374 & ~n3375 ) ;
  assign n3377 = ( x74 & n3371 ) | ( x74 & ~n3376 ) | ( n3371 & ~n3376 ) ;
  assign n3378 = ( x74 & n3179 ) | ( x74 & ~n3312 ) | ( n3179 & ~n3312 ) ;
  assign n3379 = x74 & n3179 ;
  assign n3380 = ( ~n3184 & n3378 ) | ( ~n3184 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = ( n3184 & n3378 ) | ( n3184 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3382 = ( n3184 & n3380 ) | ( n3184 & ~n3381 ) | ( n3380 & ~n3381 ) ;
  assign n3383 = ( x75 & n3377 ) | ( x75 & ~n3382 ) | ( n3377 & ~n3382 ) ;
  assign n3384 = ( x75 & n3185 ) | ( x75 & ~n3312 ) | ( n3185 & ~n3312 ) ;
  assign n3385 = x75 & n3185 ;
  assign n3386 = ( ~n3190 & n3384 ) | ( ~n3190 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3387 = ( n3190 & n3384 ) | ( n3190 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3388 = ( n3190 & n3386 ) | ( n3190 & ~n3387 ) | ( n3386 & ~n3387 ) ;
  assign n3389 = ( x76 & n3383 ) | ( x76 & ~n3388 ) | ( n3383 & ~n3388 ) ;
  assign n3390 = ( x76 & n3191 ) | ( x76 & ~n3312 ) | ( n3191 & ~n3312 ) ;
  assign n3391 = x76 & n3191 ;
  assign n3392 = ( ~n3196 & n3390 ) | ( ~n3196 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = ( n3196 & n3390 ) | ( n3196 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3394 = ( n3196 & n3392 ) | ( n3196 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = ( x77 & n3389 ) | ( x77 & ~n3394 ) | ( n3389 & ~n3394 ) ;
  assign n3396 = ( x77 & n3197 ) | ( x77 & ~n3312 ) | ( n3197 & ~n3312 ) ;
  assign n3397 = x77 & n3197 ;
  assign n3398 = ( ~n3202 & n3396 ) | ( ~n3202 & n3397 ) | ( n3396 & n3397 ) ;
  assign n3399 = ( n3202 & n3396 ) | ( n3202 & n3397 ) | ( n3396 & n3397 ) ;
  assign n3400 = ( n3202 & n3398 ) | ( n3202 & ~n3399 ) | ( n3398 & ~n3399 ) ;
  assign n3401 = ( x78 & n3395 ) | ( x78 & ~n3400 ) | ( n3395 & ~n3400 ) ;
  assign n3402 = ( x78 & n3203 ) | ( x78 & ~n3312 ) | ( n3203 & ~n3312 ) ;
  assign n3403 = x78 & n3203 ;
  assign n3404 = ( ~n3208 & n3402 ) | ( ~n3208 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3405 = ( n3208 & n3402 ) | ( n3208 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3406 = ( n3208 & n3404 ) | ( n3208 & ~n3405 ) | ( n3404 & ~n3405 ) ;
  assign n3407 = ( x79 & n3401 ) | ( x79 & ~n3406 ) | ( n3401 & ~n3406 ) ;
  assign n3408 = ( x79 & n3209 ) | ( x79 & ~n3312 ) | ( n3209 & ~n3312 ) ;
  assign n3409 = x79 & n3209 ;
  assign n3410 = ( ~n3214 & n3408 ) | ( ~n3214 & n3409 ) | ( n3408 & n3409 ) ;
  assign n3411 = ( n3214 & n3408 ) | ( n3214 & n3409 ) | ( n3408 & n3409 ) ;
  assign n3412 = ( n3214 & n3410 ) | ( n3214 & ~n3411 ) | ( n3410 & ~n3411 ) ;
  assign n3413 = ( x80 & n3407 ) | ( x80 & ~n3412 ) | ( n3407 & ~n3412 ) ;
  assign n3414 = ( x80 & n3215 ) | ( x80 & ~n3312 ) | ( n3215 & ~n3312 ) ;
  assign n3415 = x80 & n3215 ;
  assign n3416 = ( ~n3220 & n3414 ) | ( ~n3220 & n3415 ) | ( n3414 & n3415 ) ;
  assign n3417 = ( n3220 & n3414 ) | ( n3220 & n3415 ) | ( n3414 & n3415 ) ;
  assign n3418 = ( n3220 & n3416 ) | ( n3220 & ~n3417 ) | ( n3416 & ~n3417 ) ;
  assign n3419 = ( x81 & n3413 ) | ( x81 & ~n3418 ) | ( n3413 & ~n3418 ) ;
  assign n3420 = ( x81 & n3221 ) | ( x81 & ~n3312 ) | ( n3221 & ~n3312 ) ;
  assign n3421 = x81 & n3221 ;
  assign n3422 = ( ~n3226 & n3420 ) | ( ~n3226 & n3421 ) | ( n3420 & n3421 ) ;
  assign n3423 = ( n3226 & n3420 ) | ( n3226 & n3421 ) | ( n3420 & n3421 ) ;
  assign n3424 = ( n3226 & n3422 ) | ( n3226 & ~n3423 ) | ( n3422 & ~n3423 ) ;
  assign n3425 = ( x82 & n3419 ) | ( x82 & ~n3424 ) | ( n3419 & ~n3424 ) ;
  assign n3426 = ( x82 & n3227 ) | ( x82 & ~n3312 ) | ( n3227 & ~n3312 ) ;
  assign n3427 = x82 & n3227 ;
  assign n3428 = ( ~n3232 & n3426 ) | ( ~n3232 & n3427 ) | ( n3426 & n3427 ) ;
  assign n3429 = ( n3232 & n3426 ) | ( n3232 & n3427 ) | ( n3426 & n3427 ) ;
  assign n3430 = ( n3232 & n3428 ) | ( n3232 & ~n3429 ) | ( n3428 & ~n3429 ) ;
  assign n3431 = ( x83 & n3425 ) | ( x83 & ~n3430 ) | ( n3425 & ~n3430 ) ;
  assign n3432 = ( x83 & n3233 ) | ( x83 & ~n3312 ) | ( n3233 & ~n3312 ) ;
  assign n3433 = x83 & n3233 ;
  assign n3434 = ( ~n3238 & n3432 ) | ( ~n3238 & n3433 ) | ( n3432 & n3433 ) ;
  assign n3435 = ( n3238 & n3432 ) | ( n3238 & n3433 ) | ( n3432 & n3433 ) ;
  assign n3436 = ( n3238 & n3434 ) | ( n3238 & ~n3435 ) | ( n3434 & ~n3435 ) ;
  assign n3437 = ( x84 & n3431 ) | ( x84 & ~n3436 ) | ( n3431 & ~n3436 ) ;
  assign n3438 = ( x84 & n3239 ) | ( x84 & ~n3312 ) | ( n3239 & ~n3312 ) ;
  assign n3439 = x84 & n3239 ;
  assign n3440 = ( ~n3244 & n3438 ) | ( ~n3244 & n3439 ) | ( n3438 & n3439 ) ;
  assign n3441 = ( n3244 & n3438 ) | ( n3244 & n3439 ) | ( n3438 & n3439 ) ;
  assign n3442 = ( n3244 & n3440 ) | ( n3244 & ~n3441 ) | ( n3440 & ~n3441 ) ;
  assign n3443 = ( x85 & n3437 ) | ( x85 & ~n3442 ) | ( n3437 & ~n3442 ) ;
  assign n3444 = ( x85 & n3245 ) | ( x85 & ~n3312 ) | ( n3245 & ~n3312 ) ;
  assign n3445 = x85 & n3245 ;
  assign n3446 = ( ~n3250 & n3444 ) | ( ~n3250 & n3445 ) | ( n3444 & n3445 ) ;
  assign n3447 = ( n3250 & n3444 ) | ( n3250 & n3445 ) | ( n3444 & n3445 ) ;
  assign n3448 = ( n3250 & n3446 ) | ( n3250 & ~n3447 ) | ( n3446 & ~n3447 ) ;
  assign n3449 = ( x86 & n3443 ) | ( x86 & ~n3448 ) | ( n3443 & ~n3448 ) ;
  assign n3450 = ( x86 & n3251 ) | ( x86 & ~n3312 ) | ( n3251 & ~n3312 ) ;
  assign n3451 = x86 & n3251 ;
  assign n3452 = ( ~n3256 & n3450 ) | ( ~n3256 & n3451 ) | ( n3450 & n3451 ) ;
  assign n3453 = ( n3256 & n3450 ) | ( n3256 & n3451 ) | ( n3450 & n3451 ) ;
  assign n3454 = ( n3256 & n3452 ) | ( n3256 & ~n3453 ) | ( n3452 & ~n3453 ) ;
  assign n3455 = ( x87 & n3449 ) | ( x87 & ~n3454 ) | ( n3449 & ~n3454 ) ;
  assign n3456 = ( x87 & n3257 ) | ( x87 & ~n3312 ) | ( n3257 & ~n3312 ) ;
  assign n3457 = x87 & n3257 ;
  assign n3458 = ( ~n3262 & n3456 ) | ( ~n3262 & n3457 ) | ( n3456 & n3457 ) ;
  assign n3459 = ( n3262 & n3456 ) | ( n3262 & n3457 ) | ( n3456 & n3457 ) ;
  assign n3460 = ( n3262 & n3458 ) | ( n3262 & ~n3459 ) | ( n3458 & ~n3459 ) ;
  assign n3461 = ( x88 & n3455 ) | ( x88 & ~n3460 ) | ( n3455 & ~n3460 ) ;
  assign n3462 = ( x88 & n3263 ) | ( x88 & ~n3312 ) | ( n3263 & ~n3312 ) ;
  assign n3463 = x88 & n3263 ;
  assign n3464 = ( ~n3268 & n3462 ) | ( ~n3268 & n3463 ) | ( n3462 & n3463 ) ;
  assign n3465 = ( n3268 & n3462 ) | ( n3268 & n3463 ) | ( n3462 & n3463 ) ;
  assign n3466 = ( n3268 & n3464 ) | ( n3268 & ~n3465 ) | ( n3464 & ~n3465 ) ;
  assign n3467 = ( x89 & n3461 ) | ( x89 & ~n3466 ) | ( n3461 & ~n3466 ) ;
  assign n3468 = ( x89 & n3269 ) | ( x89 & ~n3312 ) | ( n3269 & ~n3312 ) ;
  assign n3469 = x89 & n3269 ;
  assign n3470 = ( ~n3274 & n3468 ) | ( ~n3274 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = ( n3274 & n3468 ) | ( n3274 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3472 = ( n3274 & n3470 ) | ( n3274 & ~n3471 ) | ( n3470 & ~n3471 ) ;
  assign n3473 = ( x90 & n3467 ) | ( x90 & ~n3472 ) | ( n3467 & ~n3472 ) ;
  assign n3474 = ( x90 & n3275 ) | ( x90 & ~n3312 ) | ( n3275 & ~n3312 ) ;
  assign n3475 = x90 & n3275 ;
  assign n3476 = ( ~n3280 & n3474 ) | ( ~n3280 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3477 = ( n3280 & n3474 ) | ( n3280 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3478 = ( n3280 & n3476 ) | ( n3280 & ~n3477 ) | ( n3476 & ~n3477 ) ;
  assign n3479 = ( x91 & n3473 ) | ( x91 & ~n3478 ) | ( n3473 & ~n3478 ) ;
  assign n3480 = ( x91 & n3281 ) | ( x91 & ~n3312 ) | ( n3281 & ~n3312 ) ;
  assign n3481 = x91 & n3281 ;
  assign n3482 = ( ~n3286 & n3480 ) | ( ~n3286 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3483 = ( n3286 & n3480 ) | ( n3286 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3484 = ( n3286 & n3482 ) | ( n3286 & ~n3483 ) | ( n3482 & ~n3483 ) ;
  assign n3485 = ( x92 & n3479 ) | ( x92 & ~n3484 ) | ( n3479 & ~n3484 ) ;
  assign n3486 = ( x92 & n3287 ) | ( x92 & ~n3312 ) | ( n3287 & ~n3312 ) ;
  assign n3487 = x92 & n3287 ;
  assign n3488 = ( ~n3292 & n3486 ) | ( ~n3292 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = ( n3292 & n3486 ) | ( n3292 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3490 = ( n3292 & n3488 ) | ( n3292 & ~n3489 ) | ( n3488 & ~n3489 ) ;
  assign n3491 = ( x93 & n3485 ) | ( x93 & ~n3490 ) | ( n3485 & ~n3490 ) ;
  assign n3492 = ( x93 & n3293 ) | ( x93 & ~n3312 ) | ( n3293 & ~n3312 ) ;
  assign n3493 = x93 & n3293 ;
  assign n3494 = ( ~n3298 & n3492 ) | ( ~n3298 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3495 = ( n3298 & n3492 ) | ( n3298 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3496 = ( n3298 & n3494 ) | ( n3298 & ~n3495 ) | ( n3494 & ~n3495 ) ;
  assign n3497 = ( x94 & n3491 ) | ( x94 & ~n3496 ) | ( n3491 & ~n3496 ) ;
  assign n3498 = ( x94 & n3299 ) | ( x94 & ~n3312 ) | ( n3299 & ~n3312 ) ;
  assign n3499 = x94 & n3299 ;
  assign n3500 = ( ~n3304 & n3498 ) | ( ~n3304 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = ( n3304 & n3498 ) | ( n3304 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3502 = ( n3304 & n3500 ) | ( n3304 & ~n3501 ) | ( n3500 & ~n3501 ) ;
  assign n3503 = ( x95 & n3497 ) | ( x95 & ~n3502 ) | ( n3497 & ~n3502 ) ;
  assign n3504 = ( x96 & ~n3317 ) | ( x96 & n3503 ) | ( ~n3317 & n3503 ) ;
  assign n3505 = n161 & n2935 ;
  assign n3506 = n3308 & n3505 ;
  assign n3507 = n389 | n3506 ;
  assign n3508 = ( x97 & n3504 ) | ( x97 & ~n3507 ) | ( n3504 & ~n3507 ) ;
  assign n3509 = n159 | n3508 ;
  assign n3510 = ( x96 & n3503 ) | ( x96 & n3509 ) | ( n3503 & n3509 ) ;
  assign n3511 = x96 | n3503 ;
  assign n3512 = ( ~n3317 & n3510 ) | ( ~n3317 & n3511 ) | ( n3510 & n3511 ) ;
  assign n3513 = ( n3317 & n3510 ) | ( n3317 & n3511 ) | ( n3510 & n3511 ) ;
  assign n3514 = ( n3317 & n3512 ) | ( n3317 & ~n3513 ) | ( n3512 & ~n3513 ) ;
  assign n3515 = ~x29 & x64 ;
  assign n3516 = ~x30 & n3509 ;
  assign n3517 = ( x30 & ~x64 ) | ( x30 & n3509 ) | ( ~x64 & n3509 ) ;
  assign n3518 = ( n3318 & ~n3516 ) | ( n3318 & n3517 ) | ( ~n3516 & n3517 ) ;
  assign n3519 = ( x65 & n3515 ) | ( x65 & ~n3518 ) | ( n3515 & ~n3518 ) ;
  assign n3520 = ( x65 & n3318 ) | ( x65 & n3509 ) | ( n3318 & n3509 ) ;
  assign n3521 = x65 | n3318 ;
  assign n3522 = ( ~n3322 & n3520 ) | ( ~n3322 & n3521 ) | ( n3520 & n3521 ) ;
  assign n3523 = ( n3322 & n3520 ) | ( n3322 & n3521 ) | ( n3520 & n3521 ) ;
  assign n3524 = ( n3322 & n3522 ) | ( n3322 & ~n3523 ) | ( n3522 & ~n3523 ) ;
  assign n3525 = ( x66 & n3519 ) | ( x66 & ~n3524 ) | ( n3519 & ~n3524 ) ;
  assign n3526 = ( x66 & n3323 ) | ( x66 & n3509 ) | ( n3323 & n3509 ) ;
  assign n3527 = x66 | n3323 ;
  assign n3528 = ( ~n3328 & n3526 ) | ( ~n3328 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3529 = ( n3328 & n3526 ) | ( n3328 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3530 = ( n3328 & n3528 ) | ( n3328 & ~n3529 ) | ( n3528 & ~n3529 ) ;
  assign n3531 = ( x67 & n3525 ) | ( x67 & ~n3530 ) | ( n3525 & ~n3530 ) ;
  assign n3532 = ( x67 & n3329 ) | ( x67 & ~n3509 ) | ( n3329 & ~n3509 ) ;
  assign n3533 = x67 & n3329 ;
  assign n3534 = ( ~n3334 & n3532 ) | ( ~n3334 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3535 = ( n3334 & n3532 ) | ( n3334 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3536 = ( n3334 & n3534 ) | ( n3334 & ~n3535 ) | ( n3534 & ~n3535 ) ;
  assign n3537 = ( x68 & n3531 ) | ( x68 & ~n3536 ) | ( n3531 & ~n3536 ) ;
  assign n3538 = ( x68 & n3335 ) | ( x68 & ~n3509 ) | ( n3335 & ~n3509 ) ;
  assign n3539 = x68 & n3335 ;
  assign n3540 = ( ~n3340 & n3538 ) | ( ~n3340 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3541 = ( n3340 & n3538 ) | ( n3340 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3542 = ( n3340 & n3540 ) | ( n3340 & ~n3541 ) | ( n3540 & ~n3541 ) ;
  assign n3543 = ( x69 & n3537 ) | ( x69 & ~n3542 ) | ( n3537 & ~n3542 ) ;
  assign n3544 = ( x69 & n3341 ) | ( x69 & ~n3509 ) | ( n3341 & ~n3509 ) ;
  assign n3545 = x69 & n3341 ;
  assign n3546 = ( ~n3346 & n3544 ) | ( ~n3346 & n3545 ) | ( n3544 & n3545 ) ;
  assign n3547 = ( n3346 & n3544 ) | ( n3346 & n3545 ) | ( n3544 & n3545 ) ;
  assign n3548 = ( n3346 & n3546 ) | ( n3346 & ~n3547 ) | ( n3546 & ~n3547 ) ;
  assign n3549 = ( x70 & n3543 ) | ( x70 & ~n3548 ) | ( n3543 & ~n3548 ) ;
  assign n3550 = ( x70 & n3347 ) | ( x70 & ~n3509 ) | ( n3347 & ~n3509 ) ;
  assign n3551 = x70 & n3347 ;
  assign n3552 = ( ~n3352 & n3550 ) | ( ~n3352 & n3551 ) | ( n3550 & n3551 ) ;
  assign n3553 = ( n3352 & n3550 ) | ( n3352 & n3551 ) | ( n3550 & n3551 ) ;
  assign n3554 = ( n3352 & n3552 ) | ( n3352 & ~n3553 ) | ( n3552 & ~n3553 ) ;
  assign n3555 = ( x71 & n3549 ) | ( x71 & ~n3554 ) | ( n3549 & ~n3554 ) ;
  assign n3556 = ( x71 & n3353 ) | ( x71 & ~n3509 ) | ( n3353 & ~n3509 ) ;
  assign n3557 = x71 & n3353 ;
  assign n3558 = ( ~n3358 & n3556 ) | ( ~n3358 & n3557 ) | ( n3556 & n3557 ) ;
  assign n3559 = ( n3358 & n3556 ) | ( n3358 & n3557 ) | ( n3556 & n3557 ) ;
  assign n3560 = ( n3358 & n3558 ) | ( n3358 & ~n3559 ) | ( n3558 & ~n3559 ) ;
  assign n3561 = ( x72 & n3555 ) | ( x72 & ~n3560 ) | ( n3555 & ~n3560 ) ;
  assign n3562 = ( x72 & n3359 ) | ( x72 & ~n3509 ) | ( n3359 & ~n3509 ) ;
  assign n3563 = x72 & n3359 ;
  assign n3564 = ( ~n3364 & n3562 ) | ( ~n3364 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ( n3364 & n3562 ) | ( n3364 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3566 = ( n3364 & n3564 ) | ( n3364 & ~n3565 ) | ( n3564 & ~n3565 ) ;
  assign n3567 = ( x73 & n3561 ) | ( x73 & ~n3566 ) | ( n3561 & ~n3566 ) ;
  assign n3568 = ( x73 & n3365 ) | ( x73 & ~n3509 ) | ( n3365 & ~n3509 ) ;
  assign n3569 = x73 & n3365 ;
  assign n3570 = ( ~n3370 & n3568 ) | ( ~n3370 & n3569 ) | ( n3568 & n3569 ) ;
  assign n3571 = ( n3370 & n3568 ) | ( n3370 & n3569 ) | ( n3568 & n3569 ) ;
  assign n3572 = ( n3370 & n3570 ) | ( n3370 & ~n3571 ) | ( n3570 & ~n3571 ) ;
  assign n3573 = ( x74 & n3567 ) | ( x74 & ~n3572 ) | ( n3567 & ~n3572 ) ;
  assign n3574 = ( x74 & n3371 ) | ( x74 & ~n3509 ) | ( n3371 & ~n3509 ) ;
  assign n3575 = x74 & n3371 ;
  assign n3576 = ( ~n3376 & n3574 ) | ( ~n3376 & n3575 ) | ( n3574 & n3575 ) ;
  assign n3577 = ( n3376 & n3574 ) | ( n3376 & n3575 ) | ( n3574 & n3575 ) ;
  assign n3578 = ( n3376 & n3576 ) | ( n3376 & ~n3577 ) | ( n3576 & ~n3577 ) ;
  assign n3579 = ( x75 & n3573 ) | ( x75 & ~n3578 ) | ( n3573 & ~n3578 ) ;
  assign n3580 = ( x75 & n3377 ) | ( x75 & ~n3509 ) | ( n3377 & ~n3509 ) ;
  assign n3581 = x75 & n3377 ;
  assign n3582 = ( ~n3382 & n3580 ) | ( ~n3382 & n3581 ) | ( n3580 & n3581 ) ;
  assign n3583 = ( n3382 & n3580 ) | ( n3382 & n3581 ) | ( n3580 & n3581 ) ;
  assign n3584 = ( n3382 & n3582 ) | ( n3382 & ~n3583 ) | ( n3582 & ~n3583 ) ;
  assign n3585 = ( x76 & n3579 ) | ( x76 & ~n3584 ) | ( n3579 & ~n3584 ) ;
  assign n3586 = ( x76 & n3383 ) | ( x76 & ~n3509 ) | ( n3383 & ~n3509 ) ;
  assign n3587 = x76 & n3383 ;
  assign n3588 = ( ~n3388 & n3586 ) | ( ~n3388 & n3587 ) | ( n3586 & n3587 ) ;
  assign n3589 = ( n3388 & n3586 ) | ( n3388 & n3587 ) | ( n3586 & n3587 ) ;
  assign n3590 = ( n3388 & n3588 ) | ( n3388 & ~n3589 ) | ( n3588 & ~n3589 ) ;
  assign n3591 = ( x77 & n3585 ) | ( x77 & ~n3590 ) | ( n3585 & ~n3590 ) ;
  assign n3592 = ( x77 & n3389 ) | ( x77 & ~n3509 ) | ( n3389 & ~n3509 ) ;
  assign n3593 = x77 & n3389 ;
  assign n3594 = ( ~n3394 & n3592 ) | ( ~n3394 & n3593 ) | ( n3592 & n3593 ) ;
  assign n3595 = ( n3394 & n3592 ) | ( n3394 & n3593 ) | ( n3592 & n3593 ) ;
  assign n3596 = ( n3394 & n3594 ) | ( n3394 & ~n3595 ) | ( n3594 & ~n3595 ) ;
  assign n3597 = ( x78 & n3591 ) | ( x78 & ~n3596 ) | ( n3591 & ~n3596 ) ;
  assign n3598 = ( x78 & n3395 ) | ( x78 & ~n3509 ) | ( n3395 & ~n3509 ) ;
  assign n3599 = x78 & n3395 ;
  assign n3600 = ( ~n3400 & n3598 ) | ( ~n3400 & n3599 ) | ( n3598 & n3599 ) ;
  assign n3601 = ( n3400 & n3598 ) | ( n3400 & n3599 ) | ( n3598 & n3599 ) ;
  assign n3602 = ( n3400 & n3600 ) | ( n3400 & ~n3601 ) | ( n3600 & ~n3601 ) ;
  assign n3603 = ( x79 & n3597 ) | ( x79 & ~n3602 ) | ( n3597 & ~n3602 ) ;
  assign n3604 = ( x79 & n3401 ) | ( x79 & ~n3509 ) | ( n3401 & ~n3509 ) ;
  assign n3605 = x79 & n3401 ;
  assign n3606 = ( ~n3406 & n3604 ) | ( ~n3406 & n3605 ) | ( n3604 & n3605 ) ;
  assign n3607 = ( n3406 & n3604 ) | ( n3406 & n3605 ) | ( n3604 & n3605 ) ;
  assign n3608 = ( n3406 & n3606 ) | ( n3406 & ~n3607 ) | ( n3606 & ~n3607 ) ;
  assign n3609 = ( x80 & n3603 ) | ( x80 & ~n3608 ) | ( n3603 & ~n3608 ) ;
  assign n3610 = ( x80 & n3407 ) | ( x80 & ~n3509 ) | ( n3407 & ~n3509 ) ;
  assign n3611 = x80 & n3407 ;
  assign n3612 = ( ~n3412 & n3610 ) | ( ~n3412 & n3611 ) | ( n3610 & n3611 ) ;
  assign n3613 = ( n3412 & n3610 ) | ( n3412 & n3611 ) | ( n3610 & n3611 ) ;
  assign n3614 = ( n3412 & n3612 ) | ( n3412 & ~n3613 ) | ( n3612 & ~n3613 ) ;
  assign n3615 = ( x81 & n3609 ) | ( x81 & ~n3614 ) | ( n3609 & ~n3614 ) ;
  assign n3616 = ( x81 & n3413 ) | ( x81 & ~n3509 ) | ( n3413 & ~n3509 ) ;
  assign n3617 = x81 & n3413 ;
  assign n3618 = ( ~n3418 & n3616 ) | ( ~n3418 & n3617 ) | ( n3616 & n3617 ) ;
  assign n3619 = ( n3418 & n3616 ) | ( n3418 & n3617 ) | ( n3616 & n3617 ) ;
  assign n3620 = ( n3418 & n3618 ) | ( n3418 & ~n3619 ) | ( n3618 & ~n3619 ) ;
  assign n3621 = ( x82 & n3615 ) | ( x82 & ~n3620 ) | ( n3615 & ~n3620 ) ;
  assign n3622 = ( x82 & n3419 ) | ( x82 & ~n3509 ) | ( n3419 & ~n3509 ) ;
  assign n3623 = x82 & n3419 ;
  assign n3624 = ( ~n3424 & n3622 ) | ( ~n3424 & n3623 ) | ( n3622 & n3623 ) ;
  assign n3625 = ( n3424 & n3622 ) | ( n3424 & n3623 ) | ( n3622 & n3623 ) ;
  assign n3626 = ( n3424 & n3624 ) | ( n3424 & ~n3625 ) | ( n3624 & ~n3625 ) ;
  assign n3627 = ( x83 & n3621 ) | ( x83 & ~n3626 ) | ( n3621 & ~n3626 ) ;
  assign n3628 = ( x83 & n3425 ) | ( x83 & ~n3509 ) | ( n3425 & ~n3509 ) ;
  assign n3629 = x83 & n3425 ;
  assign n3630 = ( ~n3430 & n3628 ) | ( ~n3430 & n3629 ) | ( n3628 & n3629 ) ;
  assign n3631 = ( n3430 & n3628 ) | ( n3430 & n3629 ) | ( n3628 & n3629 ) ;
  assign n3632 = ( n3430 & n3630 ) | ( n3430 & ~n3631 ) | ( n3630 & ~n3631 ) ;
  assign n3633 = ( x84 & n3627 ) | ( x84 & ~n3632 ) | ( n3627 & ~n3632 ) ;
  assign n3634 = ( x84 & n3431 ) | ( x84 & ~n3509 ) | ( n3431 & ~n3509 ) ;
  assign n3635 = x84 & n3431 ;
  assign n3636 = ( ~n3436 & n3634 ) | ( ~n3436 & n3635 ) | ( n3634 & n3635 ) ;
  assign n3637 = ( n3436 & n3634 ) | ( n3436 & n3635 ) | ( n3634 & n3635 ) ;
  assign n3638 = ( n3436 & n3636 ) | ( n3436 & ~n3637 ) | ( n3636 & ~n3637 ) ;
  assign n3639 = ( x85 & n3633 ) | ( x85 & ~n3638 ) | ( n3633 & ~n3638 ) ;
  assign n3640 = ( x85 & n3437 ) | ( x85 & ~n3509 ) | ( n3437 & ~n3509 ) ;
  assign n3641 = x85 & n3437 ;
  assign n3642 = ( ~n3442 & n3640 ) | ( ~n3442 & n3641 ) | ( n3640 & n3641 ) ;
  assign n3643 = ( n3442 & n3640 ) | ( n3442 & n3641 ) | ( n3640 & n3641 ) ;
  assign n3644 = ( n3442 & n3642 ) | ( n3442 & ~n3643 ) | ( n3642 & ~n3643 ) ;
  assign n3645 = ( x86 & n3639 ) | ( x86 & ~n3644 ) | ( n3639 & ~n3644 ) ;
  assign n3646 = ( x86 & n3443 ) | ( x86 & ~n3509 ) | ( n3443 & ~n3509 ) ;
  assign n3647 = x86 & n3443 ;
  assign n3648 = ( ~n3448 & n3646 ) | ( ~n3448 & n3647 ) | ( n3646 & n3647 ) ;
  assign n3649 = ( n3448 & n3646 ) | ( n3448 & n3647 ) | ( n3646 & n3647 ) ;
  assign n3650 = ( n3448 & n3648 ) | ( n3448 & ~n3649 ) | ( n3648 & ~n3649 ) ;
  assign n3651 = ( x87 & n3645 ) | ( x87 & ~n3650 ) | ( n3645 & ~n3650 ) ;
  assign n3652 = ( x87 & n3449 ) | ( x87 & ~n3509 ) | ( n3449 & ~n3509 ) ;
  assign n3653 = x87 & n3449 ;
  assign n3654 = ( ~n3454 & n3652 ) | ( ~n3454 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = ( n3454 & n3652 ) | ( n3454 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3656 = ( n3454 & n3654 ) | ( n3454 & ~n3655 ) | ( n3654 & ~n3655 ) ;
  assign n3657 = ( x88 & n3651 ) | ( x88 & ~n3656 ) | ( n3651 & ~n3656 ) ;
  assign n3658 = ( x88 & n3455 ) | ( x88 & ~n3509 ) | ( n3455 & ~n3509 ) ;
  assign n3659 = x88 & n3455 ;
  assign n3660 = ( ~n3460 & n3658 ) | ( ~n3460 & n3659 ) | ( n3658 & n3659 ) ;
  assign n3661 = ( n3460 & n3658 ) | ( n3460 & n3659 ) | ( n3658 & n3659 ) ;
  assign n3662 = ( n3460 & n3660 ) | ( n3460 & ~n3661 ) | ( n3660 & ~n3661 ) ;
  assign n3663 = ( x89 & n3657 ) | ( x89 & ~n3662 ) | ( n3657 & ~n3662 ) ;
  assign n3664 = ( x89 & n3461 ) | ( x89 & ~n3509 ) | ( n3461 & ~n3509 ) ;
  assign n3665 = x89 & n3461 ;
  assign n3666 = ( ~n3466 & n3664 ) | ( ~n3466 & n3665 ) | ( n3664 & n3665 ) ;
  assign n3667 = ( n3466 & n3664 ) | ( n3466 & n3665 ) | ( n3664 & n3665 ) ;
  assign n3668 = ( n3466 & n3666 ) | ( n3466 & ~n3667 ) | ( n3666 & ~n3667 ) ;
  assign n3669 = ( x90 & n3663 ) | ( x90 & ~n3668 ) | ( n3663 & ~n3668 ) ;
  assign n3670 = ( x90 & n3467 ) | ( x90 & ~n3509 ) | ( n3467 & ~n3509 ) ;
  assign n3671 = x90 & n3467 ;
  assign n3672 = ( ~n3472 & n3670 ) | ( ~n3472 & n3671 ) | ( n3670 & n3671 ) ;
  assign n3673 = ( n3472 & n3670 ) | ( n3472 & n3671 ) | ( n3670 & n3671 ) ;
  assign n3674 = ( n3472 & n3672 ) | ( n3472 & ~n3673 ) | ( n3672 & ~n3673 ) ;
  assign n3675 = ( x91 & n3669 ) | ( x91 & ~n3674 ) | ( n3669 & ~n3674 ) ;
  assign n3676 = ( x91 & n3473 ) | ( x91 & ~n3509 ) | ( n3473 & ~n3509 ) ;
  assign n3677 = x91 & n3473 ;
  assign n3678 = ( ~n3478 & n3676 ) | ( ~n3478 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3679 = ( n3478 & n3676 ) | ( n3478 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3680 = ( n3478 & n3678 ) | ( n3478 & ~n3679 ) | ( n3678 & ~n3679 ) ;
  assign n3681 = ( x92 & n3675 ) | ( x92 & ~n3680 ) | ( n3675 & ~n3680 ) ;
  assign n3682 = ( x92 & n3479 ) | ( x92 & ~n3509 ) | ( n3479 & ~n3509 ) ;
  assign n3683 = x92 & n3479 ;
  assign n3684 = ( ~n3484 & n3682 ) | ( ~n3484 & n3683 ) | ( n3682 & n3683 ) ;
  assign n3685 = ( n3484 & n3682 ) | ( n3484 & n3683 ) | ( n3682 & n3683 ) ;
  assign n3686 = ( n3484 & n3684 ) | ( n3484 & ~n3685 ) | ( n3684 & ~n3685 ) ;
  assign n3687 = ( x93 & n3681 ) | ( x93 & ~n3686 ) | ( n3681 & ~n3686 ) ;
  assign n3688 = ( x93 & n3485 ) | ( x93 & ~n3509 ) | ( n3485 & ~n3509 ) ;
  assign n3689 = x93 & n3485 ;
  assign n3690 = ( ~n3490 & n3688 ) | ( ~n3490 & n3689 ) | ( n3688 & n3689 ) ;
  assign n3691 = ( n3490 & n3688 ) | ( n3490 & n3689 ) | ( n3688 & n3689 ) ;
  assign n3692 = ( n3490 & n3690 ) | ( n3490 & ~n3691 ) | ( n3690 & ~n3691 ) ;
  assign n3693 = ( x94 & n3687 ) | ( x94 & ~n3692 ) | ( n3687 & ~n3692 ) ;
  assign n3694 = ( x94 & n3491 ) | ( x94 & ~n3509 ) | ( n3491 & ~n3509 ) ;
  assign n3695 = x94 & n3491 ;
  assign n3696 = ( ~n3496 & n3694 ) | ( ~n3496 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = ( n3496 & n3694 ) | ( n3496 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3698 = ( n3496 & n3696 ) | ( n3496 & ~n3697 ) | ( n3696 & ~n3697 ) ;
  assign n3699 = ( x95 & n3693 ) | ( x95 & ~n3698 ) | ( n3693 & ~n3698 ) ;
  assign n3700 = ( x95 & n3497 ) | ( x95 & ~n3509 ) | ( n3497 & ~n3509 ) ;
  assign n3701 = x95 & n3497 ;
  assign n3702 = ( ~n3502 & n3700 ) | ( ~n3502 & n3701 ) | ( n3700 & n3701 ) ;
  assign n3703 = ( n3502 & n3700 ) | ( n3502 & n3701 ) | ( n3700 & n3701 ) ;
  assign n3704 = ( n3502 & n3702 ) | ( n3502 & ~n3703 ) | ( n3702 & ~n3703 ) ;
  assign n3705 = ( x96 & n3699 ) | ( x96 & ~n3704 ) | ( n3699 & ~n3704 ) ;
  assign n3706 = ( x97 & n159 ) | ( x97 & n3504 ) | ( n159 & n3504 ) ;
  assign n3707 = x97 | n3504 ;
  assign n3708 = ( n3507 & n3706 ) | ( n3507 & ~n3707 ) | ( n3706 & ~n3707 ) ;
  assign n3709 = ( x97 & ~n3514 ) | ( x97 & n3705 ) | ( ~n3514 & n3705 ) ;
  assign n3710 = ( x98 & ~n3708 ) | ( x98 & n3709 ) | ( ~n3708 & n3709 ) ;
  assign n3711 = n158 | n3710 ;
  assign n3712 = ( x97 & n3705 ) | ( x97 & n3711 ) | ( n3705 & n3711 ) ;
  assign n3713 = x97 | n3705 ;
  assign n3714 = ( ~n3514 & n3712 ) | ( ~n3514 & n3713 ) | ( n3712 & n3713 ) ;
  assign n3715 = ( n3514 & n3712 ) | ( n3514 & n3713 ) | ( n3712 & n3713 ) ;
  assign n3716 = ( n3514 & n3714 ) | ( n3514 & ~n3715 ) | ( n3714 & ~n3715 ) ;
  assign n3717 = ~x28 & x64 ;
  assign n3718 = ~x29 & n3711 ;
  assign n3719 = ( x29 & ~x64 ) | ( x29 & n3711 ) | ( ~x64 & n3711 ) ;
  assign n3720 = ( n3515 & ~n3718 ) | ( n3515 & n3719 ) | ( ~n3718 & n3719 ) ;
  assign n3721 = ( x65 & n3717 ) | ( x65 & ~n3720 ) | ( n3717 & ~n3720 ) ;
  assign n3722 = ( x65 & n3515 ) | ( x65 & n3711 ) | ( n3515 & n3711 ) ;
  assign n3723 = x65 | n3515 ;
  assign n3724 = ( ~n3518 & n3722 ) | ( ~n3518 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = ( n3518 & n3722 ) | ( n3518 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3726 = ( n3518 & n3724 ) | ( n3518 & ~n3725 ) | ( n3724 & ~n3725 ) ;
  assign n3727 = ( x66 & n3721 ) | ( x66 & ~n3726 ) | ( n3721 & ~n3726 ) ;
  assign n3728 = ( x66 & n3519 ) | ( x66 & n3711 ) | ( n3519 & n3711 ) ;
  assign n3729 = x66 | n3519 ;
  assign n3730 = ( ~n3524 & n3728 ) | ( ~n3524 & n3729 ) | ( n3728 & n3729 ) ;
  assign n3731 = ( n3524 & n3728 ) | ( n3524 & n3729 ) | ( n3728 & n3729 ) ;
  assign n3732 = ( n3524 & n3730 ) | ( n3524 & ~n3731 ) | ( n3730 & ~n3731 ) ;
  assign n3733 = ( x67 & n3727 ) | ( x67 & ~n3732 ) | ( n3727 & ~n3732 ) ;
  assign n3734 = ( x67 & n3525 ) | ( x67 & ~n3711 ) | ( n3525 & ~n3711 ) ;
  assign n3735 = x67 & n3525 ;
  assign n3736 = ( ~n3530 & n3734 ) | ( ~n3530 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = ( n3530 & n3734 ) | ( n3530 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3738 = ( n3530 & n3736 ) | ( n3530 & ~n3737 ) | ( n3736 & ~n3737 ) ;
  assign n3739 = ( x68 & n3733 ) | ( x68 & ~n3738 ) | ( n3733 & ~n3738 ) ;
  assign n3740 = ( x68 & n3531 ) | ( x68 & ~n3711 ) | ( n3531 & ~n3711 ) ;
  assign n3741 = x68 & n3531 ;
  assign n3742 = ( ~n3536 & n3740 ) | ( ~n3536 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3743 = ( n3536 & n3740 ) | ( n3536 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3744 = ( n3536 & n3742 ) | ( n3536 & ~n3743 ) | ( n3742 & ~n3743 ) ;
  assign n3745 = ( x69 & n3739 ) | ( x69 & ~n3744 ) | ( n3739 & ~n3744 ) ;
  assign n3746 = ( x69 & n3537 ) | ( x69 & ~n3711 ) | ( n3537 & ~n3711 ) ;
  assign n3747 = x69 & n3537 ;
  assign n3748 = ( ~n3542 & n3746 ) | ( ~n3542 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3749 = ( n3542 & n3746 ) | ( n3542 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3750 = ( n3542 & n3748 ) | ( n3542 & ~n3749 ) | ( n3748 & ~n3749 ) ;
  assign n3751 = ( x70 & n3745 ) | ( x70 & ~n3750 ) | ( n3745 & ~n3750 ) ;
  assign n3752 = ( x70 & n3543 ) | ( x70 & ~n3711 ) | ( n3543 & ~n3711 ) ;
  assign n3753 = x70 & n3543 ;
  assign n3754 = ( ~n3548 & n3752 ) | ( ~n3548 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = ( n3548 & n3752 ) | ( n3548 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3756 = ( n3548 & n3754 ) | ( n3548 & ~n3755 ) | ( n3754 & ~n3755 ) ;
  assign n3757 = ( x71 & n3751 ) | ( x71 & ~n3756 ) | ( n3751 & ~n3756 ) ;
  assign n3758 = ( x71 & n3549 ) | ( x71 & ~n3711 ) | ( n3549 & ~n3711 ) ;
  assign n3759 = x71 & n3549 ;
  assign n3760 = ( ~n3554 & n3758 ) | ( ~n3554 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3761 = ( n3554 & n3758 ) | ( n3554 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3762 = ( n3554 & n3760 ) | ( n3554 & ~n3761 ) | ( n3760 & ~n3761 ) ;
  assign n3763 = ( x72 & n3757 ) | ( x72 & ~n3762 ) | ( n3757 & ~n3762 ) ;
  assign n3764 = ( x72 & n3555 ) | ( x72 & ~n3711 ) | ( n3555 & ~n3711 ) ;
  assign n3765 = x72 & n3555 ;
  assign n3766 = ( ~n3560 & n3764 ) | ( ~n3560 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3767 = ( n3560 & n3764 ) | ( n3560 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3768 = ( n3560 & n3766 ) | ( n3560 & ~n3767 ) | ( n3766 & ~n3767 ) ;
  assign n3769 = ( x73 & n3763 ) | ( x73 & ~n3768 ) | ( n3763 & ~n3768 ) ;
  assign n3770 = ( x73 & n3561 ) | ( x73 & ~n3711 ) | ( n3561 & ~n3711 ) ;
  assign n3771 = x73 & n3561 ;
  assign n3772 = ( ~n3566 & n3770 ) | ( ~n3566 & n3771 ) | ( n3770 & n3771 ) ;
  assign n3773 = ( n3566 & n3770 ) | ( n3566 & n3771 ) | ( n3770 & n3771 ) ;
  assign n3774 = ( n3566 & n3772 ) | ( n3566 & ~n3773 ) | ( n3772 & ~n3773 ) ;
  assign n3775 = ( x74 & n3769 ) | ( x74 & ~n3774 ) | ( n3769 & ~n3774 ) ;
  assign n3776 = ( x74 & n3567 ) | ( x74 & ~n3711 ) | ( n3567 & ~n3711 ) ;
  assign n3777 = x74 & n3567 ;
  assign n3778 = ( ~n3572 & n3776 ) | ( ~n3572 & n3777 ) | ( n3776 & n3777 ) ;
  assign n3779 = ( n3572 & n3776 ) | ( n3572 & n3777 ) | ( n3776 & n3777 ) ;
  assign n3780 = ( n3572 & n3778 ) | ( n3572 & ~n3779 ) | ( n3778 & ~n3779 ) ;
  assign n3781 = ( x75 & n3775 ) | ( x75 & ~n3780 ) | ( n3775 & ~n3780 ) ;
  assign n3782 = ( x75 & n3573 ) | ( x75 & ~n3711 ) | ( n3573 & ~n3711 ) ;
  assign n3783 = x75 & n3573 ;
  assign n3784 = ( ~n3578 & n3782 ) | ( ~n3578 & n3783 ) | ( n3782 & n3783 ) ;
  assign n3785 = ( n3578 & n3782 ) | ( n3578 & n3783 ) | ( n3782 & n3783 ) ;
  assign n3786 = ( n3578 & n3784 ) | ( n3578 & ~n3785 ) | ( n3784 & ~n3785 ) ;
  assign n3787 = ( x76 & n3781 ) | ( x76 & ~n3786 ) | ( n3781 & ~n3786 ) ;
  assign n3788 = ( x76 & n3579 ) | ( x76 & ~n3711 ) | ( n3579 & ~n3711 ) ;
  assign n3789 = x76 & n3579 ;
  assign n3790 = ( ~n3584 & n3788 ) | ( ~n3584 & n3789 ) | ( n3788 & n3789 ) ;
  assign n3791 = ( n3584 & n3788 ) | ( n3584 & n3789 ) | ( n3788 & n3789 ) ;
  assign n3792 = ( n3584 & n3790 ) | ( n3584 & ~n3791 ) | ( n3790 & ~n3791 ) ;
  assign n3793 = ( x77 & n3787 ) | ( x77 & ~n3792 ) | ( n3787 & ~n3792 ) ;
  assign n3794 = ( x77 & n3585 ) | ( x77 & ~n3711 ) | ( n3585 & ~n3711 ) ;
  assign n3795 = x77 & n3585 ;
  assign n3796 = ( ~n3590 & n3794 ) | ( ~n3590 & n3795 ) | ( n3794 & n3795 ) ;
  assign n3797 = ( n3590 & n3794 ) | ( n3590 & n3795 ) | ( n3794 & n3795 ) ;
  assign n3798 = ( n3590 & n3796 ) | ( n3590 & ~n3797 ) | ( n3796 & ~n3797 ) ;
  assign n3799 = ( x78 & n3793 ) | ( x78 & ~n3798 ) | ( n3793 & ~n3798 ) ;
  assign n3800 = ( x78 & n3591 ) | ( x78 & ~n3711 ) | ( n3591 & ~n3711 ) ;
  assign n3801 = x78 & n3591 ;
  assign n3802 = ( ~n3596 & n3800 ) | ( ~n3596 & n3801 ) | ( n3800 & n3801 ) ;
  assign n3803 = ( n3596 & n3800 ) | ( n3596 & n3801 ) | ( n3800 & n3801 ) ;
  assign n3804 = ( n3596 & n3802 ) | ( n3596 & ~n3803 ) | ( n3802 & ~n3803 ) ;
  assign n3805 = ( x79 & n3799 ) | ( x79 & ~n3804 ) | ( n3799 & ~n3804 ) ;
  assign n3806 = ( x79 & n3597 ) | ( x79 & ~n3711 ) | ( n3597 & ~n3711 ) ;
  assign n3807 = x79 & n3597 ;
  assign n3808 = ( ~n3602 & n3806 ) | ( ~n3602 & n3807 ) | ( n3806 & n3807 ) ;
  assign n3809 = ( n3602 & n3806 ) | ( n3602 & n3807 ) | ( n3806 & n3807 ) ;
  assign n3810 = ( n3602 & n3808 ) | ( n3602 & ~n3809 ) | ( n3808 & ~n3809 ) ;
  assign n3811 = ( x80 & n3805 ) | ( x80 & ~n3810 ) | ( n3805 & ~n3810 ) ;
  assign n3812 = ( x80 & n3603 ) | ( x80 & ~n3711 ) | ( n3603 & ~n3711 ) ;
  assign n3813 = x80 & n3603 ;
  assign n3814 = ( ~n3608 & n3812 ) | ( ~n3608 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3815 = ( n3608 & n3812 ) | ( n3608 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3816 = ( n3608 & n3814 ) | ( n3608 & ~n3815 ) | ( n3814 & ~n3815 ) ;
  assign n3817 = ( x81 & n3811 ) | ( x81 & ~n3816 ) | ( n3811 & ~n3816 ) ;
  assign n3818 = ( x81 & n3609 ) | ( x81 & ~n3711 ) | ( n3609 & ~n3711 ) ;
  assign n3819 = x81 & n3609 ;
  assign n3820 = ( ~n3614 & n3818 ) | ( ~n3614 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3821 = ( n3614 & n3818 ) | ( n3614 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3822 = ( n3614 & n3820 ) | ( n3614 & ~n3821 ) | ( n3820 & ~n3821 ) ;
  assign n3823 = ( x82 & n3817 ) | ( x82 & ~n3822 ) | ( n3817 & ~n3822 ) ;
  assign n3824 = ( x82 & n3615 ) | ( x82 & ~n3711 ) | ( n3615 & ~n3711 ) ;
  assign n3825 = x82 & n3615 ;
  assign n3826 = ( ~n3620 & n3824 ) | ( ~n3620 & n3825 ) | ( n3824 & n3825 ) ;
  assign n3827 = ( n3620 & n3824 ) | ( n3620 & n3825 ) | ( n3824 & n3825 ) ;
  assign n3828 = ( n3620 & n3826 ) | ( n3620 & ~n3827 ) | ( n3826 & ~n3827 ) ;
  assign n3829 = ( x83 & n3823 ) | ( x83 & ~n3828 ) | ( n3823 & ~n3828 ) ;
  assign n3830 = ( x83 & n3621 ) | ( x83 & ~n3711 ) | ( n3621 & ~n3711 ) ;
  assign n3831 = x83 & n3621 ;
  assign n3832 = ( ~n3626 & n3830 ) | ( ~n3626 & n3831 ) | ( n3830 & n3831 ) ;
  assign n3833 = ( n3626 & n3830 ) | ( n3626 & n3831 ) | ( n3830 & n3831 ) ;
  assign n3834 = ( n3626 & n3832 ) | ( n3626 & ~n3833 ) | ( n3832 & ~n3833 ) ;
  assign n3835 = ( x84 & n3829 ) | ( x84 & ~n3834 ) | ( n3829 & ~n3834 ) ;
  assign n3836 = ( x84 & n3627 ) | ( x84 & ~n3711 ) | ( n3627 & ~n3711 ) ;
  assign n3837 = x84 & n3627 ;
  assign n3838 = ( ~n3632 & n3836 ) | ( ~n3632 & n3837 ) | ( n3836 & n3837 ) ;
  assign n3839 = ( n3632 & n3836 ) | ( n3632 & n3837 ) | ( n3836 & n3837 ) ;
  assign n3840 = ( n3632 & n3838 ) | ( n3632 & ~n3839 ) | ( n3838 & ~n3839 ) ;
  assign n3841 = ( x85 & n3835 ) | ( x85 & ~n3840 ) | ( n3835 & ~n3840 ) ;
  assign n3842 = ( x85 & n3633 ) | ( x85 & ~n3711 ) | ( n3633 & ~n3711 ) ;
  assign n3843 = x85 & n3633 ;
  assign n3844 = ( ~n3638 & n3842 ) | ( ~n3638 & n3843 ) | ( n3842 & n3843 ) ;
  assign n3845 = ( n3638 & n3842 ) | ( n3638 & n3843 ) | ( n3842 & n3843 ) ;
  assign n3846 = ( n3638 & n3844 ) | ( n3638 & ~n3845 ) | ( n3844 & ~n3845 ) ;
  assign n3847 = ( x86 & n3841 ) | ( x86 & ~n3846 ) | ( n3841 & ~n3846 ) ;
  assign n3848 = ( x86 & n3639 ) | ( x86 & ~n3711 ) | ( n3639 & ~n3711 ) ;
  assign n3849 = x86 & n3639 ;
  assign n3850 = ( ~n3644 & n3848 ) | ( ~n3644 & n3849 ) | ( n3848 & n3849 ) ;
  assign n3851 = ( n3644 & n3848 ) | ( n3644 & n3849 ) | ( n3848 & n3849 ) ;
  assign n3852 = ( n3644 & n3850 ) | ( n3644 & ~n3851 ) | ( n3850 & ~n3851 ) ;
  assign n3853 = ( x87 & n3847 ) | ( x87 & ~n3852 ) | ( n3847 & ~n3852 ) ;
  assign n3854 = ( x87 & n3645 ) | ( x87 & ~n3711 ) | ( n3645 & ~n3711 ) ;
  assign n3855 = x87 & n3645 ;
  assign n3856 = ( ~n3650 & n3854 ) | ( ~n3650 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = ( n3650 & n3854 ) | ( n3650 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3858 = ( n3650 & n3856 ) | ( n3650 & ~n3857 ) | ( n3856 & ~n3857 ) ;
  assign n3859 = ( x88 & n3853 ) | ( x88 & ~n3858 ) | ( n3853 & ~n3858 ) ;
  assign n3860 = ( x88 & n3651 ) | ( x88 & ~n3711 ) | ( n3651 & ~n3711 ) ;
  assign n3861 = x88 & n3651 ;
  assign n3862 = ( ~n3656 & n3860 ) | ( ~n3656 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3863 = ( n3656 & n3860 ) | ( n3656 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3864 = ( n3656 & n3862 ) | ( n3656 & ~n3863 ) | ( n3862 & ~n3863 ) ;
  assign n3865 = ( x89 & n3859 ) | ( x89 & ~n3864 ) | ( n3859 & ~n3864 ) ;
  assign n3866 = ( x89 & n3657 ) | ( x89 & ~n3711 ) | ( n3657 & ~n3711 ) ;
  assign n3867 = x89 & n3657 ;
  assign n3868 = ( ~n3662 & n3866 ) | ( ~n3662 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = ( n3662 & n3866 ) | ( n3662 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3870 = ( n3662 & n3868 ) | ( n3662 & ~n3869 ) | ( n3868 & ~n3869 ) ;
  assign n3871 = ( x90 & n3865 ) | ( x90 & ~n3870 ) | ( n3865 & ~n3870 ) ;
  assign n3872 = ( x90 & n3663 ) | ( x90 & ~n3711 ) | ( n3663 & ~n3711 ) ;
  assign n3873 = x90 & n3663 ;
  assign n3874 = ( ~n3668 & n3872 ) | ( ~n3668 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = ( n3668 & n3872 ) | ( n3668 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3876 = ( n3668 & n3874 ) | ( n3668 & ~n3875 ) | ( n3874 & ~n3875 ) ;
  assign n3877 = ( x91 & n3871 ) | ( x91 & ~n3876 ) | ( n3871 & ~n3876 ) ;
  assign n3878 = ( x91 & n3669 ) | ( x91 & ~n3711 ) | ( n3669 & ~n3711 ) ;
  assign n3879 = x91 & n3669 ;
  assign n3880 = ( ~n3674 & n3878 ) | ( ~n3674 & n3879 ) | ( n3878 & n3879 ) ;
  assign n3881 = ( n3674 & n3878 ) | ( n3674 & n3879 ) | ( n3878 & n3879 ) ;
  assign n3882 = ( n3674 & n3880 ) | ( n3674 & ~n3881 ) | ( n3880 & ~n3881 ) ;
  assign n3883 = ( x92 & n3877 ) | ( x92 & ~n3882 ) | ( n3877 & ~n3882 ) ;
  assign n3884 = ( x92 & n3675 ) | ( x92 & ~n3711 ) | ( n3675 & ~n3711 ) ;
  assign n3885 = x92 & n3675 ;
  assign n3886 = ( ~n3680 & n3884 ) | ( ~n3680 & n3885 ) | ( n3884 & n3885 ) ;
  assign n3887 = ( n3680 & n3884 ) | ( n3680 & n3885 ) | ( n3884 & n3885 ) ;
  assign n3888 = ( n3680 & n3886 ) | ( n3680 & ~n3887 ) | ( n3886 & ~n3887 ) ;
  assign n3889 = ( x93 & n3883 ) | ( x93 & ~n3888 ) | ( n3883 & ~n3888 ) ;
  assign n3890 = ( x93 & n3681 ) | ( x93 & ~n3711 ) | ( n3681 & ~n3711 ) ;
  assign n3891 = x93 & n3681 ;
  assign n3892 = ( ~n3686 & n3890 ) | ( ~n3686 & n3891 ) | ( n3890 & n3891 ) ;
  assign n3893 = ( n3686 & n3890 ) | ( n3686 & n3891 ) | ( n3890 & n3891 ) ;
  assign n3894 = ( n3686 & n3892 ) | ( n3686 & ~n3893 ) | ( n3892 & ~n3893 ) ;
  assign n3895 = ( x94 & n3889 ) | ( x94 & ~n3894 ) | ( n3889 & ~n3894 ) ;
  assign n3896 = ( x94 & n3687 ) | ( x94 & ~n3711 ) | ( n3687 & ~n3711 ) ;
  assign n3897 = x94 & n3687 ;
  assign n3898 = ( ~n3692 & n3896 ) | ( ~n3692 & n3897 ) | ( n3896 & n3897 ) ;
  assign n3899 = ( n3692 & n3896 ) | ( n3692 & n3897 ) | ( n3896 & n3897 ) ;
  assign n3900 = ( n3692 & n3898 ) | ( n3692 & ~n3899 ) | ( n3898 & ~n3899 ) ;
  assign n3901 = ( x95 & n3895 ) | ( x95 & ~n3900 ) | ( n3895 & ~n3900 ) ;
  assign n3902 = ( x95 & n3693 ) | ( x95 & ~n3711 ) | ( n3693 & ~n3711 ) ;
  assign n3903 = x95 & n3693 ;
  assign n3904 = ( ~n3698 & n3902 ) | ( ~n3698 & n3903 ) | ( n3902 & n3903 ) ;
  assign n3905 = ( n3698 & n3902 ) | ( n3698 & n3903 ) | ( n3902 & n3903 ) ;
  assign n3906 = ( n3698 & n3904 ) | ( n3698 & ~n3905 ) | ( n3904 & ~n3905 ) ;
  assign n3907 = ( x96 & n3901 ) | ( x96 & ~n3906 ) | ( n3901 & ~n3906 ) ;
  assign n3908 = ( x96 & n3699 ) | ( x96 & ~n3711 ) | ( n3699 & ~n3711 ) ;
  assign n3909 = x96 & n3699 ;
  assign n3910 = ( ~n3704 & n3908 ) | ( ~n3704 & n3909 ) | ( n3908 & n3909 ) ;
  assign n3911 = ( n3704 & n3908 ) | ( n3704 & n3909 ) | ( n3908 & n3909 ) ;
  assign n3912 = ( n3704 & n3910 ) | ( n3704 & ~n3911 ) | ( n3910 & ~n3911 ) ;
  assign n3913 = ( x97 & n3907 ) | ( x97 & ~n3912 ) | ( n3907 & ~n3912 ) ;
  assign n3914 = ( ~x98 & n158 ) | ( ~x98 & n3709 ) | ( n158 & n3709 ) ;
  assign n3915 = ( ~x98 & n3708 ) | ( ~x98 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3916 = ~n3914 & n3915 ;
  assign n3917 = ( x98 & ~n3716 ) | ( x98 & n3913 ) | ( ~n3716 & n3913 ) ;
  assign n3918 = n157 | n3917 ;
  assign n3919 = x99 & ~n3708 ;
  assign n3920 = ( ~n3916 & n3918 ) | ( ~n3916 & n3919 ) | ( n3918 & n3919 ) ;
  assign n3921 = ( x98 & n3913 ) | ( x98 & ~n3920 ) | ( n3913 & ~n3920 ) ;
  assign n3922 = x98 & n3913 ;
  assign n3923 = ( ~n3716 & n3921 ) | ( ~n3716 & n3922 ) | ( n3921 & n3922 ) ;
  assign n3924 = ( n3716 & n3921 ) | ( n3716 & n3922 ) | ( n3921 & n3922 ) ;
  assign n3925 = ( n3716 & n3923 ) | ( n3716 & ~n3924 ) | ( n3923 & ~n3924 ) ;
  assign n3926 = ~x27 & x64 ;
  assign n3927 = x28 & n3920 ;
  assign n3928 = ( x28 & x64 ) | ( x28 & ~n3920 ) | ( x64 & ~n3920 ) ;
  assign n3929 = x28 & x64 ;
  assign n3930 = ( n3927 & n3928 ) | ( n3927 & ~n3929 ) | ( n3928 & ~n3929 ) ;
  assign n3931 = ( x65 & n3926 ) | ( x65 & ~n3930 ) | ( n3926 & ~n3930 ) ;
  assign n3932 = ( x65 & n3717 ) | ( x65 & n3920 ) | ( n3717 & n3920 ) ;
  assign n3933 = x65 | n3717 ;
  assign n3934 = ( ~n3720 & n3932 ) | ( ~n3720 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3935 = ( n3720 & n3932 ) | ( n3720 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3936 = ( n3720 & n3934 ) | ( n3720 & ~n3935 ) | ( n3934 & ~n3935 ) ;
  assign n3937 = ( x66 & n3931 ) | ( x66 & ~n3936 ) | ( n3931 & ~n3936 ) ;
  assign n3938 = ( x66 & n3721 ) | ( x66 & n3920 ) | ( n3721 & n3920 ) ;
  assign n3939 = x66 | n3721 ;
  assign n3940 = ( ~n3726 & n3938 ) | ( ~n3726 & n3939 ) | ( n3938 & n3939 ) ;
  assign n3941 = ( n3726 & n3938 ) | ( n3726 & n3939 ) | ( n3938 & n3939 ) ;
  assign n3942 = ( n3726 & n3940 ) | ( n3726 & ~n3941 ) | ( n3940 & ~n3941 ) ;
  assign n3943 = ( x67 & n3937 ) | ( x67 & ~n3942 ) | ( n3937 & ~n3942 ) ;
  assign n3944 = ( x67 & n3727 ) | ( x67 & ~n3920 ) | ( n3727 & ~n3920 ) ;
  assign n3945 = x67 & n3727 ;
  assign n3946 = ( ~n3732 & n3944 ) | ( ~n3732 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3947 = ( n3732 & n3944 ) | ( n3732 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3948 = ( n3732 & n3946 ) | ( n3732 & ~n3947 ) | ( n3946 & ~n3947 ) ;
  assign n3949 = ( x68 & n3943 ) | ( x68 & ~n3948 ) | ( n3943 & ~n3948 ) ;
  assign n3950 = ( x68 & n3733 ) | ( x68 & ~n3920 ) | ( n3733 & ~n3920 ) ;
  assign n3951 = x68 & n3733 ;
  assign n3952 = ( ~n3738 & n3950 ) | ( ~n3738 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3953 = ( n3738 & n3950 ) | ( n3738 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3954 = ( n3738 & n3952 ) | ( n3738 & ~n3953 ) | ( n3952 & ~n3953 ) ;
  assign n3955 = ( x69 & n3949 ) | ( x69 & ~n3954 ) | ( n3949 & ~n3954 ) ;
  assign n3956 = ( x69 & n3739 ) | ( x69 & ~n3920 ) | ( n3739 & ~n3920 ) ;
  assign n3957 = x69 & n3739 ;
  assign n3958 = ( ~n3744 & n3956 ) | ( ~n3744 & n3957 ) | ( n3956 & n3957 ) ;
  assign n3959 = ( n3744 & n3956 ) | ( n3744 & n3957 ) | ( n3956 & n3957 ) ;
  assign n3960 = ( n3744 & n3958 ) | ( n3744 & ~n3959 ) | ( n3958 & ~n3959 ) ;
  assign n3961 = ( x70 & n3955 ) | ( x70 & ~n3960 ) | ( n3955 & ~n3960 ) ;
  assign n3962 = ( x70 & n3745 ) | ( x70 & ~n3920 ) | ( n3745 & ~n3920 ) ;
  assign n3963 = x70 & n3745 ;
  assign n3964 = ( ~n3750 & n3962 ) | ( ~n3750 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3965 = ( n3750 & n3962 ) | ( n3750 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3966 = ( n3750 & n3964 ) | ( n3750 & ~n3965 ) | ( n3964 & ~n3965 ) ;
  assign n3967 = ( x71 & n3961 ) | ( x71 & ~n3966 ) | ( n3961 & ~n3966 ) ;
  assign n3968 = ( x71 & n3751 ) | ( x71 & ~n3920 ) | ( n3751 & ~n3920 ) ;
  assign n3969 = x71 & n3751 ;
  assign n3970 = ( ~n3756 & n3968 ) | ( ~n3756 & n3969 ) | ( n3968 & n3969 ) ;
  assign n3971 = ( n3756 & n3968 ) | ( n3756 & n3969 ) | ( n3968 & n3969 ) ;
  assign n3972 = ( n3756 & n3970 ) | ( n3756 & ~n3971 ) | ( n3970 & ~n3971 ) ;
  assign n3973 = ( x72 & n3967 ) | ( x72 & ~n3972 ) | ( n3967 & ~n3972 ) ;
  assign n3974 = ( x72 & n3757 ) | ( x72 & ~n3920 ) | ( n3757 & ~n3920 ) ;
  assign n3975 = x72 & n3757 ;
  assign n3976 = ( ~n3762 & n3974 ) | ( ~n3762 & n3975 ) | ( n3974 & n3975 ) ;
  assign n3977 = ( n3762 & n3974 ) | ( n3762 & n3975 ) | ( n3974 & n3975 ) ;
  assign n3978 = ( n3762 & n3976 ) | ( n3762 & ~n3977 ) | ( n3976 & ~n3977 ) ;
  assign n3979 = ( x73 & n3973 ) | ( x73 & ~n3978 ) | ( n3973 & ~n3978 ) ;
  assign n3980 = ( x73 & n3763 ) | ( x73 & ~n3920 ) | ( n3763 & ~n3920 ) ;
  assign n3981 = x73 & n3763 ;
  assign n3982 = ( ~n3768 & n3980 ) | ( ~n3768 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3983 = ( n3768 & n3980 ) | ( n3768 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3984 = ( n3768 & n3982 ) | ( n3768 & ~n3983 ) | ( n3982 & ~n3983 ) ;
  assign n3985 = ( x74 & n3979 ) | ( x74 & ~n3984 ) | ( n3979 & ~n3984 ) ;
  assign n3986 = ( x74 & n3769 ) | ( x74 & ~n3920 ) | ( n3769 & ~n3920 ) ;
  assign n3987 = x74 & n3769 ;
  assign n3988 = ( ~n3774 & n3986 ) | ( ~n3774 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3989 = ( n3774 & n3986 ) | ( n3774 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3990 = ( n3774 & n3988 ) | ( n3774 & ~n3989 ) | ( n3988 & ~n3989 ) ;
  assign n3991 = ( x75 & n3985 ) | ( x75 & ~n3990 ) | ( n3985 & ~n3990 ) ;
  assign n3992 = ( x75 & n3775 ) | ( x75 & ~n3920 ) | ( n3775 & ~n3920 ) ;
  assign n3993 = x75 & n3775 ;
  assign n3994 = ( ~n3780 & n3992 ) | ( ~n3780 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3995 = ( n3780 & n3992 ) | ( n3780 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3996 = ( n3780 & n3994 ) | ( n3780 & ~n3995 ) | ( n3994 & ~n3995 ) ;
  assign n3997 = ( x76 & n3991 ) | ( x76 & ~n3996 ) | ( n3991 & ~n3996 ) ;
  assign n3998 = ( x76 & n3781 ) | ( x76 & ~n3920 ) | ( n3781 & ~n3920 ) ;
  assign n3999 = x76 & n3781 ;
  assign n4000 = ( ~n3786 & n3998 ) | ( ~n3786 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4001 = ( n3786 & n3998 ) | ( n3786 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4002 = ( n3786 & n4000 ) | ( n3786 & ~n4001 ) | ( n4000 & ~n4001 ) ;
  assign n4003 = ( x77 & n3997 ) | ( x77 & ~n4002 ) | ( n3997 & ~n4002 ) ;
  assign n4004 = ( x77 & n3787 ) | ( x77 & ~n3920 ) | ( n3787 & ~n3920 ) ;
  assign n4005 = x77 & n3787 ;
  assign n4006 = ( ~n3792 & n4004 ) | ( ~n3792 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4007 = ( n3792 & n4004 ) | ( n3792 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4008 = ( n3792 & n4006 ) | ( n3792 & ~n4007 ) | ( n4006 & ~n4007 ) ;
  assign n4009 = ( x78 & n4003 ) | ( x78 & ~n4008 ) | ( n4003 & ~n4008 ) ;
  assign n4010 = ( x78 & n3793 ) | ( x78 & ~n3920 ) | ( n3793 & ~n3920 ) ;
  assign n4011 = x78 & n3793 ;
  assign n4012 = ( ~n3798 & n4010 ) | ( ~n3798 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4013 = ( n3798 & n4010 ) | ( n3798 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4014 = ( n3798 & n4012 ) | ( n3798 & ~n4013 ) | ( n4012 & ~n4013 ) ;
  assign n4015 = ( x79 & n4009 ) | ( x79 & ~n4014 ) | ( n4009 & ~n4014 ) ;
  assign n4016 = ( x79 & n3799 ) | ( x79 & ~n3920 ) | ( n3799 & ~n3920 ) ;
  assign n4017 = x79 & n3799 ;
  assign n4018 = ( ~n3804 & n4016 ) | ( ~n3804 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4019 = ( n3804 & n4016 ) | ( n3804 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4020 = ( n3804 & n4018 ) | ( n3804 & ~n4019 ) | ( n4018 & ~n4019 ) ;
  assign n4021 = ( x80 & n4015 ) | ( x80 & ~n4020 ) | ( n4015 & ~n4020 ) ;
  assign n4022 = ( x80 & n3805 ) | ( x80 & ~n3920 ) | ( n3805 & ~n3920 ) ;
  assign n4023 = x80 & n3805 ;
  assign n4024 = ( ~n3810 & n4022 ) | ( ~n3810 & n4023 ) | ( n4022 & n4023 ) ;
  assign n4025 = ( n3810 & n4022 ) | ( n3810 & n4023 ) | ( n4022 & n4023 ) ;
  assign n4026 = ( n3810 & n4024 ) | ( n3810 & ~n4025 ) | ( n4024 & ~n4025 ) ;
  assign n4027 = ( x81 & n4021 ) | ( x81 & ~n4026 ) | ( n4021 & ~n4026 ) ;
  assign n4028 = ( x81 & n3811 ) | ( x81 & ~n3920 ) | ( n3811 & ~n3920 ) ;
  assign n4029 = x81 & n3811 ;
  assign n4030 = ( ~n3816 & n4028 ) | ( ~n3816 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4031 = ( n3816 & n4028 ) | ( n3816 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4032 = ( n3816 & n4030 ) | ( n3816 & ~n4031 ) | ( n4030 & ~n4031 ) ;
  assign n4033 = ( x82 & n4027 ) | ( x82 & ~n4032 ) | ( n4027 & ~n4032 ) ;
  assign n4034 = ( x82 & n3817 ) | ( x82 & ~n3920 ) | ( n3817 & ~n3920 ) ;
  assign n4035 = x82 & n3817 ;
  assign n4036 = ( ~n3822 & n4034 ) | ( ~n3822 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4037 = ( n3822 & n4034 ) | ( n3822 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4038 = ( n3822 & n4036 ) | ( n3822 & ~n4037 ) | ( n4036 & ~n4037 ) ;
  assign n4039 = ( x83 & n4033 ) | ( x83 & ~n4038 ) | ( n4033 & ~n4038 ) ;
  assign n4040 = ( x83 & n3823 ) | ( x83 & ~n3920 ) | ( n3823 & ~n3920 ) ;
  assign n4041 = x83 & n3823 ;
  assign n4042 = ( ~n3828 & n4040 ) | ( ~n3828 & n4041 ) | ( n4040 & n4041 ) ;
  assign n4043 = ( n3828 & n4040 ) | ( n3828 & n4041 ) | ( n4040 & n4041 ) ;
  assign n4044 = ( n3828 & n4042 ) | ( n3828 & ~n4043 ) | ( n4042 & ~n4043 ) ;
  assign n4045 = ( x84 & n4039 ) | ( x84 & ~n4044 ) | ( n4039 & ~n4044 ) ;
  assign n4046 = ( x84 & n3829 ) | ( x84 & ~n3920 ) | ( n3829 & ~n3920 ) ;
  assign n4047 = x84 & n3829 ;
  assign n4048 = ( ~n3834 & n4046 ) | ( ~n3834 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4049 = ( n3834 & n4046 ) | ( n3834 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4050 = ( n3834 & n4048 ) | ( n3834 & ~n4049 ) | ( n4048 & ~n4049 ) ;
  assign n4051 = ( x85 & n4045 ) | ( x85 & ~n4050 ) | ( n4045 & ~n4050 ) ;
  assign n4052 = ( x85 & n3835 ) | ( x85 & ~n3920 ) | ( n3835 & ~n3920 ) ;
  assign n4053 = x85 & n3835 ;
  assign n4054 = ( ~n3840 & n4052 ) | ( ~n3840 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = ( n3840 & n4052 ) | ( n3840 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4056 = ( n3840 & n4054 ) | ( n3840 & ~n4055 ) | ( n4054 & ~n4055 ) ;
  assign n4057 = ( x86 & n4051 ) | ( x86 & ~n4056 ) | ( n4051 & ~n4056 ) ;
  assign n4058 = ( x86 & n3841 ) | ( x86 & ~n3920 ) | ( n3841 & ~n3920 ) ;
  assign n4059 = x86 & n3841 ;
  assign n4060 = ( ~n3846 & n4058 ) | ( ~n3846 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4061 = ( n3846 & n4058 ) | ( n3846 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4062 = ( n3846 & n4060 ) | ( n3846 & ~n4061 ) | ( n4060 & ~n4061 ) ;
  assign n4063 = ( x87 & n4057 ) | ( x87 & ~n4062 ) | ( n4057 & ~n4062 ) ;
  assign n4064 = ( x87 & n3847 ) | ( x87 & ~n3920 ) | ( n3847 & ~n3920 ) ;
  assign n4065 = x87 & n3847 ;
  assign n4066 = ( ~n3852 & n4064 ) | ( ~n3852 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4067 = ( n3852 & n4064 ) | ( n3852 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4068 = ( n3852 & n4066 ) | ( n3852 & ~n4067 ) | ( n4066 & ~n4067 ) ;
  assign n4069 = ( x88 & n4063 ) | ( x88 & ~n4068 ) | ( n4063 & ~n4068 ) ;
  assign n4070 = ( x88 & n3853 ) | ( x88 & ~n3920 ) | ( n3853 & ~n3920 ) ;
  assign n4071 = x88 & n3853 ;
  assign n4072 = ( ~n3858 & n4070 ) | ( ~n3858 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4073 = ( n3858 & n4070 ) | ( n3858 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4074 = ( n3858 & n4072 ) | ( n3858 & ~n4073 ) | ( n4072 & ~n4073 ) ;
  assign n4075 = ( x89 & n4069 ) | ( x89 & ~n4074 ) | ( n4069 & ~n4074 ) ;
  assign n4076 = ( x89 & n3859 ) | ( x89 & ~n3920 ) | ( n3859 & ~n3920 ) ;
  assign n4077 = x89 & n3859 ;
  assign n4078 = ( ~n3864 & n4076 ) | ( ~n3864 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4079 = ( n3864 & n4076 ) | ( n3864 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4080 = ( n3864 & n4078 ) | ( n3864 & ~n4079 ) | ( n4078 & ~n4079 ) ;
  assign n4081 = ( x90 & n4075 ) | ( x90 & ~n4080 ) | ( n4075 & ~n4080 ) ;
  assign n4082 = ( x90 & n3865 ) | ( x90 & ~n3920 ) | ( n3865 & ~n3920 ) ;
  assign n4083 = x90 & n3865 ;
  assign n4084 = ( ~n3870 & n4082 ) | ( ~n3870 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4085 = ( n3870 & n4082 ) | ( n3870 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4086 = ( n3870 & n4084 ) | ( n3870 & ~n4085 ) | ( n4084 & ~n4085 ) ;
  assign n4087 = ( x91 & n4081 ) | ( x91 & ~n4086 ) | ( n4081 & ~n4086 ) ;
  assign n4088 = ( x91 & n3871 ) | ( x91 & ~n3920 ) | ( n3871 & ~n3920 ) ;
  assign n4089 = x91 & n3871 ;
  assign n4090 = ( ~n3876 & n4088 ) | ( ~n3876 & n4089 ) | ( n4088 & n4089 ) ;
  assign n4091 = ( n3876 & n4088 ) | ( n3876 & n4089 ) | ( n4088 & n4089 ) ;
  assign n4092 = ( n3876 & n4090 ) | ( n3876 & ~n4091 ) | ( n4090 & ~n4091 ) ;
  assign n4093 = ( x92 & n4087 ) | ( x92 & ~n4092 ) | ( n4087 & ~n4092 ) ;
  assign n4094 = ( x92 & n3877 ) | ( x92 & ~n3920 ) | ( n3877 & ~n3920 ) ;
  assign n4095 = x92 & n3877 ;
  assign n4096 = ( ~n3882 & n4094 ) | ( ~n3882 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4097 = ( n3882 & n4094 ) | ( n3882 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4098 = ( n3882 & n4096 ) | ( n3882 & ~n4097 ) | ( n4096 & ~n4097 ) ;
  assign n4099 = ( x93 & n4093 ) | ( x93 & ~n4098 ) | ( n4093 & ~n4098 ) ;
  assign n4100 = ( x93 & n3883 ) | ( x93 & ~n3920 ) | ( n3883 & ~n3920 ) ;
  assign n4101 = x93 & n3883 ;
  assign n4102 = ( ~n3888 & n4100 ) | ( ~n3888 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = ( n3888 & n4100 ) | ( n3888 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4104 = ( n3888 & n4102 ) | ( n3888 & ~n4103 ) | ( n4102 & ~n4103 ) ;
  assign n4105 = ( x94 & n4099 ) | ( x94 & ~n4104 ) | ( n4099 & ~n4104 ) ;
  assign n4106 = ( x94 & n3889 ) | ( x94 & ~n3920 ) | ( n3889 & ~n3920 ) ;
  assign n4107 = x94 & n3889 ;
  assign n4108 = ( ~n3894 & n4106 ) | ( ~n3894 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = ( n3894 & n4106 ) | ( n3894 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4110 = ( n3894 & n4108 ) | ( n3894 & ~n4109 ) | ( n4108 & ~n4109 ) ;
  assign n4111 = ( x95 & n4105 ) | ( x95 & ~n4110 ) | ( n4105 & ~n4110 ) ;
  assign n4112 = ( x95 & n3895 ) | ( x95 & ~n3920 ) | ( n3895 & ~n3920 ) ;
  assign n4113 = x95 & n3895 ;
  assign n4114 = ( ~n3900 & n4112 ) | ( ~n3900 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n3900 & n4112 ) | ( n3900 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4116 = ( n3900 & n4114 ) | ( n3900 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = ( x96 & n4111 ) | ( x96 & ~n4116 ) | ( n4111 & ~n4116 ) ;
  assign n4118 = ( x96 & n3901 ) | ( x96 & ~n3920 ) | ( n3901 & ~n3920 ) ;
  assign n4119 = x96 & n3901 ;
  assign n4120 = ( ~n3906 & n4118 ) | ( ~n3906 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4121 = ( n3906 & n4118 ) | ( n3906 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4122 = ( n3906 & n4120 ) | ( n3906 & ~n4121 ) | ( n4120 & ~n4121 ) ;
  assign n4123 = ( x97 & n4117 ) | ( x97 & ~n4122 ) | ( n4117 & ~n4122 ) ;
  assign n4124 = ( x97 & n3907 ) | ( x97 & ~n3920 ) | ( n3907 & ~n3920 ) ;
  assign n4125 = x97 & n3907 ;
  assign n4126 = ( ~n3912 & n4124 ) | ( ~n3912 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = ( n3912 & n4124 ) | ( n3912 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4128 = ( n3912 & n4126 ) | ( n3912 & ~n4127 ) | ( n4126 & ~n4127 ) ;
  assign n4129 = ( x98 & n4123 ) | ( x98 & ~n4128 ) | ( n4123 & ~n4128 ) ;
  assign n4130 = ( x99 & ~n3925 ) | ( x99 & n4129 ) | ( ~n3925 & n4129 ) ;
  assign n4131 = ( n158 & n389 ) | ( n158 & n3507 ) | ( n389 & n3507 ) ;
  assign n4132 = ( n389 & n3918 ) | ( n389 & n4131 ) | ( n3918 & n4131 ) ;
  assign n4133 = ( x100 & n4130 ) | ( x100 & ~n4132 ) | ( n4130 & ~n4132 ) ;
  assign n4134 = n156 | n4133 ;
  assign n4135 = ( x99 & n4129 ) | ( x99 & n4134 ) | ( n4129 & n4134 ) ;
  assign n4136 = x99 | n4129 ;
  assign n4137 = ( ~n3925 & n4135 ) | ( ~n3925 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4138 = ( n3925 & n4135 ) | ( n3925 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4139 = ( n3925 & n4137 ) | ( n3925 & ~n4138 ) | ( n4137 & ~n4138 ) ;
  assign n4140 = ~x26 & x64 ;
  assign n4141 = ~x27 & n4134 ;
  assign n4142 = ( x27 & ~x64 ) | ( x27 & n4134 ) | ( ~x64 & n4134 ) ;
  assign n4143 = ( n3926 & ~n4141 ) | ( n3926 & n4142 ) | ( ~n4141 & n4142 ) ;
  assign n4144 = ( x65 & n4140 ) | ( x65 & ~n4143 ) | ( n4140 & ~n4143 ) ;
  assign n4145 = ( x65 & n3926 ) | ( x65 & n4134 ) | ( n3926 & n4134 ) ;
  assign n4146 = x65 | n3926 ;
  assign n4147 = ( ~n3930 & n4145 ) | ( ~n3930 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( n3930 & n4145 ) | ( n3930 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4149 = ( n3930 & n4147 ) | ( n3930 & ~n4148 ) | ( n4147 & ~n4148 ) ;
  assign n4150 = ( x66 & n4144 ) | ( x66 & ~n4149 ) | ( n4144 & ~n4149 ) ;
  assign n4151 = ( x66 & n3931 ) | ( x66 & n4134 ) | ( n3931 & n4134 ) ;
  assign n4152 = x66 | n3931 ;
  assign n4153 = ( ~n3936 & n4151 ) | ( ~n3936 & n4152 ) | ( n4151 & n4152 ) ;
  assign n4154 = ( n3936 & n4151 ) | ( n3936 & n4152 ) | ( n4151 & n4152 ) ;
  assign n4155 = ( n3936 & n4153 ) | ( n3936 & ~n4154 ) | ( n4153 & ~n4154 ) ;
  assign n4156 = ( x67 & n4150 ) | ( x67 & ~n4155 ) | ( n4150 & ~n4155 ) ;
  assign n4157 = ( x67 & n3937 ) | ( x67 & ~n4134 ) | ( n3937 & ~n4134 ) ;
  assign n4158 = x67 & n3937 ;
  assign n4159 = ( ~n3942 & n4157 ) | ( ~n3942 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4160 = ( n3942 & n4157 ) | ( n3942 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4161 = ( n3942 & n4159 ) | ( n3942 & ~n4160 ) | ( n4159 & ~n4160 ) ;
  assign n4162 = ( x68 & n4156 ) | ( x68 & ~n4161 ) | ( n4156 & ~n4161 ) ;
  assign n4163 = ( x68 & n3943 ) | ( x68 & ~n4134 ) | ( n3943 & ~n4134 ) ;
  assign n4164 = x68 & n3943 ;
  assign n4165 = ( ~n3948 & n4163 ) | ( ~n3948 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4166 = ( n3948 & n4163 ) | ( n3948 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4167 = ( n3948 & n4165 ) | ( n3948 & ~n4166 ) | ( n4165 & ~n4166 ) ;
  assign n4168 = ( x69 & n4162 ) | ( x69 & ~n4167 ) | ( n4162 & ~n4167 ) ;
  assign n4169 = ( x69 & n3949 ) | ( x69 & ~n4134 ) | ( n3949 & ~n4134 ) ;
  assign n4170 = x69 & n3949 ;
  assign n4171 = ( ~n3954 & n4169 ) | ( ~n3954 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4172 = ( n3954 & n4169 ) | ( n3954 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4173 = ( n3954 & n4171 ) | ( n3954 & ~n4172 ) | ( n4171 & ~n4172 ) ;
  assign n4174 = ( x70 & n4168 ) | ( x70 & ~n4173 ) | ( n4168 & ~n4173 ) ;
  assign n4175 = ( x70 & n3955 ) | ( x70 & ~n4134 ) | ( n3955 & ~n4134 ) ;
  assign n4176 = x70 & n3955 ;
  assign n4177 = ( ~n3960 & n4175 ) | ( ~n3960 & n4176 ) | ( n4175 & n4176 ) ;
  assign n4178 = ( n3960 & n4175 ) | ( n3960 & n4176 ) | ( n4175 & n4176 ) ;
  assign n4179 = ( n3960 & n4177 ) | ( n3960 & ~n4178 ) | ( n4177 & ~n4178 ) ;
  assign n4180 = ( x71 & n4174 ) | ( x71 & ~n4179 ) | ( n4174 & ~n4179 ) ;
  assign n4181 = ( x71 & n3961 ) | ( x71 & ~n4134 ) | ( n3961 & ~n4134 ) ;
  assign n4182 = x71 & n3961 ;
  assign n4183 = ( ~n3966 & n4181 ) | ( ~n3966 & n4182 ) | ( n4181 & n4182 ) ;
  assign n4184 = ( n3966 & n4181 ) | ( n3966 & n4182 ) | ( n4181 & n4182 ) ;
  assign n4185 = ( n3966 & n4183 ) | ( n3966 & ~n4184 ) | ( n4183 & ~n4184 ) ;
  assign n4186 = ( x72 & n4180 ) | ( x72 & ~n4185 ) | ( n4180 & ~n4185 ) ;
  assign n4187 = ( x72 & n3967 ) | ( x72 & ~n4134 ) | ( n3967 & ~n4134 ) ;
  assign n4188 = x72 & n3967 ;
  assign n4189 = ( ~n3972 & n4187 ) | ( ~n3972 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = ( n3972 & n4187 ) | ( n3972 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4191 = ( n3972 & n4189 ) | ( n3972 & ~n4190 ) | ( n4189 & ~n4190 ) ;
  assign n4192 = ( x73 & n4186 ) | ( x73 & ~n4191 ) | ( n4186 & ~n4191 ) ;
  assign n4193 = ( x73 & n3973 ) | ( x73 & ~n4134 ) | ( n3973 & ~n4134 ) ;
  assign n4194 = x73 & n3973 ;
  assign n4195 = ( ~n3978 & n4193 ) | ( ~n3978 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = ( n3978 & n4193 ) | ( n3978 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4197 = ( n3978 & n4195 ) | ( n3978 & ~n4196 ) | ( n4195 & ~n4196 ) ;
  assign n4198 = ( x74 & n4192 ) | ( x74 & ~n4197 ) | ( n4192 & ~n4197 ) ;
  assign n4199 = ( x74 & n3979 ) | ( x74 & ~n4134 ) | ( n3979 & ~n4134 ) ;
  assign n4200 = x74 & n3979 ;
  assign n4201 = ( ~n3984 & n4199 ) | ( ~n3984 & n4200 ) | ( n4199 & n4200 ) ;
  assign n4202 = ( n3984 & n4199 ) | ( n3984 & n4200 ) | ( n4199 & n4200 ) ;
  assign n4203 = ( n3984 & n4201 ) | ( n3984 & ~n4202 ) | ( n4201 & ~n4202 ) ;
  assign n4204 = ( x75 & n4198 ) | ( x75 & ~n4203 ) | ( n4198 & ~n4203 ) ;
  assign n4205 = ( x75 & n3985 ) | ( x75 & ~n4134 ) | ( n3985 & ~n4134 ) ;
  assign n4206 = x75 & n3985 ;
  assign n4207 = ( ~n3990 & n4205 ) | ( ~n3990 & n4206 ) | ( n4205 & n4206 ) ;
  assign n4208 = ( n3990 & n4205 ) | ( n3990 & n4206 ) | ( n4205 & n4206 ) ;
  assign n4209 = ( n3990 & n4207 ) | ( n3990 & ~n4208 ) | ( n4207 & ~n4208 ) ;
  assign n4210 = ( x76 & n4204 ) | ( x76 & ~n4209 ) | ( n4204 & ~n4209 ) ;
  assign n4211 = ( x76 & n3991 ) | ( x76 & ~n4134 ) | ( n3991 & ~n4134 ) ;
  assign n4212 = x76 & n3991 ;
  assign n4213 = ( ~n3996 & n4211 ) | ( ~n3996 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4214 = ( n3996 & n4211 ) | ( n3996 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4215 = ( n3996 & n4213 ) | ( n3996 & ~n4214 ) | ( n4213 & ~n4214 ) ;
  assign n4216 = ( x77 & n4210 ) | ( x77 & ~n4215 ) | ( n4210 & ~n4215 ) ;
  assign n4217 = ( x77 & n3997 ) | ( x77 & ~n4134 ) | ( n3997 & ~n4134 ) ;
  assign n4218 = x77 & n3997 ;
  assign n4219 = ( ~n4002 & n4217 ) | ( ~n4002 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4220 = ( n4002 & n4217 ) | ( n4002 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4221 = ( n4002 & n4219 ) | ( n4002 & ~n4220 ) | ( n4219 & ~n4220 ) ;
  assign n4222 = ( x78 & n4216 ) | ( x78 & ~n4221 ) | ( n4216 & ~n4221 ) ;
  assign n4223 = ( x78 & n4003 ) | ( x78 & ~n4134 ) | ( n4003 & ~n4134 ) ;
  assign n4224 = x78 & n4003 ;
  assign n4225 = ( ~n4008 & n4223 ) | ( ~n4008 & n4224 ) | ( n4223 & n4224 ) ;
  assign n4226 = ( n4008 & n4223 ) | ( n4008 & n4224 ) | ( n4223 & n4224 ) ;
  assign n4227 = ( n4008 & n4225 ) | ( n4008 & ~n4226 ) | ( n4225 & ~n4226 ) ;
  assign n4228 = ( x79 & n4222 ) | ( x79 & ~n4227 ) | ( n4222 & ~n4227 ) ;
  assign n4229 = ( x79 & n4009 ) | ( x79 & ~n4134 ) | ( n4009 & ~n4134 ) ;
  assign n4230 = x79 & n4009 ;
  assign n4231 = ( ~n4014 & n4229 ) | ( ~n4014 & n4230 ) | ( n4229 & n4230 ) ;
  assign n4232 = ( n4014 & n4229 ) | ( n4014 & n4230 ) | ( n4229 & n4230 ) ;
  assign n4233 = ( n4014 & n4231 ) | ( n4014 & ~n4232 ) | ( n4231 & ~n4232 ) ;
  assign n4234 = ( x80 & n4228 ) | ( x80 & ~n4233 ) | ( n4228 & ~n4233 ) ;
  assign n4235 = ( x80 & n4015 ) | ( x80 & ~n4134 ) | ( n4015 & ~n4134 ) ;
  assign n4236 = x80 & n4015 ;
  assign n4237 = ( ~n4020 & n4235 ) | ( ~n4020 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4238 = ( n4020 & n4235 ) | ( n4020 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4239 = ( n4020 & n4237 ) | ( n4020 & ~n4238 ) | ( n4237 & ~n4238 ) ;
  assign n4240 = ( x81 & n4234 ) | ( x81 & ~n4239 ) | ( n4234 & ~n4239 ) ;
  assign n4241 = ( x81 & n4021 ) | ( x81 & ~n4134 ) | ( n4021 & ~n4134 ) ;
  assign n4242 = x81 & n4021 ;
  assign n4243 = ( ~n4026 & n4241 ) | ( ~n4026 & n4242 ) | ( n4241 & n4242 ) ;
  assign n4244 = ( n4026 & n4241 ) | ( n4026 & n4242 ) | ( n4241 & n4242 ) ;
  assign n4245 = ( n4026 & n4243 ) | ( n4026 & ~n4244 ) | ( n4243 & ~n4244 ) ;
  assign n4246 = ( x82 & n4240 ) | ( x82 & ~n4245 ) | ( n4240 & ~n4245 ) ;
  assign n4247 = ( x82 & n4027 ) | ( x82 & ~n4134 ) | ( n4027 & ~n4134 ) ;
  assign n4248 = x82 & n4027 ;
  assign n4249 = ( ~n4032 & n4247 ) | ( ~n4032 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4250 = ( n4032 & n4247 ) | ( n4032 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4251 = ( n4032 & n4249 ) | ( n4032 & ~n4250 ) | ( n4249 & ~n4250 ) ;
  assign n4252 = ( x83 & n4246 ) | ( x83 & ~n4251 ) | ( n4246 & ~n4251 ) ;
  assign n4253 = ( x83 & n4033 ) | ( x83 & ~n4134 ) | ( n4033 & ~n4134 ) ;
  assign n4254 = x83 & n4033 ;
  assign n4255 = ( ~n4038 & n4253 ) | ( ~n4038 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4256 = ( n4038 & n4253 ) | ( n4038 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4257 = ( n4038 & n4255 ) | ( n4038 & ~n4256 ) | ( n4255 & ~n4256 ) ;
  assign n4258 = ( x84 & n4252 ) | ( x84 & ~n4257 ) | ( n4252 & ~n4257 ) ;
  assign n4259 = ( x84 & n4039 ) | ( x84 & ~n4134 ) | ( n4039 & ~n4134 ) ;
  assign n4260 = x84 & n4039 ;
  assign n4261 = ( ~n4044 & n4259 ) | ( ~n4044 & n4260 ) | ( n4259 & n4260 ) ;
  assign n4262 = ( n4044 & n4259 ) | ( n4044 & n4260 ) | ( n4259 & n4260 ) ;
  assign n4263 = ( n4044 & n4261 ) | ( n4044 & ~n4262 ) | ( n4261 & ~n4262 ) ;
  assign n4264 = ( x85 & n4258 ) | ( x85 & ~n4263 ) | ( n4258 & ~n4263 ) ;
  assign n4265 = ( x85 & n4045 ) | ( x85 & ~n4134 ) | ( n4045 & ~n4134 ) ;
  assign n4266 = x85 & n4045 ;
  assign n4267 = ( ~n4050 & n4265 ) | ( ~n4050 & n4266 ) | ( n4265 & n4266 ) ;
  assign n4268 = ( n4050 & n4265 ) | ( n4050 & n4266 ) | ( n4265 & n4266 ) ;
  assign n4269 = ( n4050 & n4267 ) | ( n4050 & ~n4268 ) | ( n4267 & ~n4268 ) ;
  assign n4270 = ( x86 & n4264 ) | ( x86 & ~n4269 ) | ( n4264 & ~n4269 ) ;
  assign n4271 = ( x86 & n4051 ) | ( x86 & ~n4134 ) | ( n4051 & ~n4134 ) ;
  assign n4272 = x86 & n4051 ;
  assign n4273 = ( ~n4056 & n4271 ) | ( ~n4056 & n4272 ) | ( n4271 & n4272 ) ;
  assign n4274 = ( n4056 & n4271 ) | ( n4056 & n4272 ) | ( n4271 & n4272 ) ;
  assign n4275 = ( n4056 & n4273 ) | ( n4056 & ~n4274 ) | ( n4273 & ~n4274 ) ;
  assign n4276 = ( x87 & n4270 ) | ( x87 & ~n4275 ) | ( n4270 & ~n4275 ) ;
  assign n4277 = ( x87 & n4057 ) | ( x87 & ~n4134 ) | ( n4057 & ~n4134 ) ;
  assign n4278 = x87 & n4057 ;
  assign n4279 = ( ~n4062 & n4277 ) | ( ~n4062 & n4278 ) | ( n4277 & n4278 ) ;
  assign n4280 = ( n4062 & n4277 ) | ( n4062 & n4278 ) | ( n4277 & n4278 ) ;
  assign n4281 = ( n4062 & n4279 ) | ( n4062 & ~n4280 ) | ( n4279 & ~n4280 ) ;
  assign n4282 = ( x88 & n4276 ) | ( x88 & ~n4281 ) | ( n4276 & ~n4281 ) ;
  assign n4283 = ( x88 & n4063 ) | ( x88 & ~n4134 ) | ( n4063 & ~n4134 ) ;
  assign n4284 = x88 & n4063 ;
  assign n4285 = ( ~n4068 & n4283 ) | ( ~n4068 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4286 = ( n4068 & n4283 ) | ( n4068 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4287 = ( n4068 & n4285 ) | ( n4068 & ~n4286 ) | ( n4285 & ~n4286 ) ;
  assign n4288 = ( x89 & n4282 ) | ( x89 & ~n4287 ) | ( n4282 & ~n4287 ) ;
  assign n4289 = ( x89 & n4069 ) | ( x89 & ~n4134 ) | ( n4069 & ~n4134 ) ;
  assign n4290 = x89 & n4069 ;
  assign n4291 = ( ~n4074 & n4289 ) | ( ~n4074 & n4290 ) | ( n4289 & n4290 ) ;
  assign n4292 = ( n4074 & n4289 ) | ( n4074 & n4290 ) | ( n4289 & n4290 ) ;
  assign n4293 = ( n4074 & n4291 ) | ( n4074 & ~n4292 ) | ( n4291 & ~n4292 ) ;
  assign n4294 = ( x90 & n4288 ) | ( x90 & ~n4293 ) | ( n4288 & ~n4293 ) ;
  assign n4295 = ( x90 & n4075 ) | ( x90 & ~n4134 ) | ( n4075 & ~n4134 ) ;
  assign n4296 = x90 & n4075 ;
  assign n4297 = ( ~n4080 & n4295 ) | ( ~n4080 & n4296 ) | ( n4295 & n4296 ) ;
  assign n4298 = ( n4080 & n4295 ) | ( n4080 & n4296 ) | ( n4295 & n4296 ) ;
  assign n4299 = ( n4080 & n4297 ) | ( n4080 & ~n4298 ) | ( n4297 & ~n4298 ) ;
  assign n4300 = ( x91 & n4294 ) | ( x91 & ~n4299 ) | ( n4294 & ~n4299 ) ;
  assign n4301 = ( x91 & n4081 ) | ( x91 & ~n4134 ) | ( n4081 & ~n4134 ) ;
  assign n4302 = x91 & n4081 ;
  assign n4303 = ( ~n4086 & n4301 ) | ( ~n4086 & n4302 ) | ( n4301 & n4302 ) ;
  assign n4304 = ( n4086 & n4301 ) | ( n4086 & n4302 ) | ( n4301 & n4302 ) ;
  assign n4305 = ( n4086 & n4303 ) | ( n4086 & ~n4304 ) | ( n4303 & ~n4304 ) ;
  assign n4306 = ( x92 & n4300 ) | ( x92 & ~n4305 ) | ( n4300 & ~n4305 ) ;
  assign n4307 = ( x92 & n4087 ) | ( x92 & ~n4134 ) | ( n4087 & ~n4134 ) ;
  assign n4308 = x92 & n4087 ;
  assign n4309 = ( ~n4092 & n4307 ) | ( ~n4092 & n4308 ) | ( n4307 & n4308 ) ;
  assign n4310 = ( n4092 & n4307 ) | ( n4092 & n4308 ) | ( n4307 & n4308 ) ;
  assign n4311 = ( n4092 & n4309 ) | ( n4092 & ~n4310 ) | ( n4309 & ~n4310 ) ;
  assign n4312 = ( x93 & n4306 ) | ( x93 & ~n4311 ) | ( n4306 & ~n4311 ) ;
  assign n4313 = ( x93 & n4093 ) | ( x93 & ~n4134 ) | ( n4093 & ~n4134 ) ;
  assign n4314 = x93 & n4093 ;
  assign n4315 = ( ~n4098 & n4313 ) | ( ~n4098 & n4314 ) | ( n4313 & n4314 ) ;
  assign n4316 = ( n4098 & n4313 ) | ( n4098 & n4314 ) | ( n4313 & n4314 ) ;
  assign n4317 = ( n4098 & n4315 ) | ( n4098 & ~n4316 ) | ( n4315 & ~n4316 ) ;
  assign n4318 = ( x94 & n4312 ) | ( x94 & ~n4317 ) | ( n4312 & ~n4317 ) ;
  assign n4319 = ( x94 & n4099 ) | ( x94 & ~n4134 ) | ( n4099 & ~n4134 ) ;
  assign n4320 = x94 & n4099 ;
  assign n4321 = ( ~n4104 & n4319 ) | ( ~n4104 & n4320 ) | ( n4319 & n4320 ) ;
  assign n4322 = ( n4104 & n4319 ) | ( n4104 & n4320 ) | ( n4319 & n4320 ) ;
  assign n4323 = ( n4104 & n4321 ) | ( n4104 & ~n4322 ) | ( n4321 & ~n4322 ) ;
  assign n4324 = ( x95 & n4318 ) | ( x95 & ~n4323 ) | ( n4318 & ~n4323 ) ;
  assign n4325 = ( x95 & n4105 ) | ( x95 & ~n4134 ) | ( n4105 & ~n4134 ) ;
  assign n4326 = x95 & n4105 ;
  assign n4327 = ( ~n4110 & n4325 ) | ( ~n4110 & n4326 ) | ( n4325 & n4326 ) ;
  assign n4328 = ( n4110 & n4325 ) | ( n4110 & n4326 ) | ( n4325 & n4326 ) ;
  assign n4329 = ( n4110 & n4327 ) | ( n4110 & ~n4328 ) | ( n4327 & ~n4328 ) ;
  assign n4330 = ( x96 & n4324 ) | ( x96 & ~n4329 ) | ( n4324 & ~n4329 ) ;
  assign n4331 = ( x96 & n4111 ) | ( x96 & ~n4134 ) | ( n4111 & ~n4134 ) ;
  assign n4332 = x96 & n4111 ;
  assign n4333 = ( ~n4116 & n4331 ) | ( ~n4116 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4334 = ( n4116 & n4331 ) | ( n4116 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4335 = ( n4116 & n4333 ) | ( n4116 & ~n4334 ) | ( n4333 & ~n4334 ) ;
  assign n4336 = ( x97 & n4330 ) | ( x97 & ~n4335 ) | ( n4330 & ~n4335 ) ;
  assign n4337 = ( x97 & n4117 ) | ( x97 & ~n4134 ) | ( n4117 & ~n4134 ) ;
  assign n4338 = x97 & n4117 ;
  assign n4339 = ( ~n4122 & n4337 ) | ( ~n4122 & n4338 ) | ( n4337 & n4338 ) ;
  assign n4340 = ( n4122 & n4337 ) | ( n4122 & n4338 ) | ( n4337 & n4338 ) ;
  assign n4341 = ( n4122 & n4339 ) | ( n4122 & ~n4340 ) | ( n4339 & ~n4340 ) ;
  assign n4342 = ( x98 & n4336 ) | ( x98 & ~n4341 ) | ( n4336 & ~n4341 ) ;
  assign n4343 = ( x98 & n4123 ) | ( x98 & ~n4134 ) | ( n4123 & ~n4134 ) ;
  assign n4344 = x98 & n4123 ;
  assign n4345 = ( ~n4128 & n4343 ) | ( ~n4128 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = ( n4128 & n4343 ) | ( n4128 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4347 = ( n4128 & n4345 ) | ( n4128 & ~n4346 ) | ( n4345 & ~n4346 ) ;
  assign n4348 = ( x99 & n4342 ) | ( x99 & ~n4347 ) | ( n4342 & ~n4347 ) ;
  assign n4349 = ( x100 & n156 ) | ( x100 & n4130 ) | ( n156 & n4130 ) ;
  assign n4350 = x100 | n4130 ;
  assign n4351 = ( n4132 & n4349 ) | ( n4132 & ~n4350 ) | ( n4349 & ~n4350 ) ;
  assign n4352 = ( x100 & ~n4139 ) | ( x100 & n4348 ) | ( ~n4139 & n4348 ) ;
  assign n4353 = ( x101 & ~n4351 ) | ( x101 & n4352 ) | ( ~n4351 & n4352 ) ;
  assign n4354 = n155 | n4353 ;
  assign n4355 = ( x100 & n4348 ) | ( x100 & n4354 ) | ( n4348 & n4354 ) ;
  assign n4356 = x100 | n4348 ;
  assign n4357 = ( ~n4139 & n4355 ) | ( ~n4139 & n4356 ) | ( n4355 & n4356 ) ;
  assign n4358 = ( n4139 & n4355 ) | ( n4139 & n4356 ) | ( n4355 & n4356 ) ;
  assign n4359 = ( n4139 & n4357 ) | ( n4139 & ~n4358 ) | ( n4357 & ~n4358 ) ;
  assign n4360 = ~x25 & x64 ;
  assign n4361 = ~x26 & n4354 ;
  assign n4362 = ( x26 & ~x64 ) | ( x26 & n4354 ) | ( ~x64 & n4354 ) ;
  assign n4363 = ( n4140 & ~n4361 ) | ( n4140 & n4362 ) | ( ~n4361 & n4362 ) ;
  assign n4364 = ( x65 & n4360 ) | ( x65 & ~n4363 ) | ( n4360 & ~n4363 ) ;
  assign n4365 = ( x65 & n4140 ) | ( x65 & n4354 ) | ( n4140 & n4354 ) ;
  assign n4366 = x65 | n4140 ;
  assign n4367 = ( ~n4143 & n4365 ) | ( ~n4143 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4368 = ( n4143 & n4365 ) | ( n4143 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4369 = ( n4143 & n4367 ) | ( n4143 & ~n4368 ) | ( n4367 & ~n4368 ) ;
  assign n4370 = ( x66 & n4364 ) | ( x66 & ~n4369 ) | ( n4364 & ~n4369 ) ;
  assign n4371 = ( x66 & n4144 ) | ( x66 & n4354 ) | ( n4144 & n4354 ) ;
  assign n4372 = x66 | n4144 ;
  assign n4373 = ( ~n4149 & n4371 ) | ( ~n4149 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4374 = ( n4149 & n4371 ) | ( n4149 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4375 = ( n4149 & n4373 ) | ( n4149 & ~n4374 ) | ( n4373 & ~n4374 ) ;
  assign n4376 = ( x67 & n4370 ) | ( x67 & ~n4375 ) | ( n4370 & ~n4375 ) ;
  assign n4377 = ( x67 & n4150 ) | ( x67 & ~n4354 ) | ( n4150 & ~n4354 ) ;
  assign n4378 = x67 & n4150 ;
  assign n4379 = ( ~n4155 & n4377 ) | ( ~n4155 & n4378 ) | ( n4377 & n4378 ) ;
  assign n4380 = ( n4155 & n4377 ) | ( n4155 & n4378 ) | ( n4377 & n4378 ) ;
  assign n4381 = ( n4155 & n4379 ) | ( n4155 & ~n4380 ) | ( n4379 & ~n4380 ) ;
  assign n4382 = ( x68 & n4376 ) | ( x68 & ~n4381 ) | ( n4376 & ~n4381 ) ;
  assign n4383 = ( x68 & n4156 ) | ( x68 & ~n4354 ) | ( n4156 & ~n4354 ) ;
  assign n4384 = x68 & n4156 ;
  assign n4385 = ( ~n4161 & n4383 ) | ( ~n4161 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4386 = ( n4161 & n4383 ) | ( n4161 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4387 = ( n4161 & n4385 ) | ( n4161 & ~n4386 ) | ( n4385 & ~n4386 ) ;
  assign n4388 = ( x69 & n4382 ) | ( x69 & ~n4387 ) | ( n4382 & ~n4387 ) ;
  assign n4389 = ( x69 & n4162 ) | ( x69 & ~n4354 ) | ( n4162 & ~n4354 ) ;
  assign n4390 = x69 & n4162 ;
  assign n4391 = ( ~n4167 & n4389 ) | ( ~n4167 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4392 = ( n4167 & n4389 ) | ( n4167 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4393 = ( n4167 & n4391 ) | ( n4167 & ~n4392 ) | ( n4391 & ~n4392 ) ;
  assign n4394 = ( x70 & n4388 ) | ( x70 & ~n4393 ) | ( n4388 & ~n4393 ) ;
  assign n4395 = ( x70 & n4168 ) | ( x70 & ~n4354 ) | ( n4168 & ~n4354 ) ;
  assign n4396 = x70 & n4168 ;
  assign n4397 = ( ~n4173 & n4395 ) | ( ~n4173 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = ( n4173 & n4395 ) | ( n4173 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4399 = ( n4173 & n4397 ) | ( n4173 & ~n4398 ) | ( n4397 & ~n4398 ) ;
  assign n4400 = ( x71 & n4394 ) | ( x71 & ~n4399 ) | ( n4394 & ~n4399 ) ;
  assign n4401 = ( x71 & n4174 ) | ( x71 & ~n4354 ) | ( n4174 & ~n4354 ) ;
  assign n4402 = x71 & n4174 ;
  assign n4403 = ( ~n4179 & n4401 ) | ( ~n4179 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4404 = ( n4179 & n4401 ) | ( n4179 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4405 = ( n4179 & n4403 ) | ( n4179 & ~n4404 ) | ( n4403 & ~n4404 ) ;
  assign n4406 = ( x72 & n4400 ) | ( x72 & ~n4405 ) | ( n4400 & ~n4405 ) ;
  assign n4407 = ( x72 & n4180 ) | ( x72 & ~n4354 ) | ( n4180 & ~n4354 ) ;
  assign n4408 = x72 & n4180 ;
  assign n4409 = ( ~n4185 & n4407 ) | ( ~n4185 & n4408 ) | ( n4407 & n4408 ) ;
  assign n4410 = ( n4185 & n4407 ) | ( n4185 & n4408 ) | ( n4407 & n4408 ) ;
  assign n4411 = ( n4185 & n4409 ) | ( n4185 & ~n4410 ) | ( n4409 & ~n4410 ) ;
  assign n4412 = ( x73 & n4406 ) | ( x73 & ~n4411 ) | ( n4406 & ~n4411 ) ;
  assign n4413 = ( x73 & n4186 ) | ( x73 & ~n4354 ) | ( n4186 & ~n4354 ) ;
  assign n4414 = x73 & n4186 ;
  assign n4415 = ( ~n4191 & n4413 ) | ( ~n4191 & n4414 ) | ( n4413 & n4414 ) ;
  assign n4416 = ( n4191 & n4413 ) | ( n4191 & n4414 ) | ( n4413 & n4414 ) ;
  assign n4417 = ( n4191 & n4415 ) | ( n4191 & ~n4416 ) | ( n4415 & ~n4416 ) ;
  assign n4418 = ( x74 & n4412 ) | ( x74 & ~n4417 ) | ( n4412 & ~n4417 ) ;
  assign n4419 = ( x74 & n4192 ) | ( x74 & ~n4354 ) | ( n4192 & ~n4354 ) ;
  assign n4420 = x74 & n4192 ;
  assign n4421 = ( ~n4197 & n4419 ) | ( ~n4197 & n4420 ) | ( n4419 & n4420 ) ;
  assign n4422 = ( n4197 & n4419 ) | ( n4197 & n4420 ) | ( n4419 & n4420 ) ;
  assign n4423 = ( n4197 & n4421 ) | ( n4197 & ~n4422 ) | ( n4421 & ~n4422 ) ;
  assign n4424 = ( x75 & n4418 ) | ( x75 & ~n4423 ) | ( n4418 & ~n4423 ) ;
  assign n4425 = ( x75 & n4198 ) | ( x75 & ~n4354 ) | ( n4198 & ~n4354 ) ;
  assign n4426 = x75 & n4198 ;
  assign n4427 = ( ~n4203 & n4425 ) | ( ~n4203 & n4426 ) | ( n4425 & n4426 ) ;
  assign n4428 = ( n4203 & n4425 ) | ( n4203 & n4426 ) | ( n4425 & n4426 ) ;
  assign n4429 = ( n4203 & n4427 ) | ( n4203 & ~n4428 ) | ( n4427 & ~n4428 ) ;
  assign n4430 = ( x76 & n4424 ) | ( x76 & ~n4429 ) | ( n4424 & ~n4429 ) ;
  assign n4431 = ( x76 & n4204 ) | ( x76 & ~n4354 ) | ( n4204 & ~n4354 ) ;
  assign n4432 = x76 & n4204 ;
  assign n4433 = ( ~n4209 & n4431 ) | ( ~n4209 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4434 = ( n4209 & n4431 ) | ( n4209 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4435 = ( n4209 & n4433 ) | ( n4209 & ~n4434 ) | ( n4433 & ~n4434 ) ;
  assign n4436 = ( x77 & n4430 ) | ( x77 & ~n4435 ) | ( n4430 & ~n4435 ) ;
  assign n4437 = ( x77 & n4210 ) | ( x77 & ~n4354 ) | ( n4210 & ~n4354 ) ;
  assign n4438 = x77 & n4210 ;
  assign n4439 = ( ~n4215 & n4437 ) | ( ~n4215 & n4438 ) | ( n4437 & n4438 ) ;
  assign n4440 = ( n4215 & n4437 ) | ( n4215 & n4438 ) | ( n4437 & n4438 ) ;
  assign n4441 = ( n4215 & n4439 ) | ( n4215 & ~n4440 ) | ( n4439 & ~n4440 ) ;
  assign n4442 = ( x78 & n4436 ) | ( x78 & ~n4441 ) | ( n4436 & ~n4441 ) ;
  assign n4443 = ( x78 & n4216 ) | ( x78 & ~n4354 ) | ( n4216 & ~n4354 ) ;
  assign n4444 = x78 & n4216 ;
  assign n4445 = ( ~n4221 & n4443 ) | ( ~n4221 & n4444 ) | ( n4443 & n4444 ) ;
  assign n4446 = ( n4221 & n4443 ) | ( n4221 & n4444 ) | ( n4443 & n4444 ) ;
  assign n4447 = ( n4221 & n4445 ) | ( n4221 & ~n4446 ) | ( n4445 & ~n4446 ) ;
  assign n4448 = ( x79 & n4442 ) | ( x79 & ~n4447 ) | ( n4442 & ~n4447 ) ;
  assign n4449 = ( x79 & n4222 ) | ( x79 & ~n4354 ) | ( n4222 & ~n4354 ) ;
  assign n4450 = x79 & n4222 ;
  assign n4451 = ( ~n4227 & n4449 ) | ( ~n4227 & n4450 ) | ( n4449 & n4450 ) ;
  assign n4452 = ( n4227 & n4449 ) | ( n4227 & n4450 ) | ( n4449 & n4450 ) ;
  assign n4453 = ( n4227 & n4451 ) | ( n4227 & ~n4452 ) | ( n4451 & ~n4452 ) ;
  assign n4454 = ( x80 & n4448 ) | ( x80 & ~n4453 ) | ( n4448 & ~n4453 ) ;
  assign n4455 = ( x80 & n4228 ) | ( x80 & ~n4354 ) | ( n4228 & ~n4354 ) ;
  assign n4456 = x80 & n4228 ;
  assign n4457 = ( ~n4233 & n4455 ) | ( ~n4233 & n4456 ) | ( n4455 & n4456 ) ;
  assign n4458 = ( n4233 & n4455 ) | ( n4233 & n4456 ) | ( n4455 & n4456 ) ;
  assign n4459 = ( n4233 & n4457 ) | ( n4233 & ~n4458 ) | ( n4457 & ~n4458 ) ;
  assign n4460 = ( x81 & n4454 ) | ( x81 & ~n4459 ) | ( n4454 & ~n4459 ) ;
  assign n4461 = ( x81 & n4234 ) | ( x81 & ~n4354 ) | ( n4234 & ~n4354 ) ;
  assign n4462 = x81 & n4234 ;
  assign n4463 = ( ~n4239 & n4461 ) | ( ~n4239 & n4462 ) | ( n4461 & n4462 ) ;
  assign n4464 = ( n4239 & n4461 ) | ( n4239 & n4462 ) | ( n4461 & n4462 ) ;
  assign n4465 = ( n4239 & n4463 ) | ( n4239 & ~n4464 ) | ( n4463 & ~n4464 ) ;
  assign n4466 = ( x82 & n4460 ) | ( x82 & ~n4465 ) | ( n4460 & ~n4465 ) ;
  assign n4467 = ( x82 & n4240 ) | ( x82 & ~n4354 ) | ( n4240 & ~n4354 ) ;
  assign n4468 = x82 & n4240 ;
  assign n4469 = ( ~n4245 & n4467 ) | ( ~n4245 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4470 = ( n4245 & n4467 ) | ( n4245 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4471 = ( n4245 & n4469 ) | ( n4245 & ~n4470 ) | ( n4469 & ~n4470 ) ;
  assign n4472 = ( x83 & n4466 ) | ( x83 & ~n4471 ) | ( n4466 & ~n4471 ) ;
  assign n4473 = ( x83 & n4246 ) | ( x83 & ~n4354 ) | ( n4246 & ~n4354 ) ;
  assign n4474 = x83 & n4246 ;
  assign n4475 = ( ~n4251 & n4473 ) | ( ~n4251 & n4474 ) | ( n4473 & n4474 ) ;
  assign n4476 = ( n4251 & n4473 ) | ( n4251 & n4474 ) | ( n4473 & n4474 ) ;
  assign n4477 = ( n4251 & n4475 ) | ( n4251 & ~n4476 ) | ( n4475 & ~n4476 ) ;
  assign n4478 = ( x84 & n4472 ) | ( x84 & ~n4477 ) | ( n4472 & ~n4477 ) ;
  assign n4479 = ( x84 & n4252 ) | ( x84 & ~n4354 ) | ( n4252 & ~n4354 ) ;
  assign n4480 = x84 & n4252 ;
  assign n4481 = ( ~n4257 & n4479 ) | ( ~n4257 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = ( n4257 & n4479 ) | ( n4257 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4483 = ( n4257 & n4481 ) | ( n4257 & ~n4482 ) | ( n4481 & ~n4482 ) ;
  assign n4484 = ( x85 & n4478 ) | ( x85 & ~n4483 ) | ( n4478 & ~n4483 ) ;
  assign n4485 = ( x85 & n4258 ) | ( x85 & ~n4354 ) | ( n4258 & ~n4354 ) ;
  assign n4486 = x85 & n4258 ;
  assign n4487 = ( ~n4263 & n4485 ) | ( ~n4263 & n4486 ) | ( n4485 & n4486 ) ;
  assign n4488 = ( n4263 & n4485 ) | ( n4263 & n4486 ) | ( n4485 & n4486 ) ;
  assign n4489 = ( n4263 & n4487 ) | ( n4263 & ~n4488 ) | ( n4487 & ~n4488 ) ;
  assign n4490 = ( x86 & n4484 ) | ( x86 & ~n4489 ) | ( n4484 & ~n4489 ) ;
  assign n4491 = ( x86 & n4264 ) | ( x86 & ~n4354 ) | ( n4264 & ~n4354 ) ;
  assign n4492 = x86 & n4264 ;
  assign n4493 = ( ~n4269 & n4491 ) | ( ~n4269 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4494 = ( n4269 & n4491 ) | ( n4269 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4495 = ( n4269 & n4493 ) | ( n4269 & ~n4494 ) | ( n4493 & ~n4494 ) ;
  assign n4496 = ( x87 & n4490 ) | ( x87 & ~n4495 ) | ( n4490 & ~n4495 ) ;
  assign n4497 = ( x87 & n4270 ) | ( x87 & ~n4354 ) | ( n4270 & ~n4354 ) ;
  assign n4498 = x87 & n4270 ;
  assign n4499 = ( ~n4275 & n4497 ) | ( ~n4275 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4500 = ( n4275 & n4497 ) | ( n4275 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4501 = ( n4275 & n4499 ) | ( n4275 & ~n4500 ) | ( n4499 & ~n4500 ) ;
  assign n4502 = ( x88 & n4496 ) | ( x88 & ~n4501 ) | ( n4496 & ~n4501 ) ;
  assign n4503 = ( x88 & n4276 ) | ( x88 & ~n4354 ) | ( n4276 & ~n4354 ) ;
  assign n4504 = x88 & n4276 ;
  assign n4505 = ( ~n4281 & n4503 ) | ( ~n4281 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4506 = ( n4281 & n4503 ) | ( n4281 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4507 = ( n4281 & n4505 ) | ( n4281 & ~n4506 ) | ( n4505 & ~n4506 ) ;
  assign n4508 = ( x89 & n4502 ) | ( x89 & ~n4507 ) | ( n4502 & ~n4507 ) ;
  assign n4509 = ( x89 & n4282 ) | ( x89 & ~n4354 ) | ( n4282 & ~n4354 ) ;
  assign n4510 = x89 & n4282 ;
  assign n4511 = ( ~n4287 & n4509 ) | ( ~n4287 & n4510 ) | ( n4509 & n4510 ) ;
  assign n4512 = ( n4287 & n4509 ) | ( n4287 & n4510 ) | ( n4509 & n4510 ) ;
  assign n4513 = ( n4287 & n4511 ) | ( n4287 & ~n4512 ) | ( n4511 & ~n4512 ) ;
  assign n4514 = ( x90 & n4508 ) | ( x90 & ~n4513 ) | ( n4508 & ~n4513 ) ;
  assign n4515 = ( x90 & n4288 ) | ( x90 & ~n4354 ) | ( n4288 & ~n4354 ) ;
  assign n4516 = x90 & n4288 ;
  assign n4517 = ( ~n4293 & n4515 ) | ( ~n4293 & n4516 ) | ( n4515 & n4516 ) ;
  assign n4518 = ( n4293 & n4515 ) | ( n4293 & n4516 ) | ( n4515 & n4516 ) ;
  assign n4519 = ( n4293 & n4517 ) | ( n4293 & ~n4518 ) | ( n4517 & ~n4518 ) ;
  assign n4520 = ( x91 & n4514 ) | ( x91 & ~n4519 ) | ( n4514 & ~n4519 ) ;
  assign n4521 = ( x91 & n4294 ) | ( x91 & ~n4354 ) | ( n4294 & ~n4354 ) ;
  assign n4522 = x91 & n4294 ;
  assign n4523 = ( ~n4299 & n4521 ) | ( ~n4299 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4524 = ( n4299 & n4521 ) | ( n4299 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4525 = ( n4299 & n4523 ) | ( n4299 & ~n4524 ) | ( n4523 & ~n4524 ) ;
  assign n4526 = ( x92 & n4520 ) | ( x92 & ~n4525 ) | ( n4520 & ~n4525 ) ;
  assign n4527 = ( x92 & n4300 ) | ( x92 & ~n4354 ) | ( n4300 & ~n4354 ) ;
  assign n4528 = x92 & n4300 ;
  assign n4529 = ( ~n4305 & n4527 ) | ( ~n4305 & n4528 ) | ( n4527 & n4528 ) ;
  assign n4530 = ( n4305 & n4527 ) | ( n4305 & n4528 ) | ( n4527 & n4528 ) ;
  assign n4531 = ( n4305 & n4529 ) | ( n4305 & ~n4530 ) | ( n4529 & ~n4530 ) ;
  assign n4532 = ( x93 & n4526 ) | ( x93 & ~n4531 ) | ( n4526 & ~n4531 ) ;
  assign n4533 = ( x93 & n4306 ) | ( x93 & ~n4354 ) | ( n4306 & ~n4354 ) ;
  assign n4534 = x93 & n4306 ;
  assign n4535 = ( ~n4311 & n4533 ) | ( ~n4311 & n4534 ) | ( n4533 & n4534 ) ;
  assign n4536 = ( n4311 & n4533 ) | ( n4311 & n4534 ) | ( n4533 & n4534 ) ;
  assign n4537 = ( n4311 & n4535 ) | ( n4311 & ~n4536 ) | ( n4535 & ~n4536 ) ;
  assign n4538 = ( x94 & n4532 ) | ( x94 & ~n4537 ) | ( n4532 & ~n4537 ) ;
  assign n4539 = ( x94 & n4312 ) | ( x94 & ~n4354 ) | ( n4312 & ~n4354 ) ;
  assign n4540 = x94 & n4312 ;
  assign n4541 = ( ~n4317 & n4539 ) | ( ~n4317 & n4540 ) | ( n4539 & n4540 ) ;
  assign n4542 = ( n4317 & n4539 ) | ( n4317 & n4540 ) | ( n4539 & n4540 ) ;
  assign n4543 = ( n4317 & n4541 ) | ( n4317 & ~n4542 ) | ( n4541 & ~n4542 ) ;
  assign n4544 = ( x95 & n4538 ) | ( x95 & ~n4543 ) | ( n4538 & ~n4543 ) ;
  assign n4545 = ( x95 & n4318 ) | ( x95 & ~n4354 ) | ( n4318 & ~n4354 ) ;
  assign n4546 = x95 & n4318 ;
  assign n4547 = ( ~n4323 & n4545 ) | ( ~n4323 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4548 = ( n4323 & n4545 ) | ( n4323 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4549 = ( n4323 & n4547 ) | ( n4323 & ~n4548 ) | ( n4547 & ~n4548 ) ;
  assign n4550 = ( x96 & n4544 ) | ( x96 & ~n4549 ) | ( n4544 & ~n4549 ) ;
  assign n4551 = ( x96 & n4324 ) | ( x96 & ~n4354 ) | ( n4324 & ~n4354 ) ;
  assign n4552 = x96 & n4324 ;
  assign n4553 = ( ~n4329 & n4551 ) | ( ~n4329 & n4552 ) | ( n4551 & n4552 ) ;
  assign n4554 = ( n4329 & n4551 ) | ( n4329 & n4552 ) | ( n4551 & n4552 ) ;
  assign n4555 = ( n4329 & n4553 ) | ( n4329 & ~n4554 ) | ( n4553 & ~n4554 ) ;
  assign n4556 = ( x97 & n4550 ) | ( x97 & ~n4555 ) | ( n4550 & ~n4555 ) ;
  assign n4557 = ( x97 & n4330 ) | ( x97 & ~n4354 ) | ( n4330 & ~n4354 ) ;
  assign n4558 = x97 & n4330 ;
  assign n4559 = ( ~n4335 & n4557 ) | ( ~n4335 & n4558 ) | ( n4557 & n4558 ) ;
  assign n4560 = ( n4335 & n4557 ) | ( n4335 & n4558 ) | ( n4557 & n4558 ) ;
  assign n4561 = ( n4335 & n4559 ) | ( n4335 & ~n4560 ) | ( n4559 & ~n4560 ) ;
  assign n4562 = ( x98 & n4556 ) | ( x98 & ~n4561 ) | ( n4556 & ~n4561 ) ;
  assign n4563 = ( x98 & n4336 ) | ( x98 & ~n4354 ) | ( n4336 & ~n4354 ) ;
  assign n4564 = x98 & n4336 ;
  assign n4565 = ( ~n4341 & n4563 ) | ( ~n4341 & n4564 ) | ( n4563 & n4564 ) ;
  assign n4566 = ( n4341 & n4563 ) | ( n4341 & n4564 ) | ( n4563 & n4564 ) ;
  assign n4567 = ( n4341 & n4565 ) | ( n4341 & ~n4566 ) | ( n4565 & ~n4566 ) ;
  assign n4568 = ( x99 & n4562 ) | ( x99 & ~n4567 ) | ( n4562 & ~n4567 ) ;
  assign n4569 = ( x99 & n4342 ) | ( x99 & ~n4354 ) | ( n4342 & ~n4354 ) ;
  assign n4570 = x99 & n4342 ;
  assign n4571 = ( ~n4347 & n4569 ) | ( ~n4347 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = ( n4347 & n4569 ) | ( n4347 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4573 = ( n4347 & n4571 ) | ( n4347 & ~n4572 ) | ( n4571 & ~n4572 ) ;
  assign n4574 = ( x100 & n4568 ) | ( x100 & ~n4573 ) | ( n4568 & ~n4573 ) ;
  assign n4575 = ( x101 & ~n4359 ) | ( x101 & n4574 ) | ( ~n4359 & n4574 ) ;
  assign n4576 = ( x101 & x102 ) | ( x101 & ~n4352 ) | ( x102 & ~n4352 ) ;
  assign n4577 = ( ~x101 & x102 ) | ( ~x101 & n4352 ) | ( x102 & n4352 ) ;
  assign n4578 = n4576 | n4577 ;
  assign n4579 = ~n154 & n4351 ;
  assign n4580 = ~n4578 & n4579 ;
  assign n4581 = n155 & ~n4579 ;
  assign n4582 = ( n4575 & ~n4580 ) | ( n4575 & n4581 ) | ( ~n4580 & n4581 ) ;
  assign n4583 = ( x101 & n4574 ) | ( x101 & ~n4582 ) | ( n4574 & ~n4582 ) ;
  assign n4584 = x101 & n4574 ;
  assign n4585 = ( ~n4359 & n4583 ) | ( ~n4359 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4586 = ( n4359 & n4583 ) | ( n4359 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4587 = ( n4359 & n4585 ) | ( n4359 & ~n4586 ) | ( n4585 & ~n4586 ) ;
  assign n4588 = ~x24 & x64 ;
  assign n4589 = x25 & n4582 ;
  assign n4590 = ( x25 & x64 ) | ( x25 & ~n4582 ) | ( x64 & ~n4582 ) ;
  assign n4591 = x25 & x64 ;
  assign n4592 = ( n4589 & n4590 ) | ( n4589 & ~n4591 ) | ( n4590 & ~n4591 ) ;
  assign n4593 = ( x65 & n4588 ) | ( x65 & ~n4592 ) | ( n4588 & ~n4592 ) ;
  assign n4594 = ( x65 & n4360 ) | ( x65 & n4582 ) | ( n4360 & n4582 ) ;
  assign n4595 = x65 | n4360 ;
  assign n4596 = ( ~n4363 & n4594 ) | ( ~n4363 & n4595 ) | ( n4594 & n4595 ) ;
  assign n4597 = ( n4363 & n4594 ) | ( n4363 & n4595 ) | ( n4594 & n4595 ) ;
  assign n4598 = ( n4363 & n4596 ) | ( n4363 & ~n4597 ) | ( n4596 & ~n4597 ) ;
  assign n4599 = ( x66 & n4593 ) | ( x66 & ~n4598 ) | ( n4593 & ~n4598 ) ;
  assign n4600 = ( x66 & n4364 ) | ( x66 & n4582 ) | ( n4364 & n4582 ) ;
  assign n4601 = x66 | n4364 ;
  assign n4602 = ( ~n4369 & n4600 ) | ( ~n4369 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4603 = ( n4369 & n4600 ) | ( n4369 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4604 = ( n4369 & n4602 ) | ( n4369 & ~n4603 ) | ( n4602 & ~n4603 ) ;
  assign n4605 = ( x67 & n4599 ) | ( x67 & ~n4604 ) | ( n4599 & ~n4604 ) ;
  assign n4606 = ( x67 & n4370 ) | ( x67 & ~n4582 ) | ( n4370 & ~n4582 ) ;
  assign n4607 = x67 & n4370 ;
  assign n4608 = ( ~n4375 & n4606 ) | ( ~n4375 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4609 = ( n4375 & n4606 ) | ( n4375 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4610 = ( n4375 & n4608 ) | ( n4375 & ~n4609 ) | ( n4608 & ~n4609 ) ;
  assign n4611 = ( x68 & n4605 ) | ( x68 & ~n4610 ) | ( n4605 & ~n4610 ) ;
  assign n4612 = ( x68 & n4376 ) | ( x68 & ~n4582 ) | ( n4376 & ~n4582 ) ;
  assign n4613 = x68 & n4376 ;
  assign n4614 = ( ~n4381 & n4612 ) | ( ~n4381 & n4613 ) | ( n4612 & n4613 ) ;
  assign n4615 = ( n4381 & n4612 ) | ( n4381 & n4613 ) | ( n4612 & n4613 ) ;
  assign n4616 = ( n4381 & n4614 ) | ( n4381 & ~n4615 ) | ( n4614 & ~n4615 ) ;
  assign n4617 = ( x69 & n4611 ) | ( x69 & ~n4616 ) | ( n4611 & ~n4616 ) ;
  assign n4618 = ( x69 & n4382 ) | ( x69 & ~n4582 ) | ( n4382 & ~n4582 ) ;
  assign n4619 = x69 & n4382 ;
  assign n4620 = ( ~n4387 & n4618 ) | ( ~n4387 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4621 = ( n4387 & n4618 ) | ( n4387 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4622 = ( n4387 & n4620 ) | ( n4387 & ~n4621 ) | ( n4620 & ~n4621 ) ;
  assign n4623 = ( x70 & n4617 ) | ( x70 & ~n4622 ) | ( n4617 & ~n4622 ) ;
  assign n4624 = ( x70 & n4388 ) | ( x70 & ~n4582 ) | ( n4388 & ~n4582 ) ;
  assign n4625 = x70 & n4388 ;
  assign n4626 = ( ~n4393 & n4624 ) | ( ~n4393 & n4625 ) | ( n4624 & n4625 ) ;
  assign n4627 = ( n4393 & n4624 ) | ( n4393 & n4625 ) | ( n4624 & n4625 ) ;
  assign n4628 = ( n4393 & n4626 ) | ( n4393 & ~n4627 ) | ( n4626 & ~n4627 ) ;
  assign n4629 = ( x71 & n4623 ) | ( x71 & ~n4628 ) | ( n4623 & ~n4628 ) ;
  assign n4630 = ( x71 & n4394 ) | ( x71 & ~n4582 ) | ( n4394 & ~n4582 ) ;
  assign n4631 = x71 & n4394 ;
  assign n4632 = ( ~n4399 & n4630 ) | ( ~n4399 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4633 = ( n4399 & n4630 ) | ( n4399 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4634 = ( n4399 & n4632 ) | ( n4399 & ~n4633 ) | ( n4632 & ~n4633 ) ;
  assign n4635 = ( x72 & n4629 ) | ( x72 & ~n4634 ) | ( n4629 & ~n4634 ) ;
  assign n4636 = ( x72 & n4400 ) | ( x72 & ~n4582 ) | ( n4400 & ~n4582 ) ;
  assign n4637 = x72 & n4400 ;
  assign n4638 = ( ~n4405 & n4636 ) | ( ~n4405 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4639 = ( n4405 & n4636 ) | ( n4405 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4640 = ( n4405 & n4638 ) | ( n4405 & ~n4639 ) | ( n4638 & ~n4639 ) ;
  assign n4641 = ( x73 & n4635 ) | ( x73 & ~n4640 ) | ( n4635 & ~n4640 ) ;
  assign n4642 = ( x73 & n4406 ) | ( x73 & ~n4582 ) | ( n4406 & ~n4582 ) ;
  assign n4643 = x73 & n4406 ;
  assign n4644 = ( ~n4411 & n4642 ) | ( ~n4411 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4645 = ( n4411 & n4642 ) | ( n4411 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4646 = ( n4411 & n4644 ) | ( n4411 & ~n4645 ) | ( n4644 & ~n4645 ) ;
  assign n4647 = ( x74 & n4641 ) | ( x74 & ~n4646 ) | ( n4641 & ~n4646 ) ;
  assign n4648 = ( x74 & n4412 ) | ( x74 & ~n4582 ) | ( n4412 & ~n4582 ) ;
  assign n4649 = x74 & n4412 ;
  assign n4650 = ( ~n4417 & n4648 ) | ( ~n4417 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4651 = ( n4417 & n4648 ) | ( n4417 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4652 = ( n4417 & n4650 ) | ( n4417 & ~n4651 ) | ( n4650 & ~n4651 ) ;
  assign n4653 = ( x75 & n4647 ) | ( x75 & ~n4652 ) | ( n4647 & ~n4652 ) ;
  assign n4654 = ( x75 & n4418 ) | ( x75 & ~n4582 ) | ( n4418 & ~n4582 ) ;
  assign n4655 = x75 & n4418 ;
  assign n4656 = ( ~n4423 & n4654 ) | ( ~n4423 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = ( n4423 & n4654 ) | ( n4423 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4658 = ( n4423 & n4656 ) | ( n4423 & ~n4657 ) | ( n4656 & ~n4657 ) ;
  assign n4659 = ( x76 & n4653 ) | ( x76 & ~n4658 ) | ( n4653 & ~n4658 ) ;
  assign n4660 = ( x76 & n4424 ) | ( x76 & ~n4582 ) | ( n4424 & ~n4582 ) ;
  assign n4661 = x76 & n4424 ;
  assign n4662 = ( ~n4429 & n4660 ) | ( ~n4429 & n4661 ) | ( n4660 & n4661 ) ;
  assign n4663 = ( n4429 & n4660 ) | ( n4429 & n4661 ) | ( n4660 & n4661 ) ;
  assign n4664 = ( n4429 & n4662 ) | ( n4429 & ~n4663 ) | ( n4662 & ~n4663 ) ;
  assign n4665 = ( x77 & n4659 ) | ( x77 & ~n4664 ) | ( n4659 & ~n4664 ) ;
  assign n4666 = ( x77 & n4430 ) | ( x77 & ~n4582 ) | ( n4430 & ~n4582 ) ;
  assign n4667 = x77 & n4430 ;
  assign n4668 = ( ~n4435 & n4666 ) | ( ~n4435 & n4667 ) | ( n4666 & n4667 ) ;
  assign n4669 = ( n4435 & n4666 ) | ( n4435 & n4667 ) | ( n4666 & n4667 ) ;
  assign n4670 = ( n4435 & n4668 ) | ( n4435 & ~n4669 ) | ( n4668 & ~n4669 ) ;
  assign n4671 = ( x78 & n4665 ) | ( x78 & ~n4670 ) | ( n4665 & ~n4670 ) ;
  assign n4672 = ( x78 & n4436 ) | ( x78 & ~n4582 ) | ( n4436 & ~n4582 ) ;
  assign n4673 = x78 & n4436 ;
  assign n4674 = ( ~n4441 & n4672 ) | ( ~n4441 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4675 = ( n4441 & n4672 ) | ( n4441 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4676 = ( n4441 & n4674 ) | ( n4441 & ~n4675 ) | ( n4674 & ~n4675 ) ;
  assign n4677 = ( x79 & n4671 ) | ( x79 & ~n4676 ) | ( n4671 & ~n4676 ) ;
  assign n4678 = ( x79 & n4442 ) | ( x79 & ~n4582 ) | ( n4442 & ~n4582 ) ;
  assign n4679 = x79 & n4442 ;
  assign n4680 = ( ~n4447 & n4678 ) | ( ~n4447 & n4679 ) | ( n4678 & n4679 ) ;
  assign n4681 = ( n4447 & n4678 ) | ( n4447 & n4679 ) | ( n4678 & n4679 ) ;
  assign n4682 = ( n4447 & n4680 ) | ( n4447 & ~n4681 ) | ( n4680 & ~n4681 ) ;
  assign n4683 = ( x80 & n4677 ) | ( x80 & ~n4682 ) | ( n4677 & ~n4682 ) ;
  assign n4684 = ( x80 & n4448 ) | ( x80 & ~n4582 ) | ( n4448 & ~n4582 ) ;
  assign n4685 = x80 & n4448 ;
  assign n4686 = ( ~n4453 & n4684 ) | ( ~n4453 & n4685 ) | ( n4684 & n4685 ) ;
  assign n4687 = ( n4453 & n4684 ) | ( n4453 & n4685 ) | ( n4684 & n4685 ) ;
  assign n4688 = ( n4453 & n4686 ) | ( n4453 & ~n4687 ) | ( n4686 & ~n4687 ) ;
  assign n4689 = ( x81 & n4683 ) | ( x81 & ~n4688 ) | ( n4683 & ~n4688 ) ;
  assign n4690 = ( x81 & n4454 ) | ( x81 & ~n4582 ) | ( n4454 & ~n4582 ) ;
  assign n4691 = x81 & n4454 ;
  assign n4692 = ( ~n4459 & n4690 ) | ( ~n4459 & n4691 ) | ( n4690 & n4691 ) ;
  assign n4693 = ( n4459 & n4690 ) | ( n4459 & n4691 ) | ( n4690 & n4691 ) ;
  assign n4694 = ( n4459 & n4692 ) | ( n4459 & ~n4693 ) | ( n4692 & ~n4693 ) ;
  assign n4695 = ( x82 & n4689 ) | ( x82 & ~n4694 ) | ( n4689 & ~n4694 ) ;
  assign n4696 = ( x82 & n4460 ) | ( x82 & ~n4582 ) | ( n4460 & ~n4582 ) ;
  assign n4697 = x82 & n4460 ;
  assign n4698 = ( ~n4465 & n4696 ) | ( ~n4465 & n4697 ) | ( n4696 & n4697 ) ;
  assign n4699 = ( n4465 & n4696 ) | ( n4465 & n4697 ) | ( n4696 & n4697 ) ;
  assign n4700 = ( n4465 & n4698 ) | ( n4465 & ~n4699 ) | ( n4698 & ~n4699 ) ;
  assign n4701 = ( x83 & n4695 ) | ( x83 & ~n4700 ) | ( n4695 & ~n4700 ) ;
  assign n4702 = ( x83 & n4466 ) | ( x83 & ~n4582 ) | ( n4466 & ~n4582 ) ;
  assign n4703 = x83 & n4466 ;
  assign n4704 = ( ~n4471 & n4702 ) | ( ~n4471 & n4703 ) | ( n4702 & n4703 ) ;
  assign n4705 = ( n4471 & n4702 ) | ( n4471 & n4703 ) | ( n4702 & n4703 ) ;
  assign n4706 = ( n4471 & n4704 ) | ( n4471 & ~n4705 ) | ( n4704 & ~n4705 ) ;
  assign n4707 = ( x84 & n4701 ) | ( x84 & ~n4706 ) | ( n4701 & ~n4706 ) ;
  assign n4708 = ( x84 & n4472 ) | ( x84 & ~n4582 ) | ( n4472 & ~n4582 ) ;
  assign n4709 = x84 & n4472 ;
  assign n4710 = ( ~n4477 & n4708 ) | ( ~n4477 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4711 = ( n4477 & n4708 ) | ( n4477 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4712 = ( n4477 & n4710 ) | ( n4477 & ~n4711 ) | ( n4710 & ~n4711 ) ;
  assign n4713 = ( x85 & n4707 ) | ( x85 & ~n4712 ) | ( n4707 & ~n4712 ) ;
  assign n4714 = ( x85 & n4478 ) | ( x85 & ~n4582 ) | ( n4478 & ~n4582 ) ;
  assign n4715 = x85 & n4478 ;
  assign n4716 = ( ~n4483 & n4714 ) | ( ~n4483 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4717 = ( n4483 & n4714 ) | ( n4483 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4718 = ( n4483 & n4716 ) | ( n4483 & ~n4717 ) | ( n4716 & ~n4717 ) ;
  assign n4719 = ( x86 & n4713 ) | ( x86 & ~n4718 ) | ( n4713 & ~n4718 ) ;
  assign n4720 = ( x86 & n4484 ) | ( x86 & ~n4582 ) | ( n4484 & ~n4582 ) ;
  assign n4721 = x86 & n4484 ;
  assign n4722 = ( ~n4489 & n4720 ) | ( ~n4489 & n4721 ) | ( n4720 & n4721 ) ;
  assign n4723 = ( n4489 & n4720 ) | ( n4489 & n4721 ) | ( n4720 & n4721 ) ;
  assign n4724 = ( n4489 & n4722 ) | ( n4489 & ~n4723 ) | ( n4722 & ~n4723 ) ;
  assign n4725 = ( x87 & n4719 ) | ( x87 & ~n4724 ) | ( n4719 & ~n4724 ) ;
  assign n4726 = ( x87 & n4490 ) | ( x87 & ~n4582 ) | ( n4490 & ~n4582 ) ;
  assign n4727 = x87 & n4490 ;
  assign n4728 = ( ~n4495 & n4726 ) | ( ~n4495 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4729 = ( n4495 & n4726 ) | ( n4495 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4730 = ( n4495 & n4728 ) | ( n4495 & ~n4729 ) | ( n4728 & ~n4729 ) ;
  assign n4731 = ( x88 & n4725 ) | ( x88 & ~n4730 ) | ( n4725 & ~n4730 ) ;
  assign n4732 = ( x88 & n4496 ) | ( x88 & ~n4582 ) | ( n4496 & ~n4582 ) ;
  assign n4733 = x88 & n4496 ;
  assign n4734 = ( ~n4501 & n4732 ) | ( ~n4501 & n4733 ) | ( n4732 & n4733 ) ;
  assign n4735 = ( n4501 & n4732 ) | ( n4501 & n4733 ) | ( n4732 & n4733 ) ;
  assign n4736 = ( n4501 & n4734 ) | ( n4501 & ~n4735 ) | ( n4734 & ~n4735 ) ;
  assign n4737 = ( x89 & n4731 ) | ( x89 & ~n4736 ) | ( n4731 & ~n4736 ) ;
  assign n4738 = ( x89 & n4502 ) | ( x89 & ~n4582 ) | ( n4502 & ~n4582 ) ;
  assign n4739 = x89 & n4502 ;
  assign n4740 = ( ~n4507 & n4738 ) | ( ~n4507 & n4739 ) | ( n4738 & n4739 ) ;
  assign n4741 = ( n4507 & n4738 ) | ( n4507 & n4739 ) | ( n4738 & n4739 ) ;
  assign n4742 = ( n4507 & n4740 ) | ( n4507 & ~n4741 ) | ( n4740 & ~n4741 ) ;
  assign n4743 = ( x90 & n4737 ) | ( x90 & ~n4742 ) | ( n4737 & ~n4742 ) ;
  assign n4744 = ( x90 & n4508 ) | ( x90 & ~n4582 ) | ( n4508 & ~n4582 ) ;
  assign n4745 = x90 & n4508 ;
  assign n4746 = ( ~n4513 & n4744 ) | ( ~n4513 & n4745 ) | ( n4744 & n4745 ) ;
  assign n4747 = ( n4513 & n4744 ) | ( n4513 & n4745 ) | ( n4744 & n4745 ) ;
  assign n4748 = ( n4513 & n4746 ) | ( n4513 & ~n4747 ) | ( n4746 & ~n4747 ) ;
  assign n4749 = ( x91 & n4743 ) | ( x91 & ~n4748 ) | ( n4743 & ~n4748 ) ;
  assign n4750 = ( x91 & n4514 ) | ( x91 & ~n4582 ) | ( n4514 & ~n4582 ) ;
  assign n4751 = x91 & n4514 ;
  assign n4752 = ( ~n4519 & n4750 ) | ( ~n4519 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4753 = ( n4519 & n4750 ) | ( n4519 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4754 = ( n4519 & n4752 ) | ( n4519 & ~n4753 ) | ( n4752 & ~n4753 ) ;
  assign n4755 = ( x92 & n4749 ) | ( x92 & ~n4754 ) | ( n4749 & ~n4754 ) ;
  assign n4756 = ( x92 & n4520 ) | ( x92 & ~n4582 ) | ( n4520 & ~n4582 ) ;
  assign n4757 = x92 & n4520 ;
  assign n4758 = ( ~n4525 & n4756 ) | ( ~n4525 & n4757 ) | ( n4756 & n4757 ) ;
  assign n4759 = ( n4525 & n4756 ) | ( n4525 & n4757 ) | ( n4756 & n4757 ) ;
  assign n4760 = ( n4525 & n4758 ) | ( n4525 & ~n4759 ) | ( n4758 & ~n4759 ) ;
  assign n4761 = ( x93 & n4755 ) | ( x93 & ~n4760 ) | ( n4755 & ~n4760 ) ;
  assign n4762 = ( x93 & n4526 ) | ( x93 & ~n4582 ) | ( n4526 & ~n4582 ) ;
  assign n4763 = x93 & n4526 ;
  assign n4764 = ( ~n4531 & n4762 ) | ( ~n4531 & n4763 ) | ( n4762 & n4763 ) ;
  assign n4765 = ( n4531 & n4762 ) | ( n4531 & n4763 ) | ( n4762 & n4763 ) ;
  assign n4766 = ( n4531 & n4764 ) | ( n4531 & ~n4765 ) | ( n4764 & ~n4765 ) ;
  assign n4767 = ( x94 & n4761 ) | ( x94 & ~n4766 ) | ( n4761 & ~n4766 ) ;
  assign n4768 = ( x94 & n4532 ) | ( x94 & ~n4582 ) | ( n4532 & ~n4582 ) ;
  assign n4769 = x94 & n4532 ;
  assign n4770 = ( ~n4537 & n4768 ) | ( ~n4537 & n4769 ) | ( n4768 & n4769 ) ;
  assign n4771 = ( n4537 & n4768 ) | ( n4537 & n4769 ) | ( n4768 & n4769 ) ;
  assign n4772 = ( n4537 & n4770 ) | ( n4537 & ~n4771 ) | ( n4770 & ~n4771 ) ;
  assign n4773 = ( x95 & n4767 ) | ( x95 & ~n4772 ) | ( n4767 & ~n4772 ) ;
  assign n4774 = ( x95 & n4538 ) | ( x95 & ~n4582 ) | ( n4538 & ~n4582 ) ;
  assign n4775 = x95 & n4538 ;
  assign n4776 = ( ~n4543 & n4774 ) | ( ~n4543 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4777 = ( n4543 & n4774 ) | ( n4543 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4778 = ( n4543 & n4776 ) | ( n4543 & ~n4777 ) | ( n4776 & ~n4777 ) ;
  assign n4779 = ( x96 & n4773 ) | ( x96 & ~n4778 ) | ( n4773 & ~n4778 ) ;
  assign n4780 = ( x96 & n4544 ) | ( x96 & ~n4582 ) | ( n4544 & ~n4582 ) ;
  assign n4781 = x96 & n4544 ;
  assign n4782 = ( ~n4549 & n4780 ) | ( ~n4549 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4783 = ( n4549 & n4780 ) | ( n4549 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4784 = ( n4549 & n4782 ) | ( n4549 & ~n4783 ) | ( n4782 & ~n4783 ) ;
  assign n4785 = ( x97 & n4779 ) | ( x97 & ~n4784 ) | ( n4779 & ~n4784 ) ;
  assign n4786 = ( x97 & n4550 ) | ( x97 & ~n4582 ) | ( n4550 & ~n4582 ) ;
  assign n4787 = x97 & n4550 ;
  assign n4788 = ( ~n4555 & n4786 ) | ( ~n4555 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4789 = ( n4555 & n4786 ) | ( n4555 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4790 = ( n4555 & n4788 ) | ( n4555 & ~n4789 ) | ( n4788 & ~n4789 ) ;
  assign n4791 = ( x98 & n4785 ) | ( x98 & ~n4790 ) | ( n4785 & ~n4790 ) ;
  assign n4792 = ( x98 & n4556 ) | ( x98 & ~n4582 ) | ( n4556 & ~n4582 ) ;
  assign n4793 = x98 & n4556 ;
  assign n4794 = ( ~n4561 & n4792 ) | ( ~n4561 & n4793 ) | ( n4792 & n4793 ) ;
  assign n4795 = ( n4561 & n4792 ) | ( n4561 & n4793 ) | ( n4792 & n4793 ) ;
  assign n4796 = ( n4561 & n4794 ) | ( n4561 & ~n4795 ) | ( n4794 & ~n4795 ) ;
  assign n4797 = ( x99 & n4791 ) | ( x99 & ~n4796 ) | ( n4791 & ~n4796 ) ;
  assign n4798 = ( x99 & n4562 ) | ( x99 & ~n4582 ) | ( n4562 & ~n4582 ) ;
  assign n4799 = x99 & n4562 ;
  assign n4800 = ( ~n4567 & n4798 ) | ( ~n4567 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4801 = ( n4567 & n4798 ) | ( n4567 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4802 = ( n4567 & n4800 ) | ( n4567 & ~n4801 ) | ( n4800 & ~n4801 ) ;
  assign n4803 = ( x100 & n4797 ) | ( x100 & ~n4802 ) | ( n4797 & ~n4802 ) ;
  assign n4804 = ( x100 & n4568 ) | ( x100 & ~n4582 ) | ( n4568 & ~n4582 ) ;
  assign n4805 = x100 & n4568 ;
  assign n4806 = ( ~n4573 & n4804 ) | ( ~n4573 & n4805 ) | ( n4804 & n4805 ) ;
  assign n4807 = ( n4573 & n4804 ) | ( n4573 & n4805 ) | ( n4804 & n4805 ) ;
  assign n4808 = ( n4573 & n4806 ) | ( n4573 & ~n4807 ) | ( n4806 & ~n4807 ) ;
  assign n4809 = ( x101 & n4803 ) | ( x101 & ~n4808 ) | ( n4803 & ~n4808 ) ;
  assign n4810 = ( x102 & ~n4587 ) | ( x102 & n4809 ) | ( ~n4587 & n4809 ) ;
  assign n4811 = n155 & n4575 ;
  assign n4812 = ~n154 & n4578 ;
  assign n4813 = n4575 | n4812 ;
  assign n4814 = ( n4351 & n4811 ) | ( n4351 & ~n4813 ) | ( n4811 & ~n4813 ) ;
  assign n4815 = ( x103 & n4810 ) | ( x103 & ~n4814 ) | ( n4810 & ~n4814 ) ;
  assign n4816 = n153 | n4815 ;
  assign n4817 = ( x102 & n4809 ) | ( x102 & n4816 ) | ( n4809 & n4816 ) ;
  assign n4818 = x102 | n4809 ;
  assign n4819 = ( ~n4587 & n4817 ) | ( ~n4587 & n4818 ) | ( n4817 & n4818 ) ;
  assign n4820 = ( n4587 & n4817 ) | ( n4587 & n4818 ) | ( n4817 & n4818 ) ;
  assign n4821 = ( n4587 & n4819 ) | ( n4587 & ~n4820 ) | ( n4819 & ~n4820 ) ;
  assign n4822 = ~x23 & x64 ;
  assign n4823 = ~x24 & n4816 ;
  assign n4824 = ( x24 & ~x64 ) | ( x24 & n4816 ) | ( ~x64 & n4816 ) ;
  assign n4825 = ( n4588 & ~n4823 ) | ( n4588 & n4824 ) | ( ~n4823 & n4824 ) ;
  assign n4826 = ( x65 & n4822 ) | ( x65 & ~n4825 ) | ( n4822 & ~n4825 ) ;
  assign n4827 = ( x65 & n4588 ) | ( x65 & n4816 ) | ( n4588 & n4816 ) ;
  assign n4828 = x65 | n4588 ;
  assign n4829 = ( ~n4592 & n4827 ) | ( ~n4592 & n4828 ) | ( n4827 & n4828 ) ;
  assign n4830 = ( n4592 & n4827 ) | ( n4592 & n4828 ) | ( n4827 & n4828 ) ;
  assign n4831 = ( n4592 & n4829 ) | ( n4592 & ~n4830 ) | ( n4829 & ~n4830 ) ;
  assign n4832 = ( x66 & n4826 ) | ( x66 & ~n4831 ) | ( n4826 & ~n4831 ) ;
  assign n4833 = ( x66 & n4593 ) | ( x66 & n4816 ) | ( n4593 & n4816 ) ;
  assign n4834 = x66 | n4593 ;
  assign n4835 = ( ~n4598 & n4833 ) | ( ~n4598 & n4834 ) | ( n4833 & n4834 ) ;
  assign n4836 = ( n4598 & n4833 ) | ( n4598 & n4834 ) | ( n4833 & n4834 ) ;
  assign n4837 = ( n4598 & n4835 ) | ( n4598 & ~n4836 ) | ( n4835 & ~n4836 ) ;
  assign n4838 = ( x67 & n4832 ) | ( x67 & ~n4837 ) | ( n4832 & ~n4837 ) ;
  assign n4839 = ( x67 & n4599 ) | ( x67 & ~n4816 ) | ( n4599 & ~n4816 ) ;
  assign n4840 = x67 & n4599 ;
  assign n4841 = ( ~n4604 & n4839 ) | ( ~n4604 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4842 = ( n4604 & n4839 ) | ( n4604 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4843 = ( n4604 & n4841 ) | ( n4604 & ~n4842 ) | ( n4841 & ~n4842 ) ;
  assign n4844 = ( x68 & n4838 ) | ( x68 & ~n4843 ) | ( n4838 & ~n4843 ) ;
  assign n4845 = ( x68 & n4605 ) | ( x68 & ~n4816 ) | ( n4605 & ~n4816 ) ;
  assign n4846 = x68 & n4605 ;
  assign n4847 = ( ~n4610 & n4845 ) | ( ~n4610 & n4846 ) | ( n4845 & n4846 ) ;
  assign n4848 = ( n4610 & n4845 ) | ( n4610 & n4846 ) | ( n4845 & n4846 ) ;
  assign n4849 = ( n4610 & n4847 ) | ( n4610 & ~n4848 ) | ( n4847 & ~n4848 ) ;
  assign n4850 = ( x69 & n4844 ) | ( x69 & ~n4849 ) | ( n4844 & ~n4849 ) ;
  assign n4851 = ( x69 & n4611 ) | ( x69 & ~n4816 ) | ( n4611 & ~n4816 ) ;
  assign n4852 = x69 & n4611 ;
  assign n4853 = ( ~n4616 & n4851 ) | ( ~n4616 & n4852 ) | ( n4851 & n4852 ) ;
  assign n4854 = ( n4616 & n4851 ) | ( n4616 & n4852 ) | ( n4851 & n4852 ) ;
  assign n4855 = ( n4616 & n4853 ) | ( n4616 & ~n4854 ) | ( n4853 & ~n4854 ) ;
  assign n4856 = ( x70 & n4850 ) | ( x70 & ~n4855 ) | ( n4850 & ~n4855 ) ;
  assign n4857 = ( x70 & n4617 ) | ( x70 & ~n4816 ) | ( n4617 & ~n4816 ) ;
  assign n4858 = x70 & n4617 ;
  assign n4859 = ( ~n4622 & n4857 ) | ( ~n4622 & n4858 ) | ( n4857 & n4858 ) ;
  assign n4860 = ( n4622 & n4857 ) | ( n4622 & n4858 ) | ( n4857 & n4858 ) ;
  assign n4861 = ( n4622 & n4859 ) | ( n4622 & ~n4860 ) | ( n4859 & ~n4860 ) ;
  assign n4862 = ( x71 & n4856 ) | ( x71 & ~n4861 ) | ( n4856 & ~n4861 ) ;
  assign n4863 = ( x71 & n4623 ) | ( x71 & ~n4816 ) | ( n4623 & ~n4816 ) ;
  assign n4864 = x71 & n4623 ;
  assign n4865 = ( ~n4628 & n4863 ) | ( ~n4628 & n4864 ) | ( n4863 & n4864 ) ;
  assign n4866 = ( n4628 & n4863 ) | ( n4628 & n4864 ) | ( n4863 & n4864 ) ;
  assign n4867 = ( n4628 & n4865 ) | ( n4628 & ~n4866 ) | ( n4865 & ~n4866 ) ;
  assign n4868 = ( x72 & n4862 ) | ( x72 & ~n4867 ) | ( n4862 & ~n4867 ) ;
  assign n4869 = ( x72 & n4629 ) | ( x72 & ~n4816 ) | ( n4629 & ~n4816 ) ;
  assign n4870 = x72 & n4629 ;
  assign n4871 = ( ~n4634 & n4869 ) | ( ~n4634 & n4870 ) | ( n4869 & n4870 ) ;
  assign n4872 = ( n4634 & n4869 ) | ( n4634 & n4870 ) | ( n4869 & n4870 ) ;
  assign n4873 = ( n4634 & n4871 ) | ( n4634 & ~n4872 ) | ( n4871 & ~n4872 ) ;
  assign n4874 = ( x73 & n4868 ) | ( x73 & ~n4873 ) | ( n4868 & ~n4873 ) ;
  assign n4875 = ( x73 & n4635 ) | ( x73 & ~n4816 ) | ( n4635 & ~n4816 ) ;
  assign n4876 = x73 & n4635 ;
  assign n4877 = ( ~n4640 & n4875 ) | ( ~n4640 & n4876 ) | ( n4875 & n4876 ) ;
  assign n4878 = ( n4640 & n4875 ) | ( n4640 & n4876 ) | ( n4875 & n4876 ) ;
  assign n4879 = ( n4640 & n4877 ) | ( n4640 & ~n4878 ) | ( n4877 & ~n4878 ) ;
  assign n4880 = ( x74 & n4874 ) | ( x74 & ~n4879 ) | ( n4874 & ~n4879 ) ;
  assign n4881 = ( x74 & n4641 ) | ( x74 & ~n4816 ) | ( n4641 & ~n4816 ) ;
  assign n4882 = x74 & n4641 ;
  assign n4883 = ( ~n4646 & n4881 ) | ( ~n4646 & n4882 ) | ( n4881 & n4882 ) ;
  assign n4884 = ( n4646 & n4881 ) | ( n4646 & n4882 ) | ( n4881 & n4882 ) ;
  assign n4885 = ( n4646 & n4883 ) | ( n4646 & ~n4884 ) | ( n4883 & ~n4884 ) ;
  assign n4886 = ( x75 & n4880 ) | ( x75 & ~n4885 ) | ( n4880 & ~n4885 ) ;
  assign n4887 = ( x75 & n4647 ) | ( x75 & ~n4816 ) | ( n4647 & ~n4816 ) ;
  assign n4888 = x75 & n4647 ;
  assign n4889 = ( ~n4652 & n4887 ) | ( ~n4652 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4890 = ( n4652 & n4887 ) | ( n4652 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4891 = ( n4652 & n4889 ) | ( n4652 & ~n4890 ) | ( n4889 & ~n4890 ) ;
  assign n4892 = ( x76 & n4886 ) | ( x76 & ~n4891 ) | ( n4886 & ~n4891 ) ;
  assign n4893 = ( x76 & n4653 ) | ( x76 & ~n4816 ) | ( n4653 & ~n4816 ) ;
  assign n4894 = x76 & n4653 ;
  assign n4895 = ( ~n4658 & n4893 ) | ( ~n4658 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4896 = ( n4658 & n4893 ) | ( n4658 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4897 = ( n4658 & n4895 ) | ( n4658 & ~n4896 ) | ( n4895 & ~n4896 ) ;
  assign n4898 = ( x77 & n4892 ) | ( x77 & ~n4897 ) | ( n4892 & ~n4897 ) ;
  assign n4899 = ( x77 & n4659 ) | ( x77 & ~n4816 ) | ( n4659 & ~n4816 ) ;
  assign n4900 = x77 & n4659 ;
  assign n4901 = ( ~n4664 & n4899 ) | ( ~n4664 & n4900 ) | ( n4899 & n4900 ) ;
  assign n4902 = ( n4664 & n4899 ) | ( n4664 & n4900 ) | ( n4899 & n4900 ) ;
  assign n4903 = ( n4664 & n4901 ) | ( n4664 & ~n4902 ) | ( n4901 & ~n4902 ) ;
  assign n4904 = ( x78 & n4898 ) | ( x78 & ~n4903 ) | ( n4898 & ~n4903 ) ;
  assign n4905 = ( x78 & n4665 ) | ( x78 & ~n4816 ) | ( n4665 & ~n4816 ) ;
  assign n4906 = x78 & n4665 ;
  assign n4907 = ( ~n4670 & n4905 ) | ( ~n4670 & n4906 ) | ( n4905 & n4906 ) ;
  assign n4908 = ( n4670 & n4905 ) | ( n4670 & n4906 ) | ( n4905 & n4906 ) ;
  assign n4909 = ( n4670 & n4907 ) | ( n4670 & ~n4908 ) | ( n4907 & ~n4908 ) ;
  assign n4910 = ( x79 & n4904 ) | ( x79 & ~n4909 ) | ( n4904 & ~n4909 ) ;
  assign n4911 = ( x79 & n4671 ) | ( x79 & ~n4816 ) | ( n4671 & ~n4816 ) ;
  assign n4912 = x79 & n4671 ;
  assign n4913 = ( ~n4676 & n4911 ) | ( ~n4676 & n4912 ) | ( n4911 & n4912 ) ;
  assign n4914 = ( n4676 & n4911 ) | ( n4676 & n4912 ) | ( n4911 & n4912 ) ;
  assign n4915 = ( n4676 & n4913 ) | ( n4676 & ~n4914 ) | ( n4913 & ~n4914 ) ;
  assign n4916 = ( x80 & n4910 ) | ( x80 & ~n4915 ) | ( n4910 & ~n4915 ) ;
  assign n4917 = ( x80 & n4677 ) | ( x80 & ~n4816 ) | ( n4677 & ~n4816 ) ;
  assign n4918 = x80 & n4677 ;
  assign n4919 = ( ~n4682 & n4917 ) | ( ~n4682 & n4918 ) | ( n4917 & n4918 ) ;
  assign n4920 = ( n4682 & n4917 ) | ( n4682 & n4918 ) | ( n4917 & n4918 ) ;
  assign n4921 = ( n4682 & n4919 ) | ( n4682 & ~n4920 ) | ( n4919 & ~n4920 ) ;
  assign n4922 = ( x81 & n4916 ) | ( x81 & ~n4921 ) | ( n4916 & ~n4921 ) ;
  assign n4923 = ( x81 & n4683 ) | ( x81 & ~n4816 ) | ( n4683 & ~n4816 ) ;
  assign n4924 = x81 & n4683 ;
  assign n4925 = ( ~n4688 & n4923 ) | ( ~n4688 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4926 = ( n4688 & n4923 ) | ( n4688 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4927 = ( n4688 & n4925 ) | ( n4688 & ~n4926 ) | ( n4925 & ~n4926 ) ;
  assign n4928 = ( x82 & n4922 ) | ( x82 & ~n4927 ) | ( n4922 & ~n4927 ) ;
  assign n4929 = ( x82 & n4689 ) | ( x82 & ~n4816 ) | ( n4689 & ~n4816 ) ;
  assign n4930 = x82 & n4689 ;
  assign n4931 = ( ~n4694 & n4929 ) | ( ~n4694 & n4930 ) | ( n4929 & n4930 ) ;
  assign n4932 = ( n4694 & n4929 ) | ( n4694 & n4930 ) | ( n4929 & n4930 ) ;
  assign n4933 = ( n4694 & n4931 ) | ( n4694 & ~n4932 ) | ( n4931 & ~n4932 ) ;
  assign n4934 = ( x83 & n4928 ) | ( x83 & ~n4933 ) | ( n4928 & ~n4933 ) ;
  assign n4935 = ( x83 & n4695 ) | ( x83 & ~n4816 ) | ( n4695 & ~n4816 ) ;
  assign n4936 = x83 & n4695 ;
  assign n4937 = ( ~n4700 & n4935 ) | ( ~n4700 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4938 = ( n4700 & n4935 ) | ( n4700 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4939 = ( n4700 & n4937 ) | ( n4700 & ~n4938 ) | ( n4937 & ~n4938 ) ;
  assign n4940 = ( x84 & n4934 ) | ( x84 & ~n4939 ) | ( n4934 & ~n4939 ) ;
  assign n4941 = ( x84 & n4701 ) | ( x84 & ~n4816 ) | ( n4701 & ~n4816 ) ;
  assign n4942 = x84 & n4701 ;
  assign n4943 = ( ~n4706 & n4941 ) | ( ~n4706 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4944 = ( n4706 & n4941 ) | ( n4706 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4945 = ( n4706 & n4943 ) | ( n4706 & ~n4944 ) | ( n4943 & ~n4944 ) ;
  assign n4946 = ( x85 & n4940 ) | ( x85 & ~n4945 ) | ( n4940 & ~n4945 ) ;
  assign n4947 = ( x85 & n4707 ) | ( x85 & ~n4816 ) | ( n4707 & ~n4816 ) ;
  assign n4948 = x85 & n4707 ;
  assign n4949 = ( ~n4712 & n4947 ) | ( ~n4712 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4950 = ( n4712 & n4947 ) | ( n4712 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4951 = ( n4712 & n4949 ) | ( n4712 & ~n4950 ) | ( n4949 & ~n4950 ) ;
  assign n4952 = ( x86 & n4946 ) | ( x86 & ~n4951 ) | ( n4946 & ~n4951 ) ;
  assign n4953 = ( x86 & n4713 ) | ( x86 & ~n4816 ) | ( n4713 & ~n4816 ) ;
  assign n4954 = x86 & n4713 ;
  assign n4955 = ( ~n4718 & n4953 ) | ( ~n4718 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4956 = ( n4718 & n4953 ) | ( n4718 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4957 = ( n4718 & n4955 ) | ( n4718 & ~n4956 ) | ( n4955 & ~n4956 ) ;
  assign n4958 = ( x87 & n4952 ) | ( x87 & ~n4957 ) | ( n4952 & ~n4957 ) ;
  assign n4959 = ( x87 & n4719 ) | ( x87 & ~n4816 ) | ( n4719 & ~n4816 ) ;
  assign n4960 = x87 & n4719 ;
  assign n4961 = ( ~n4724 & n4959 ) | ( ~n4724 & n4960 ) | ( n4959 & n4960 ) ;
  assign n4962 = ( n4724 & n4959 ) | ( n4724 & n4960 ) | ( n4959 & n4960 ) ;
  assign n4963 = ( n4724 & n4961 ) | ( n4724 & ~n4962 ) | ( n4961 & ~n4962 ) ;
  assign n4964 = ( x88 & n4958 ) | ( x88 & ~n4963 ) | ( n4958 & ~n4963 ) ;
  assign n4965 = ( x88 & n4725 ) | ( x88 & ~n4816 ) | ( n4725 & ~n4816 ) ;
  assign n4966 = x88 & n4725 ;
  assign n4967 = ( ~n4730 & n4965 ) | ( ~n4730 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4968 = ( n4730 & n4965 ) | ( n4730 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4969 = ( n4730 & n4967 ) | ( n4730 & ~n4968 ) | ( n4967 & ~n4968 ) ;
  assign n4970 = ( x89 & n4964 ) | ( x89 & ~n4969 ) | ( n4964 & ~n4969 ) ;
  assign n4971 = ( x89 & n4731 ) | ( x89 & ~n4816 ) | ( n4731 & ~n4816 ) ;
  assign n4972 = x89 & n4731 ;
  assign n4973 = ( ~n4736 & n4971 ) | ( ~n4736 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = ( n4736 & n4971 ) | ( n4736 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4975 = ( n4736 & n4973 ) | ( n4736 & ~n4974 ) | ( n4973 & ~n4974 ) ;
  assign n4976 = ( x90 & n4970 ) | ( x90 & ~n4975 ) | ( n4970 & ~n4975 ) ;
  assign n4977 = ( x90 & n4737 ) | ( x90 & ~n4816 ) | ( n4737 & ~n4816 ) ;
  assign n4978 = x90 & n4737 ;
  assign n4979 = ( ~n4742 & n4977 ) | ( ~n4742 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4980 = ( n4742 & n4977 ) | ( n4742 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4981 = ( n4742 & n4979 ) | ( n4742 & ~n4980 ) | ( n4979 & ~n4980 ) ;
  assign n4982 = ( x91 & n4976 ) | ( x91 & ~n4981 ) | ( n4976 & ~n4981 ) ;
  assign n4983 = ( x91 & n4743 ) | ( x91 & ~n4816 ) | ( n4743 & ~n4816 ) ;
  assign n4984 = x91 & n4743 ;
  assign n4985 = ( ~n4748 & n4983 ) | ( ~n4748 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4986 = ( n4748 & n4983 ) | ( n4748 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4987 = ( n4748 & n4985 ) | ( n4748 & ~n4986 ) | ( n4985 & ~n4986 ) ;
  assign n4988 = ( x92 & n4982 ) | ( x92 & ~n4987 ) | ( n4982 & ~n4987 ) ;
  assign n4989 = ( x92 & n4749 ) | ( x92 & ~n4816 ) | ( n4749 & ~n4816 ) ;
  assign n4990 = x92 & n4749 ;
  assign n4991 = ( ~n4754 & n4989 ) | ( ~n4754 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = ( n4754 & n4989 ) | ( n4754 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4993 = ( n4754 & n4991 ) | ( n4754 & ~n4992 ) | ( n4991 & ~n4992 ) ;
  assign n4994 = ( x93 & n4988 ) | ( x93 & ~n4993 ) | ( n4988 & ~n4993 ) ;
  assign n4995 = ( x93 & n4755 ) | ( x93 & ~n4816 ) | ( n4755 & ~n4816 ) ;
  assign n4996 = x93 & n4755 ;
  assign n4997 = ( ~n4760 & n4995 ) | ( ~n4760 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4998 = ( n4760 & n4995 ) | ( n4760 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4999 = ( n4760 & n4997 ) | ( n4760 & ~n4998 ) | ( n4997 & ~n4998 ) ;
  assign n5000 = ( x94 & n4994 ) | ( x94 & ~n4999 ) | ( n4994 & ~n4999 ) ;
  assign n5001 = ( x94 & n4761 ) | ( x94 & ~n4816 ) | ( n4761 & ~n4816 ) ;
  assign n5002 = x94 & n4761 ;
  assign n5003 = ( ~n4766 & n5001 ) | ( ~n4766 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5004 = ( n4766 & n5001 ) | ( n4766 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5005 = ( n4766 & n5003 ) | ( n4766 & ~n5004 ) | ( n5003 & ~n5004 ) ;
  assign n5006 = ( x95 & n5000 ) | ( x95 & ~n5005 ) | ( n5000 & ~n5005 ) ;
  assign n5007 = ( x95 & n4767 ) | ( x95 & ~n4816 ) | ( n4767 & ~n4816 ) ;
  assign n5008 = x95 & n4767 ;
  assign n5009 = ( ~n4772 & n5007 ) | ( ~n4772 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5010 = ( n4772 & n5007 ) | ( n4772 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5011 = ( n4772 & n5009 ) | ( n4772 & ~n5010 ) | ( n5009 & ~n5010 ) ;
  assign n5012 = ( x96 & n5006 ) | ( x96 & ~n5011 ) | ( n5006 & ~n5011 ) ;
  assign n5013 = ( x96 & n4773 ) | ( x96 & ~n4816 ) | ( n4773 & ~n4816 ) ;
  assign n5014 = x96 & n4773 ;
  assign n5015 = ( ~n4778 & n5013 ) | ( ~n4778 & n5014 ) | ( n5013 & n5014 ) ;
  assign n5016 = ( n4778 & n5013 ) | ( n4778 & n5014 ) | ( n5013 & n5014 ) ;
  assign n5017 = ( n4778 & n5015 ) | ( n4778 & ~n5016 ) | ( n5015 & ~n5016 ) ;
  assign n5018 = ( x97 & n5012 ) | ( x97 & ~n5017 ) | ( n5012 & ~n5017 ) ;
  assign n5019 = ( x97 & n4779 ) | ( x97 & ~n4816 ) | ( n4779 & ~n4816 ) ;
  assign n5020 = x97 & n4779 ;
  assign n5021 = ( ~n4784 & n5019 ) | ( ~n4784 & n5020 ) | ( n5019 & n5020 ) ;
  assign n5022 = ( n4784 & n5019 ) | ( n4784 & n5020 ) | ( n5019 & n5020 ) ;
  assign n5023 = ( n4784 & n5021 ) | ( n4784 & ~n5022 ) | ( n5021 & ~n5022 ) ;
  assign n5024 = ( x98 & n5018 ) | ( x98 & ~n5023 ) | ( n5018 & ~n5023 ) ;
  assign n5025 = ( x98 & n4785 ) | ( x98 & ~n4816 ) | ( n4785 & ~n4816 ) ;
  assign n5026 = x98 & n4785 ;
  assign n5027 = ( ~n4790 & n5025 ) | ( ~n4790 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5028 = ( n4790 & n5025 ) | ( n4790 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5029 = ( n4790 & n5027 ) | ( n4790 & ~n5028 ) | ( n5027 & ~n5028 ) ;
  assign n5030 = ( x99 & n5024 ) | ( x99 & ~n5029 ) | ( n5024 & ~n5029 ) ;
  assign n5031 = ( x99 & n4791 ) | ( x99 & ~n4816 ) | ( n4791 & ~n4816 ) ;
  assign n5032 = x99 & n4791 ;
  assign n5033 = ( ~n4796 & n5031 ) | ( ~n4796 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5034 = ( n4796 & n5031 ) | ( n4796 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5035 = ( n4796 & n5033 ) | ( n4796 & ~n5034 ) | ( n5033 & ~n5034 ) ;
  assign n5036 = ( x100 & n5030 ) | ( x100 & ~n5035 ) | ( n5030 & ~n5035 ) ;
  assign n5037 = ( x100 & n4797 ) | ( x100 & ~n4816 ) | ( n4797 & ~n4816 ) ;
  assign n5038 = x100 & n4797 ;
  assign n5039 = ( ~n4802 & n5037 ) | ( ~n4802 & n5038 ) | ( n5037 & n5038 ) ;
  assign n5040 = ( n4802 & n5037 ) | ( n4802 & n5038 ) | ( n5037 & n5038 ) ;
  assign n5041 = ( n4802 & n5039 ) | ( n4802 & ~n5040 ) | ( n5039 & ~n5040 ) ;
  assign n5042 = ( x101 & n5036 ) | ( x101 & ~n5041 ) | ( n5036 & ~n5041 ) ;
  assign n5043 = ( x101 & n4803 ) | ( x101 & ~n4816 ) | ( n4803 & ~n4816 ) ;
  assign n5044 = x101 & n4803 ;
  assign n5045 = ( ~n4808 & n5043 ) | ( ~n4808 & n5044 ) | ( n5043 & n5044 ) ;
  assign n5046 = ( n4808 & n5043 ) | ( n4808 & n5044 ) | ( n5043 & n5044 ) ;
  assign n5047 = ( n4808 & n5045 ) | ( n4808 & ~n5046 ) | ( n5045 & ~n5046 ) ;
  assign n5048 = ( x102 & n5042 ) | ( x102 & ~n5047 ) | ( n5042 & ~n5047 ) ;
  assign n5049 = ( x103 & ~n153 ) | ( x103 & n4810 ) | ( ~n153 & n4810 ) ;
  assign n5050 = x103 & n4810 ;
  assign n5051 = ( n4814 & ~n5049 ) | ( n4814 & n5050 ) | ( ~n5049 & n5050 ) ;
  assign n5052 = ( x103 & ~n4821 ) | ( x103 & n5048 ) | ( ~n4821 & n5048 ) ;
  assign n5053 = ( x104 & ~n5051 ) | ( x104 & n5052 ) | ( ~n5051 & n5052 ) ;
  assign n5054 = n152 | n5053 ;
  assign n5055 = ( x103 & n5048 ) | ( x103 & n5054 ) | ( n5048 & n5054 ) ;
  assign n5056 = x103 | n5048 ;
  assign n5057 = ( ~n4821 & n5055 ) | ( ~n4821 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5058 = ( n4821 & n5055 ) | ( n4821 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5059 = ( n4821 & n5057 ) | ( n4821 & ~n5058 ) | ( n5057 & ~n5058 ) ;
  assign n5060 = ~x22 & x64 ;
  assign n5061 = ~x23 & n5054 ;
  assign n5062 = ( x23 & ~x64 ) | ( x23 & n5054 ) | ( ~x64 & n5054 ) ;
  assign n5063 = ( n4822 & ~n5061 ) | ( n4822 & n5062 ) | ( ~n5061 & n5062 ) ;
  assign n5064 = ( x65 & n5060 ) | ( x65 & ~n5063 ) | ( n5060 & ~n5063 ) ;
  assign n5065 = ( x65 & n4822 ) | ( x65 & n5054 ) | ( n4822 & n5054 ) ;
  assign n5066 = x65 | n4822 ;
  assign n5067 = ( ~n4825 & n5065 ) | ( ~n4825 & n5066 ) | ( n5065 & n5066 ) ;
  assign n5068 = ( n4825 & n5065 ) | ( n4825 & n5066 ) | ( n5065 & n5066 ) ;
  assign n5069 = ( n4825 & n5067 ) | ( n4825 & ~n5068 ) | ( n5067 & ~n5068 ) ;
  assign n5070 = ( x66 & n5064 ) | ( x66 & ~n5069 ) | ( n5064 & ~n5069 ) ;
  assign n5071 = ( x66 & n4826 ) | ( x66 & n5054 ) | ( n4826 & n5054 ) ;
  assign n5072 = x66 | n4826 ;
  assign n5073 = ( ~n4831 & n5071 ) | ( ~n4831 & n5072 ) | ( n5071 & n5072 ) ;
  assign n5074 = ( n4831 & n5071 ) | ( n4831 & n5072 ) | ( n5071 & n5072 ) ;
  assign n5075 = ( n4831 & n5073 ) | ( n4831 & ~n5074 ) | ( n5073 & ~n5074 ) ;
  assign n5076 = ( x67 & n5070 ) | ( x67 & ~n5075 ) | ( n5070 & ~n5075 ) ;
  assign n5077 = ( x67 & n4832 ) | ( x67 & ~n5054 ) | ( n4832 & ~n5054 ) ;
  assign n5078 = x67 & n4832 ;
  assign n5079 = ( ~n4837 & n5077 ) | ( ~n4837 & n5078 ) | ( n5077 & n5078 ) ;
  assign n5080 = ( n4837 & n5077 ) | ( n4837 & n5078 ) | ( n5077 & n5078 ) ;
  assign n5081 = ( n4837 & n5079 ) | ( n4837 & ~n5080 ) | ( n5079 & ~n5080 ) ;
  assign n5082 = ( x68 & n5076 ) | ( x68 & ~n5081 ) | ( n5076 & ~n5081 ) ;
  assign n5083 = ( x68 & n4838 ) | ( x68 & ~n5054 ) | ( n4838 & ~n5054 ) ;
  assign n5084 = x68 & n4838 ;
  assign n5085 = ( ~n4843 & n5083 ) | ( ~n4843 & n5084 ) | ( n5083 & n5084 ) ;
  assign n5086 = ( n4843 & n5083 ) | ( n4843 & n5084 ) | ( n5083 & n5084 ) ;
  assign n5087 = ( n4843 & n5085 ) | ( n4843 & ~n5086 ) | ( n5085 & ~n5086 ) ;
  assign n5088 = ( x69 & n5082 ) | ( x69 & ~n5087 ) | ( n5082 & ~n5087 ) ;
  assign n5089 = ( x69 & n4844 ) | ( x69 & ~n5054 ) | ( n4844 & ~n5054 ) ;
  assign n5090 = x69 & n4844 ;
  assign n5091 = ( ~n4849 & n5089 ) | ( ~n4849 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5092 = ( n4849 & n5089 ) | ( n4849 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5093 = ( n4849 & n5091 ) | ( n4849 & ~n5092 ) | ( n5091 & ~n5092 ) ;
  assign n5094 = ( x70 & n5088 ) | ( x70 & ~n5093 ) | ( n5088 & ~n5093 ) ;
  assign n5095 = ( x70 & n4850 ) | ( x70 & ~n5054 ) | ( n4850 & ~n5054 ) ;
  assign n5096 = x70 & n4850 ;
  assign n5097 = ( ~n4855 & n5095 ) | ( ~n4855 & n5096 ) | ( n5095 & n5096 ) ;
  assign n5098 = ( n4855 & n5095 ) | ( n4855 & n5096 ) | ( n5095 & n5096 ) ;
  assign n5099 = ( n4855 & n5097 ) | ( n4855 & ~n5098 ) | ( n5097 & ~n5098 ) ;
  assign n5100 = ( x71 & n5094 ) | ( x71 & ~n5099 ) | ( n5094 & ~n5099 ) ;
  assign n5101 = ( x71 & n4856 ) | ( x71 & ~n5054 ) | ( n4856 & ~n5054 ) ;
  assign n5102 = x71 & n4856 ;
  assign n5103 = ( ~n4861 & n5101 ) | ( ~n4861 & n5102 ) | ( n5101 & n5102 ) ;
  assign n5104 = ( n4861 & n5101 ) | ( n4861 & n5102 ) | ( n5101 & n5102 ) ;
  assign n5105 = ( n4861 & n5103 ) | ( n4861 & ~n5104 ) | ( n5103 & ~n5104 ) ;
  assign n5106 = ( x72 & n5100 ) | ( x72 & ~n5105 ) | ( n5100 & ~n5105 ) ;
  assign n5107 = ( x72 & n4862 ) | ( x72 & ~n5054 ) | ( n4862 & ~n5054 ) ;
  assign n5108 = x72 & n4862 ;
  assign n5109 = ( ~n4867 & n5107 ) | ( ~n4867 & n5108 ) | ( n5107 & n5108 ) ;
  assign n5110 = ( n4867 & n5107 ) | ( n4867 & n5108 ) | ( n5107 & n5108 ) ;
  assign n5111 = ( n4867 & n5109 ) | ( n4867 & ~n5110 ) | ( n5109 & ~n5110 ) ;
  assign n5112 = ( x73 & n5106 ) | ( x73 & ~n5111 ) | ( n5106 & ~n5111 ) ;
  assign n5113 = ( x73 & n4868 ) | ( x73 & ~n5054 ) | ( n4868 & ~n5054 ) ;
  assign n5114 = x73 & n4868 ;
  assign n5115 = ( ~n4873 & n5113 ) | ( ~n4873 & n5114 ) | ( n5113 & n5114 ) ;
  assign n5116 = ( n4873 & n5113 ) | ( n4873 & n5114 ) | ( n5113 & n5114 ) ;
  assign n5117 = ( n4873 & n5115 ) | ( n4873 & ~n5116 ) | ( n5115 & ~n5116 ) ;
  assign n5118 = ( x74 & n5112 ) | ( x74 & ~n5117 ) | ( n5112 & ~n5117 ) ;
  assign n5119 = ( x74 & n4874 ) | ( x74 & ~n5054 ) | ( n4874 & ~n5054 ) ;
  assign n5120 = x74 & n4874 ;
  assign n5121 = ( ~n4879 & n5119 ) | ( ~n4879 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5122 = ( n4879 & n5119 ) | ( n4879 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5123 = ( n4879 & n5121 ) | ( n4879 & ~n5122 ) | ( n5121 & ~n5122 ) ;
  assign n5124 = ( x75 & n5118 ) | ( x75 & ~n5123 ) | ( n5118 & ~n5123 ) ;
  assign n5125 = ( x75 & n4880 ) | ( x75 & ~n5054 ) | ( n4880 & ~n5054 ) ;
  assign n5126 = x75 & n4880 ;
  assign n5127 = ( ~n4885 & n5125 ) | ( ~n4885 & n5126 ) | ( n5125 & n5126 ) ;
  assign n5128 = ( n4885 & n5125 ) | ( n4885 & n5126 ) | ( n5125 & n5126 ) ;
  assign n5129 = ( n4885 & n5127 ) | ( n4885 & ~n5128 ) | ( n5127 & ~n5128 ) ;
  assign n5130 = ( x76 & n5124 ) | ( x76 & ~n5129 ) | ( n5124 & ~n5129 ) ;
  assign n5131 = ( x76 & n4886 ) | ( x76 & ~n5054 ) | ( n4886 & ~n5054 ) ;
  assign n5132 = x76 & n4886 ;
  assign n5133 = ( ~n4891 & n5131 ) | ( ~n4891 & n5132 ) | ( n5131 & n5132 ) ;
  assign n5134 = ( n4891 & n5131 ) | ( n4891 & n5132 ) | ( n5131 & n5132 ) ;
  assign n5135 = ( n4891 & n5133 ) | ( n4891 & ~n5134 ) | ( n5133 & ~n5134 ) ;
  assign n5136 = ( x77 & n5130 ) | ( x77 & ~n5135 ) | ( n5130 & ~n5135 ) ;
  assign n5137 = ( x77 & n4892 ) | ( x77 & ~n5054 ) | ( n4892 & ~n5054 ) ;
  assign n5138 = x77 & n4892 ;
  assign n5139 = ( ~n4897 & n5137 ) | ( ~n4897 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5140 = ( n4897 & n5137 ) | ( n4897 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5141 = ( n4897 & n5139 ) | ( n4897 & ~n5140 ) | ( n5139 & ~n5140 ) ;
  assign n5142 = ( x78 & n5136 ) | ( x78 & ~n5141 ) | ( n5136 & ~n5141 ) ;
  assign n5143 = ( x78 & n4898 ) | ( x78 & ~n5054 ) | ( n4898 & ~n5054 ) ;
  assign n5144 = x78 & n4898 ;
  assign n5145 = ( ~n4903 & n5143 ) | ( ~n4903 & n5144 ) | ( n5143 & n5144 ) ;
  assign n5146 = ( n4903 & n5143 ) | ( n4903 & n5144 ) | ( n5143 & n5144 ) ;
  assign n5147 = ( n4903 & n5145 ) | ( n4903 & ~n5146 ) | ( n5145 & ~n5146 ) ;
  assign n5148 = ( x79 & n5142 ) | ( x79 & ~n5147 ) | ( n5142 & ~n5147 ) ;
  assign n5149 = ( x79 & n4904 ) | ( x79 & ~n5054 ) | ( n4904 & ~n5054 ) ;
  assign n5150 = x79 & n4904 ;
  assign n5151 = ( ~n4909 & n5149 ) | ( ~n4909 & n5150 ) | ( n5149 & n5150 ) ;
  assign n5152 = ( n4909 & n5149 ) | ( n4909 & n5150 ) | ( n5149 & n5150 ) ;
  assign n5153 = ( n4909 & n5151 ) | ( n4909 & ~n5152 ) | ( n5151 & ~n5152 ) ;
  assign n5154 = ( x80 & n5148 ) | ( x80 & ~n5153 ) | ( n5148 & ~n5153 ) ;
  assign n5155 = ( x80 & n4910 ) | ( x80 & ~n5054 ) | ( n4910 & ~n5054 ) ;
  assign n5156 = x80 & n4910 ;
  assign n5157 = ( ~n4915 & n5155 ) | ( ~n4915 & n5156 ) | ( n5155 & n5156 ) ;
  assign n5158 = ( n4915 & n5155 ) | ( n4915 & n5156 ) | ( n5155 & n5156 ) ;
  assign n5159 = ( n4915 & n5157 ) | ( n4915 & ~n5158 ) | ( n5157 & ~n5158 ) ;
  assign n5160 = ( x81 & n5154 ) | ( x81 & ~n5159 ) | ( n5154 & ~n5159 ) ;
  assign n5161 = ( x81 & n4916 ) | ( x81 & ~n5054 ) | ( n4916 & ~n5054 ) ;
  assign n5162 = x81 & n4916 ;
  assign n5163 = ( ~n4921 & n5161 ) | ( ~n4921 & n5162 ) | ( n5161 & n5162 ) ;
  assign n5164 = ( n4921 & n5161 ) | ( n4921 & n5162 ) | ( n5161 & n5162 ) ;
  assign n5165 = ( n4921 & n5163 ) | ( n4921 & ~n5164 ) | ( n5163 & ~n5164 ) ;
  assign n5166 = ( x82 & n5160 ) | ( x82 & ~n5165 ) | ( n5160 & ~n5165 ) ;
  assign n5167 = ( x82 & n4922 ) | ( x82 & ~n5054 ) | ( n4922 & ~n5054 ) ;
  assign n5168 = x82 & n4922 ;
  assign n5169 = ( ~n4927 & n5167 ) | ( ~n4927 & n5168 ) | ( n5167 & n5168 ) ;
  assign n5170 = ( n4927 & n5167 ) | ( n4927 & n5168 ) | ( n5167 & n5168 ) ;
  assign n5171 = ( n4927 & n5169 ) | ( n4927 & ~n5170 ) | ( n5169 & ~n5170 ) ;
  assign n5172 = ( x83 & n5166 ) | ( x83 & ~n5171 ) | ( n5166 & ~n5171 ) ;
  assign n5173 = ( x83 & n4928 ) | ( x83 & ~n5054 ) | ( n4928 & ~n5054 ) ;
  assign n5174 = x83 & n4928 ;
  assign n5175 = ( ~n4933 & n5173 ) | ( ~n4933 & n5174 ) | ( n5173 & n5174 ) ;
  assign n5176 = ( n4933 & n5173 ) | ( n4933 & n5174 ) | ( n5173 & n5174 ) ;
  assign n5177 = ( n4933 & n5175 ) | ( n4933 & ~n5176 ) | ( n5175 & ~n5176 ) ;
  assign n5178 = ( x84 & n5172 ) | ( x84 & ~n5177 ) | ( n5172 & ~n5177 ) ;
  assign n5179 = ( x84 & n4934 ) | ( x84 & ~n5054 ) | ( n4934 & ~n5054 ) ;
  assign n5180 = x84 & n4934 ;
  assign n5181 = ( ~n4939 & n5179 ) | ( ~n4939 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5182 = ( n4939 & n5179 ) | ( n4939 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5183 = ( n4939 & n5181 ) | ( n4939 & ~n5182 ) | ( n5181 & ~n5182 ) ;
  assign n5184 = ( x85 & n5178 ) | ( x85 & ~n5183 ) | ( n5178 & ~n5183 ) ;
  assign n5185 = ( x85 & n4940 ) | ( x85 & ~n5054 ) | ( n4940 & ~n5054 ) ;
  assign n5186 = x85 & n4940 ;
  assign n5187 = ( ~n4945 & n5185 ) | ( ~n4945 & n5186 ) | ( n5185 & n5186 ) ;
  assign n5188 = ( n4945 & n5185 ) | ( n4945 & n5186 ) | ( n5185 & n5186 ) ;
  assign n5189 = ( n4945 & n5187 ) | ( n4945 & ~n5188 ) | ( n5187 & ~n5188 ) ;
  assign n5190 = ( x86 & n5184 ) | ( x86 & ~n5189 ) | ( n5184 & ~n5189 ) ;
  assign n5191 = ( x86 & n4946 ) | ( x86 & ~n5054 ) | ( n4946 & ~n5054 ) ;
  assign n5192 = x86 & n4946 ;
  assign n5193 = ( ~n4951 & n5191 ) | ( ~n4951 & n5192 ) | ( n5191 & n5192 ) ;
  assign n5194 = ( n4951 & n5191 ) | ( n4951 & n5192 ) | ( n5191 & n5192 ) ;
  assign n5195 = ( n4951 & n5193 ) | ( n4951 & ~n5194 ) | ( n5193 & ~n5194 ) ;
  assign n5196 = ( x87 & n5190 ) | ( x87 & ~n5195 ) | ( n5190 & ~n5195 ) ;
  assign n5197 = ( x87 & n4952 ) | ( x87 & ~n5054 ) | ( n4952 & ~n5054 ) ;
  assign n5198 = x87 & n4952 ;
  assign n5199 = ( ~n4957 & n5197 ) | ( ~n4957 & n5198 ) | ( n5197 & n5198 ) ;
  assign n5200 = ( n4957 & n5197 ) | ( n4957 & n5198 ) | ( n5197 & n5198 ) ;
  assign n5201 = ( n4957 & n5199 ) | ( n4957 & ~n5200 ) | ( n5199 & ~n5200 ) ;
  assign n5202 = ( x88 & n5196 ) | ( x88 & ~n5201 ) | ( n5196 & ~n5201 ) ;
  assign n5203 = ( x88 & n4958 ) | ( x88 & ~n5054 ) | ( n4958 & ~n5054 ) ;
  assign n5204 = x88 & n4958 ;
  assign n5205 = ( ~n4963 & n5203 ) | ( ~n4963 & n5204 ) | ( n5203 & n5204 ) ;
  assign n5206 = ( n4963 & n5203 ) | ( n4963 & n5204 ) | ( n5203 & n5204 ) ;
  assign n5207 = ( n4963 & n5205 ) | ( n4963 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = ( x89 & n5202 ) | ( x89 & ~n5207 ) | ( n5202 & ~n5207 ) ;
  assign n5209 = ( x89 & n4964 ) | ( x89 & ~n5054 ) | ( n4964 & ~n5054 ) ;
  assign n5210 = x89 & n4964 ;
  assign n5211 = ( ~n4969 & n5209 ) | ( ~n4969 & n5210 ) | ( n5209 & n5210 ) ;
  assign n5212 = ( n4969 & n5209 ) | ( n4969 & n5210 ) | ( n5209 & n5210 ) ;
  assign n5213 = ( n4969 & n5211 ) | ( n4969 & ~n5212 ) | ( n5211 & ~n5212 ) ;
  assign n5214 = ( x90 & n5208 ) | ( x90 & ~n5213 ) | ( n5208 & ~n5213 ) ;
  assign n5215 = ( x90 & n4970 ) | ( x90 & ~n5054 ) | ( n4970 & ~n5054 ) ;
  assign n5216 = x90 & n4970 ;
  assign n5217 = ( ~n4975 & n5215 ) | ( ~n4975 & n5216 ) | ( n5215 & n5216 ) ;
  assign n5218 = ( n4975 & n5215 ) | ( n4975 & n5216 ) | ( n5215 & n5216 ) ;
  assign n5219 = ( n4975 & n5217 ) | ( n4975 & ~n5218 ) | ( n5217 & ~n5218 ) ;
  assign n5220 = ( x91 & n5214 ) | ( x91 & ~n5219 ) | ( n5214 & ~n5219 ) ;
  assign n5221 = ( x91 & n4976 ) | ( x91 & ~n5054 ) | ( n4976 & ~n5054 ) ;
  assign n5222 = x91 & n4976 ;
  assign n5223 = ( ~n4981 & n5221 ) | ( ~n4981 & n5222 ) | ( n5221 & n5222 ) ;
  assign n5224 = ( n4981 & n5221 ) | ( n4981 & n5222 ) | ( n5221 & n5222 ) ;
  assign n5225 = ( n4981 & n5223 ) | ( n4981 & ~n5224 ) | ( n5223 & ~n5224 ) ;
  assign n5226 = ( x92 & n5220 ) | ( x92 & ~n5225 ) | ( n5220 & ~n5225 ) ;
  assign n5227 = ( x92 & n4982 ) | ( x92 & ~n5054 ) | ( n4982 & ~n5054 ) ;
  assign n5228 = x92 & n4982 ;
  assign n5229 = ( ~n4987 & n5227 ) | ( ~n4987 & n5228 ) | ( n5227 & n5228 ) ;
  assign n5230 = ( n4987 & n5227 ) | ( n4987 & n5228 ) | ( n5227 & n5228 ) ;
  assign n5231 = ( n4987 & n5229 ) | ( n4987 & ~n5230 ) | ( n5229 & ~n5230 ) ;
  assign n5232 = ( x93 & n5226 ) | ( x93 & ~n5231 ) | ( n5226 & ~n5231 ) ;
  assign n5233 = ( x93 & n4988 ) | ( x93 & ~n5054 ) | ( n4988 & ~n5054 ) ;
  assign n5234 = x93 & n4988 ;
  assign n5235 = ( ~n4993 & n5233 ) | ( ~n4993 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5236 = ( n4993 & n5233 ) | ( n4993 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5237 = ( n4993 & n5235 ) | ( n4993 & ~n5236 ) | ( n5235 & ~n5236 ) ;
  assign n5238 = ( x94 & n5232 ) | ( x94 & ~n5237 ) | ( n5232 & ~n5237 ) ;
  assign n5239 = ( x94 & n4994 ) | ( x94 & ~n5054 ) | ( n4994 & ~n5054 ) ;
  assign n5240 = x94 & n4994 ;
  assign n5241 = ( ~n4999 & n5239 ) | ( ~n4999 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5242 = ( n4999 & n5239 ) | ( n4999 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5243 = ( n4999 & n5241 ) | ( n4999 & ~n5242 ) | ( n5241 & ~n5242 ) ;
  assign n5244 = ( x95 & n5238 ) | ( x95 & ~n5243 ) | ( n5238 & ~n5243 ) ;
  assign n5245 = ( x95 & n5000 ) | ( x95 & ~n5054 ) | ( n5000 & ~n5054 ) ;
  assign n5246 = x95 & n5000 ;
  assign n5247 = ( ~n5005 & n5245 ) | ( ~n5005 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5248 = ( n5005 & n5245 ) | ( n5005 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5249 = ( n5005 & n5247 ) | ( n5005 & ~n5248 ) | ( n5247 & ~n5248 ) ;
  assign n5250 = ( x96 & n5244 ) | ( x96 & ~n5249 ) | ( n5244 & ~n5249 ) ;
  assign n5251 = ( x96 & n5006 ) | ( x96 & ~n5054 ) | ( n5006 & ~n5054 ) ;
  assign n5252 = x96 & n5006 ;
  assign n5253 = ( ~n5011 & n5251 ) | ( ~n5011 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5254 = ( n5011 & n5251 ) | ( n5011 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5255 = ( n5011 & n5253 ) | ( n5011 & ~n5254 ) | ( n5253 & ~n5254 ) ;
  assign n5256 = ( x97 & n5250 ) | ( x97 & ~n5255 ) | ( n5250 & ~n5255 ) ;
  assign n5257 = ( x97 & n5012 ) | ( x97 & ~n5054 ) | ( n5012 & ~n5054 ) ;
  assign n5258 = x97 & n5012 ;
  assign n5259 = ( ~n5017 & n5257 ) | ( ~n5017 & n5258 ) | ( n5257 & n5258 ) ;
  assign n5260 = ( n5017 & n5257 ) | ( n5017 & n5258 ) | ( n5257 & n5258 ) ;
  assign n5261 = ( n5017 & n5259 ) | ( n5017 & ~n5260 ) | ( n5259 & ~n5260 ) ;
  assign n5262 = ( x98 & n5256 ) | ( x98 & ~n5261 ) | ( n5256 & ~n5261 ) ;
  assign n5263 = ( x98 & n5018 ) | ( x98 & ~n5054 ) | ( n5018 & ~n5054 ) ;
  assign n5264 = x98 & n5018 ;
  assign n5265 = ( ~n5023 & n5263 ) | ( ~n5023 & n5264 ) | ( n5263 & n5264 ) ;
  assign n5266 = ( n5023 & n5263 ) | ( n5023 & n5264 ) | ( n5263 & n5264 ) ;
  assign n5267 = ( n5023 & n5265 ) | ( n5023 & ~n5266 ) | ( n5265 & ~n5266 ) ;
  assign n5268 = ( x99 & n5262 ) | ( x99 & ~n5267 ) | ( n5262 & ~n5267 ) ;
  assign n5269 = ( x99 & n5024 ) | ( x99 & ~n5054 ) | ( n5024 & ~n5054 ) ;
  assign n5270 = x99 & n5024 ;
  assign n5271 = ( ~n5029 & n5269 ) | ( ~n5029 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5272 = ( n5029 & n5269 ) | ( n5029 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5273 = ( n5029 & n5271 ) | ( n5029 & ~n5272 ) | ( n5271 & ~n5272 ) ;
  assign n5274 = ( x100 & n5268 ) | ( x100 & ~n5273 ) | ( n5268 & ~n5273 ) ;
  assign n5275 = ( x100 & n5030 ) | ( x100 & ~n5054 ) | ( n5030 & ~n5054 ) ;
  assign n5276 = x100 & n5030 ;
  assign n5277 = ( ~n5035 & n5275 ) | ( ~n5035 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5278 = ( n5035 & n5275 ) | ( n5035 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5279 = ( n5035 & n5277 ) | ( n5035 & ~n5278 ) | ( n5277 & ~n5278 ) ;
  assign n5280 = ( x101 & n5274 ) | ( x101 & ~n5279 ) | ( n5274 & ~n5279 ) ;
  assign n5281 = ( x101 & n5036 ) | ( x101 & ~n5054 ) | ( n5036 & ~n5054 ) ;
  assign n5282 = x101 & n5036 ;
  assign n5283 = ( ~n5041 & n5281 ) | ( ~n5041 & n5282 ) | ( n5281 & n5282 ) ;
  assign n5284 = ( n5041 & n5281 ) | ( n5041 & n5282 ) | ( n5281 & n5282 ) ;
  assign n5285 = ( n5041 & n5283 ) | ( n5041 & ~n5284 ) | ( n5283 & ~n5284 ) ;
  assign n5286 = ( x102 & n5280 ) | ( x102 & ~n5285 ) | ( n5280 & ~n5285 ) ;
  assign n5287 = ( x102 & n5042 ) | ( x102 & ~n5054 ) | ( n5042 & ~n5054 ) ;
  assign n5288 = x102 & n5042 ;
  assign n5289 = ( ~n5047 & n5287 ) | ( ~n5047 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5290 = ( n5047 & n5287 ) | ( n5047 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5291 = ( n5047 & n5289 ) | ( n5047 & ~n5290 ) | ( n5289 & ~n5290 ) ;
  assign n5292 = ( x103 & n5286 ) | ( x103 & ~n5291 ) | ( n5286 & ~n5291 ) ;
  assign n5293 = ( n151 & n152 ) | ( n151 & ~n5051 ) | ( n152 & ~n5051 ) ;
  assign n5294 = ( x104 & ~n5059 ) | ( x104 & n5292 ) | ( ~n5059 & n5292 ) ;
  assign n5295 = n5293 | n5294 ;
  assign n5296 = ( ~x104 & n152 ) | ( ~x104 & n5052 ) | ( n152 & n5052 ) ;
  assign n5297 = ( ~x104 & n5051 ) | ( ~x104 & n5052 ) | ( n5051 & n5052 ) ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = n5295 & ~n5298 ;
  assign n5300 = ( x104 & n5292 ) | ( x104 & ~n5299 ) | ( n5292 & ~n5299 ) ;
  assign n5301 = x104 & n5292 ;
  assign n5302 = ( ~n5059 & n5300 ) | ( ~n5059 & n5301 ) | ( n5300 & n5301 ) ;
  assign n5303 = ( n5059 & n5300 ) | ( n5059 & n5301 ) | ( n5300 & n5301 ) ;
  assign n5304 = ( n5059 & n5302 ) | ( n5059 & ~n5303 ) | ( n5302 & ~n5303 ) ;
  assign n5305 = ~x21 & x64 ;
  assign n5306 = x22 & n5299 ;
  assign n5307 = ( x22 & x64 ) | ( x22 & ~n5299 ) | ( x64 & ~n5299 ) ;
  assign n5308 = x22 & x64 ;
  assign n5309 = ( n5306 & n5307 ) | ( n5306 & ~n5308 ) | ( n5307 & ~n5308 ) ;
  assign n5310 = ( x65 & n5305 ) | ( x65 & ~n5309 ) | ( n5305 & ~n5309 ) ;
  assign n5311 = ( x65 & n5060 ) | ( x65 & n5299 ) | ( n5060 & n5299 ) ;
  assign n5312 = x65 | n5060 ;
  assign n5313 = ( ~n5063 & n5311 ) | ( ~n5063 & n5312 ) | ( n5311 & n5312 ) ;
  assign n5314 = ( n5063 & n5311 ) | ( n5063 & n5312 ) | ( n5311 & n5312 ) ;
  assign n5315 = ( n5063 & n5313 ) | ( n5063 & ~n5314 ) | ( n5313 & ~n5314 ) ;
  assign n5316 = ( x66 & n5310 ) | ( x66 & ~n5315 ) | ( n5310 & ~n5315 ) ;
  assign n5317 = ( x66 & n5064 ) | ( x66 & n5299 ) | ( n5064 & n5299 ) ;
  assign n5318 = x66 | n5064 ;
  assign n5319 = ( ~n5069 & n5317 ) | ( ~n5069 & n5318 ) | ( n5317 & n5318 ) ;
  assign n5320 = ( n5069 & n5317 ) | ( n5069 & n5318 ) | ( n5317 & n5318 ) ;
  assign n5321 = ( n5069 & n5319 ) | ( n5069 & ~n5320 ) | ( n5319 & ~n5320 ) ;
  assign n5322 = ( x67 & n5316 ) | ( x67 & ~n5321 ) | ( n5316 & ~n5321 ) ;
  assign n5323 = ( x67 & n5070 ) | ( x67 & ~n5299 ) | ( n5070 & ~n5299 ) ;
  assign n5324 = x67 & n5070 ;
  assign n5325 = ( ~n5075 & n5323 ) | ( ~n5075 & n5324 ) | ( n5323 & n5324 ) ;
  assign n5326 = ( n5075 & n5323 ) | ( n5075 & n5324 ) | ( n5323 & n5324 ) ;
  assign n5327 = ( n5075 & n5325 ) | ( n5075 & ~n5326 ) | ( n5325 & ~n5326 ) ;
  assign n5328 = ( x68 & n5322 ) | ( x68 & ~n5327 ) | ( n5322 & ~n5327 ) ;
  assign n5329 = ( x68 & n5076 ) | ( x68 & ~n5299 ) | ( n5076 & ~n5299 ) ;
  assign n5330 = x68 & n5076 ;
  assign n5331 = ( ~n5081 & n5329 ) | ( ~n5081 & n5330 ) | ( n5329 & n5330 ) ;
  assign n5332 = ( n5081 & n5329 ) | ( n5081 & n5330 ) | ( n5329 & n5330 ) ;
  assign n5333 = ( n5081 & n5331 ) | ( n5081 & ~n5332 ) | ( n5331 & ~n5332 ) ;
  assign n5334 = ( x69 & n5328 ) | ( x69 & ~n5333 ) | ( n5328 & ~n5333 ) ;
  assign n5335 = ( x69 & n5082 ) | ( x69 & ~n5299 ) | ( n5082 & ~n5299 ) ;
  assign n5336 = x69 & n5082 ;
  assign n5337 = ( ~n5087 & n5335 ) | ( ~n5087 & n5336 ) | ( n5335 & n5336 ) ;
  assign n5338 = ( n5087 & n5335 ) | ( n5087 & n5336 ) | ( n5335 & n5336 ) ;
  assign n5339 = ( n5087 & n5337 ) | ( n5087 & ~n5338 ) | ( n5337 & ~n5338 ) ;
  assign n5340 = ( x70 & n5334 ) | ( x70 & ~n5339 ) | ( n5334 & ~n5339 ) ;
  assign n5341 = ( x70 & n5088 ) | ( x70 & ~n5299 ) | ( n5088 & ~n5299 ) ;
  assign n5342 = x70 & n5088 ;
  assign n5343 = ( ~n5093 & n5341 ) | ( ~n5093 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = ( n5093 & n5341 ) | ( n5093 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5345 = ( n5093 & n5343 ) | ( n5093 & ~n5344 ) | ( n5343 & ~n5344 ) ;
  assign n5346 = ( x71 & n5340 ) | ( x71 & ~n5345 ) | ( n5340 & ~n5345 ) ;
  assign n5347 = ( x71 & n5094 ) | ( x71 & ~n5299 ) | ( n5094 & ~n5299 ) ;
  assign n5348 = x71 & n5094 ;
  assign n5349 = ( ~n5099 & n5347 ) | ( ~n5099 & n5348 ) | ( n5347 & n5348 ) ;
  assign n5350 = ( n5099 & n5347 ) | ( n5099 & n5348 ) | ( n5347 & n5348 ) ;
  assign n5351 = ( n5099 & n5349 ) | ( n5099 & ~n5350 ) | ( n5349 & ~n5350 ) ;
  assign n5352 = ( x72 & n5346 ) | ( x72 & ~n5351 ) | ( n5346 & ~n5351 ) ;
  assign n5353 = ( x72 & n5100 ) | ( x72 & ~n5299 ) | ( n5100 & ~n5299 ) ;
  assign n5354 = x72 & n5100 ;
  assign n5355 = ( ~n5105 & n5353 ) | ( ~n5105 & n5354 ) | ( n5353 & n5354 ) ;
  assign n5356 = ( n5105 & n5353 ) | ( n5105 & n5354 ) | ( n5353 & n5354 ) ;
  assign n5357 = ( n5105 & n5355 ) | ( n5105 & ~n5356 ) | ( n5355 & ~n5356 ) ;
  assign n5358 = ( x73 & n5352 ) | ( x73 & ~n5357 ) | ( n5352 & ~n5357 ) ;
  assign n5359 = ( x73 & n5106 ) | ( x73 & ~n5299 ) | ( n5106 & ~n5299 ) ;
  assign n5360 = x73 & n5106 ;
  assign n5361 = ( ~n5111 & n5359 ) | ( ~n5111 & n5360 ) | ( n5359 & n5360 ) ;
  assign n5362 = ( n5111 & n5359 ) | ( n5111 & n5360 ) | ( n5359 & n5360 ) ;
  assign n5363 = ( n5111 & n5361 ) | ( n5111 & ~n5362 ) | ( n5361 & ~n5362 ) ;
  assign n5364 = ( x74 & n5358 ) | ( x74 & ~n5363 ) | ( n5358 & ~n5363 ) ;
  assign n5365 = ( x74 & n5112 ) | ( x74 & ~n5299 ) | ( n5112 & ~n5299 ) ;
  assign n5366 = x74 & n5112 ;
  assign n5367 = ( ~n5117 & n5365 ) | ( ~n5117 & n5366 ) | ( n5365 & n5366 ) ;
  assign n5368 = ( n5117 & n5365 ) | ( n5117 & n5366 ) | ( n5365 & n5366 ) ;
  assign n5369 = ( n5117 & n5367 ) | ( n5117 & ~n5368 ) | ( n5367 & ~n5368 ) ;
  assign n5370 = ( x75 & n5364 ) | ( x75 & ~n5369 ) | ( n5364 & ~n5369 ) ;
  assign n5371 = ( x75 & n5118 ) | ( x75 & ~n5299 ) | ( n5118 & ~n5299 ) ;
  assign n5372 = x75 & n5118 ;
  assign n5373 = ( ~n5123 & n5371 ) | ( ~n5123 & n5372 ) | ( n5371 & n5372 ) ;
  assign n5374 = ( n5123 & n5371 ) | ( n5123 & n5372 ) | ( n5371 & n5372 ) ;
  assign n5375 = ( n5123 & n5373 ) | ( n5123 & ~n5374 ) | ( n5373 & ~n5374 ) ;
  assign n5376 = ( x76 & n5370 ) | ( x76 & ~n5375 ) | ( n5370 & ~n5375 ) ;
  assign n5377 = ( x76 & n5124 ) | ( x76 & ~n5299 ) | ( n5124 & ~n5299 ) ;
  assign n5378 = x76 & n5124 ;
  assign n5379 = ( ~n5129 & n5377 ) | ( ~n5129 & n5378 ) | ( n5377 & n5378 ) ;
  assign n5380 = ( n5129 & n5377 ) | ( n5129 & n5378 ) | ( n5377 & n5378 ) ;
  assign n5381 = ( n5129 & n5379 ) | ( n5129 & ~n5380 ) | ( n5379 & ~n5380 ) ;
  assign n5382 = ( x77 & n5376 ) | ( x77 & ~n5381 ) | ( n5376 & ~n5381 ) ;
  assign n5383 = ( x77 & n5130 ) | ( x77 & ~n5299 ) | ( n5130 & ~n5299 ) ;
  assign n5384 = x77 & n5130 ;
  assign n5385 = ( ~n5135 & n5383 ) | ( ~n5135 & n5384 ) | ( n5383 & n5384 ) ;
  assign n5386 = ( n5135 & n5383 ) | ( n5135 & n5384 ) | ( n5383 & n5384 ) ;
  assign n5387 = ( n5135 & n5385 ) | ( n5135 & ~n5386 ) | ( n5385 & ~n5386 ) ;
  assign n5388 = ( x78 & n5382 ) | ( x78 & ~n5387 ) | ( n5382 & ~n5387 ) ;
  assign n5389 = ( x78 & n5136 ) | ( x78 & ~n5299 ) | ( n5136 & ~n5299 ) ;
  assign n5390 = x78 & n5136 ;
  assign n5391 = ( ~n5141 & n5389 ) | ( ~n5141 & n5390 ) | ( n5389 & n5390 ) ;
  assign n5392 = ( n5141 & n5389 ) | ( n5141 & n5390 ) | ( n5389 & n5390 ) ;
  assign n5393 = ( n5141 & n5391 ) | ( n5141 & ~n5392 ) | ( n5391 & ~n5392 ) ;
  assign n5394 = ( x79 & n5388 ) | ( x79 & ~n5393 ) | ( n5388 & ~n5393 ) ;
  assign n5395 = ( x79 & n5142 ) | ( x79 & ~n5299 ) | ( n5142 & ~n5299 ) ;
  assign n5396 = x79 & n5142 ;
  assign n5397 = ( ~n5147 & n5395 ) | ( ~n5147 & n5396 ) | ( n5395 & n5396 ) ;
  assign n5398 = ( n5147 & n5395 ) | ( n5147 & n5396 ) | ( n5395 & n5396 ) ;
  assign n5399 = ( n5147 & n5397 ) | ( n5147 & ~n5398 ) | ( n5397 & ~n5398 ) ;
  assign n5400 = ( x80 & n5394 ) | ( x80 & ~n5399 ) | ( n5394 & ~n5399 ) ;
  assign n5401 = ( x80 & n5148 ) | ( x80 & ~n5299 ) | ( n5148 & ~n5299 ) ;
  assign n5402 = x80 & n5148 ;
  assign n5403 = ( ~n5153 & n5401 ) | ( ~n5153 & n5402 ) | ( n5401 & n5402 ) ;
  assign n5404 = ( n5153 & n5401 ) | ( n5153 & n5402 ) | ( n5401 & n5402 ) ;
  assign n5405 = ( n5153 & n5403 ) | ( n5153 & ~n5404 ) | ( n5403 & ~n5404 ) ;
  assign n5406 = ( x81 & n5400 ) | ( x81 & ~n5405 ) | ( n5400 & ~n5405 ) ;
  assign n5407 = ( x81 & n5154 ) | ( x81 & ~n5299 ) | ( n5154 & ~n5299 ) ;
  assign n5408 = x81 & n5154 ;
  assign n5409 = ( ~n5159 & n5407 ) | ( ~n5159 & n5408 ) | ( n5407 & n5408 ) ;
  assign n5410 = ( n5159 & n5407 ) | ( n5159 & n5408 ) | ( n5407 & n5408 ) ;
  assign n5411 = ( n5159 & n5409 ) | ( n5159 & ~n5410 ) | ( n5409 & ~n5410 ) ;
  assign n5412 = ( x82 & n5406 ) | ( x82 & ~n5411 ) | ( n5406 & ~n5411 ) ;
  assign n5413 = ( x82 & n5160 ) | ( x82 & ~n5299 ) | ( n5160 & ~n5299 ) ;
  assign n5414 = x82 & n5160 ;
  assign n5415 = ( ~n5165 & n5413 ) | ( ~n5165 & n5414 ) | ( n5413 & n5414 ) ;
  assign n5416 = ( n5165 & n5413 ) | ( n5165 & n5414 ) | ( n5413 & n5414 ) ;
  assign n5417 = ( n5165 & n5415 ) | ( n5165 & ~n5416 ) | ( n5415 & ~n5416 ) ;
  assign n5418 = ( x83 & n5412 ) | ( x83 & ~n5417 ) | ( n5412 & ~n5417 ) ;
  assign n5419 = ( x83 & n5166 ) | ( x83 & ~n5299 ) | ( n5166 & ~n5299 ) ;
  assign n5420 = x83 & n5166 ;
  assign n5421 = ( ~n5171 & n5419 ) | ( ~n5171 & n5420 ) | ( n5419 & n5420 ) ;
  assign n5422 = ( n5171 & n5419 ) | ( n5171 & n5420 ) | ( n5419 & n5420 ) ;
  assign n5423 = ( n5171 & n5421 ) | ( n5171 & ~n5422 ) | ( n5421 & ~n5422 ) ;
  assign n5424 = ( x84 & n5418 ) | ( x84 & ~n5423 ) | ( n5418 & ~n5423 ) ;
  assign n5425 = ( x84 & n5172 ) | ( x84 & ~n5299 ) | ( n5172 & ~n5299 ) ;
  assign n5426 = x84 & n5172 ;
  assign n5427 = ( ~n5177 & n5425 ) | ( ~n5177 & n5426 ) | ( n5425 & n5426 ) ;
  assign n5428 = ( n5177 & n5425 ) | ( n5177 & n5426 ) | ( n5425 & n5426 ) ;
  assign n5429 = ( n5177 & n5427 ) | ( n5177 & ~n5428 ) | ( n5427 & ~n5428 ) ;
  assign n5430 = ( x85 & n5424 ) | ( x85 & ~n5429 ) | ( n5424 & ~n5429 ) ;
  assign n5431 = ( x85 & n5178 ) | ( x85 & ~n5299 ) | ( n5178 & ~n5299 ) ;
  assign n5432 = x85 & n5178 ;
  assign n5433 = ( ~n5183 & n5431 ) | ( ~n5183 & n5432 ) | ( n5431 & n5432 ) ;
  assign n5434 = ( n5183 & n5431 ) | ( n5183 & n5432 ) | ( n5431 & n5432 ) ;
  assign n5435 = ( n5183 & n5433 ) | ( n5183 & ~n5434 ) | ( n5433 & ~n5434 ) ;
  assign n5436 = ( x86 & n5430 ) | ( x86 & ~n5435 ) | ( n5430 & ~n5435 ) ;
  assign n5437 = ( x86 & n5184 ) | ( x86 & ~n5299 ) | ( n5184 & ~n5299 ) ;
  assign n5438 = x86 & n5184 ;
  assign n5439 = ( ~n5189 & n5437 ) | ( ~n5189 & n5438 ) | ( n5437 & n5438 ) ;
  assign n5440 = ( n5189 & n5437 ) | ( n5189 & n5438 ) | ( n5437 & n5438 ) ;
  assign n5441 = ( n5189 & n5439 ) | ( n5189 & ~n5440 ) | ( n5439 & ~n5440 ) ;
  assign n5442 = ( x87 & n5436 ) | ( x87 & ~n5441 ) | ( n5436 & ~n5441 ) ;
  assign n5443 = ( x87 & n5190 ) | ( x87 & ~n5299 ) | ( n5190 & ~n5299 ) ;
  assign n5444 = x87 & n5190 ;
  assign n5445 = ( ~n5195 & n5443 ) | ( ~n5195 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5446 = ( n5195 & n5443 ) | ( n5195 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5447 = ( n5195 & n5445 ) | ( n5195 & ~n5446 ) | ( n5445 & ~n5446 ) ;
  assign n5448 = ( x88 & n5442 ) | ( x88 & ~n5447 ) | ( n5442 & ~n5447 ) ;
  assign n5449 = ( x88 & n5196 ) | ( x88 & ~n5299 ) | ( n5196 & ~n5299 ) ;
  assign n5450 = x88 & n5196 ;
  assign n5451 = ( ~n5201 & n5449 ) | ( ~n5201 & n5450 ) | ( n5449 & n5450 ) ;
  assign n5452 = ( n5201 & n5449 ) | ( n5201 & n5450 ) | ( n5449 & n5450 ) ;
  assign n5453 = ( n5201 & n5451 ) | ( n5201 & ~n5452 ) | ( n5451 & ~n5452 ) ;
  assign n5454 = ( x89 & n5448 ) | ( x89 & ~n5453 ) | ( n5448 & ~n5453 ) ;
  assign n5455 = ( x89 & n5202 ) | ( x89 & ~n5299 ) | ( n5202 & ~n5299 ) ;
  assign n5456 = x89 & n5202 ;
  assign n5457 = ( ~n5207 & n5455 ) | ( ~n5207 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5458 = ( n5207 & n5455 ) | ( n5207 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5459 = ( n5207 & n5457 ) | ( n5207 & ~n5458 ) | ( n5457 & ~n5458 ) ;
  assign n5460 = ( x90 & n5454 ) | ( x90 & ~n5459 ) | ( n5454 & ~n5459 ) ;
  assign n5461 = ( x90 & n5208 ) | ( x90 & ~n5299 ) | ( n5208 & ~n5299 ) ;
  assign n5462 = x90 & n5208 ;
  assign n5463 = ( ~n5213 & n5461 ) | ( ~n5213 & n5462 ) | ( n5461 & n5462 ) ;
  assign n5464 = ( n5213 & n5461 ) | ( n5213 & n5462 ) | ( n5461 & n5462 ) ;
  assign n5465 = ( n5213 & n5463 ) | ( n5213 & ~n5464 ) | ( n5463 & ~n5464 ) ;
  assign n5466 = ( x91 & n5460 ) | ( x91 & ~n5465 ) | ( n5460 & ~n5465 ) ;
  assign n5467 = ( x91 & n5214 ) | ( x91 & ~n5299 ) | ( n5214 & ~n5299 ) ;
  assign n5468 = x91 & n5214 ;
  assign n5469 = ( ~n5219 & n5467 ) | ( ~n5219 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5470 = ( n5219 & n5467 ) | ( n5219 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5471 = ( n5219 & n5469 ) | ( n5219 & ~n5470 ) | ( n5469 & ~n5470 ) ;
  assign n5472 = ( x92 & n5466 ) | ( x92 & ~n5471 ) | ( n5466 & ~n5471 ) ;
  assign n5473 = ( x92 & n5220 ) | ( x92 & ~n5299 ) | ( n5220 & ~n5299 ) ;
  assign n5474 = x92 & n5220 ;
  assign n5475 = ( ~n5225 & n5473 ) | ( ~n5225 & n5474 ) | ( n5473 & n5474 ) ;
  assign n5476 = ( n5225 & n5473 ) | ( n5225 & n5474 ) | ( n5473 & n5474 ) ;
  assign n5477 = ( n5225 & n5475 ) | ( n5225 & ~n5476 ) | ( n5475 & ~n5476 ) ;
  assign n5478 = ( x93 & n5472 ) | ( x93 & ~n5477 ) | ( n5472 & ~n5477 ) ;
  assign n5479 = ( x93 & n5226 ) | ( x93 & ~n5299 ) | ( n5226 & ~n5299 ) ;
  assign n5480 = x93 & n5226 ;
  assign n5481 = ( ~n5231 & n5479 ) | ( ~n5231 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5482 = ( n5231 & n5479 ) | ( n5231 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5483 = ( n5231 & n5481 ) | ( n5231 & ~n5482 ) | ( n5481 & ~n5482 ) ;
  assign n5484 = ( x94 & n5478 ) | ( x94 & ~n5483 ) | ( n5478 & ~n5483 ) ;
  assign n5485 = ( x94 & n5232 ) | ( x94 & ~n5299 ) | ( n5232 & ~n5299 ) ;
  assign n5486 = x94 & n5232 ;
  assign n5487 = ( ~n5237 & n5485 ) | ( ~n5237 & n5486 ) | ( n5485 & n5486 ) ;
  assign n5488 = ( n5237 & n5485 ) | ( n5237 & n5486 ) | ( n5485 & n5486 ) ;
  assign n5489 = ( n5237 & n5487 ) | ( n5237 & ~n5488 ) | ( n5487 & ~n5488 ) ;
  assign n5490 = ( x95 & n5484 ) | ( x95 & ~n5489 ) | ( n5484 & ~n5489 ) ;
  assign n5491 = ( x95 & n5238 ) | ( x95 & ~n5299 ) | ( n5238 & ~n5299 ) ;
  assign n5492 = x95 & n5238 ;
  assign n5493 = ( ~n5243 & n5491 ) | ( ~n5243 & n5492 ) | ( n5491 & n5492 ) ;
  assign n5494 = ( n5243 & n5491 ) | ( n5243 & n5492 ) | ( n5491 & n5492 ) ;
  assign n5495 = ( n5243 & n5493 ) | ( n5243 & ~n5494 ) | ( n5493 & ~n5494 ) ;
  assign n5496 = ( x96 & n5490 ) | ( x96 & ~n5495 ) | ( n5490 & ~n5495 ) ;
  assign n5497 = ( x96 & n5244 ) | ( x96 & ~n5299 ) | ( n5244 & ~n5299 ) ;
  assign n5498 = x96 & n5244 ;
  assign n5499 = ( ~n5249 & n5497 ) | ( ~n5249 & n5498 ) | ( n5497 & n5498 ) ;
  assign n5500 = ( n5249 & n5497 ) | ( n5249 & n5498 ) | ( n5497 & n5498 ) ;
  assign n5501 = ( n5249 & n5499 ) | ( n5249 & ~n5500 ) | ( n5499 & ~n5500 ) ;
  assign n5502 = ( x97 & n5496 ) | ( x97 & ~n5501 ) | ( n5496 & ~n5501 ) ;
  assign n5503 = ( x97 & n5250 ) | ( x97 & ~n5299 ) | ( n5250 & ~n5299 ) ;
  assign n5504 = x97 & n5250 ;
  assign n5505 = ( ~n5255 & n5503 ) | ( ~n5255 & n5504 ) | ( n5503 & n5504 ) ;
  assign n5506 = ( n5255 & n5503 ) | ( n5255 & n5504 ) | ( n5503 & n5504 ) ;
  assign n5507 = ( n5255 & n5505 ) | ( n5255 & ~n5506 ) | ( n5505 & ~n5506 ) ;
  assign n5508 = ( x98 & n5502 ) | ( x98 & ~n5507 ) | ( n5502 & ~n5507 ) ;
  assign n5509 = ( x98 & n5256 ) | ( x98 & ~n5299 ) | ( n5256 & ~n5299 ) ;
  assign n5510 = x98 & n5256 ;
  assign n5511 = ( ~n5261 & n5509 ) | ( ~n5261 & n5510 ) | ( n5509 & n5510 ) ;
  assign n5512 = ( n5261 & n5509 ) | ( n5261 & n5510 ) | ( n5509 & n5510 ) ;
  assign n5513 = ( n5261 & n5511 ) | ( n5261 & ~n5512 ) | ( n5511 & ~n5512 ) ;
  assign n5514 = ( x99 & n5508 ) | ( x99 & ~n5513 ) | ( n5508 & ~n5513 ) ;
  assign n5515 = ( x99 & n5262 ) | ( x99 & ~n5299 ) | ( n5262 & ~n5299 ) ;
  assign n5516 = x99 & n5262 ;
  assign n5517 = ( ~n5267 & n5515 ) | ( ~n5267 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5518 = ( n5267 & n5515 ) | ( n5267 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5519 = ( n5267 & n5517 ) | ( n5267 & ~n5518 ) | ( n5517 & ~n5518 ) ;
  assign n5520 = ( x100 & n5514 ) | ( x100 & ~n5519 ) | ( n5514 & ~n5519 ) ;
  assign n5521 = ( x100 & n5268 ) | ( x100 & ~n5299 ) | ( n5268 & ~n5299 ) ;
  assign n5522 = x100 & n5268 ;
  assign n5523 = ( ~n5273 & n5521 ) | ( ~n5273 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5524 = ( n5273 & n5521 ) | ( n5273 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5525 = ( n5273 & n5523 ) | ( n5273 & ~n5524 ) | ( n5523 & ~n5524 ) ;
  assign n5526 = ( x101 & n5520 ) | ( x101 & ~n5525 ) | ( n5520 & ~n5525 ) ;
  assign n5527 = ( x101 & n5274 ) | ( x101 & ~n5299 ) | ( n5274 & ~n5299 ) ;
  assign n5528 = x101 & n5274 ;
  assign n5529 = ( ~n5279 & n5527 ) | ( ~n5279 & n5528 ) | ( n5527 & n5528 ) ;
  assign n5530 = ( n5279 & n5527 ) | ( n5279 & n5528 ) | ( n5527 & n5528 ) ;
  assign n5531 = ( n5279 & n5529 ) | ( n5279 & ~n5530 ) | ( n5529 & ~n5530 ) ;
  assign n5532 = ( x102 & n5526 ) | ( x102 & ~n5531 ) | ( n5526 & ~n5531 ) ;
  assign n5533 = ( x102 & n5280 ) | ( x102 & ~n5299 ) | ( n5280 & ~n5299 ) ;
  assign n5534 = x102 & n5280 ;
  assign n5535 = ( ~n5285 & n5533 ) | ( ~n5285 & n5534 ) | ( n5533 & n5534 ) ;
  assign n5536 = ( n5285 & n5533 ) | ( n5285 & n5534 ) | ( n5533 & n5534 ) ;
  assign n5537 = ( n5285 & n5535 ) | ( n5285 & ~n5536 ) | ( n5535 & ~n5536 ) ;
  assign n5538 = ( x103 & n5532 ) | ( x103 & ~n5537 ) | ( n5532 & ~n5537 ) ;
  assign n5539 = ( x103 & n5286 ) | ( x103 & ~n5299 ) | ( n5286 & ~n5299 ) ;
  assign n5540 = x103 & n5286 ;
  assign n5541 = ( ~n5291 & n5539 ) | ( ~n5291 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = ( n5291 & n5539 ) | ( n5291 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5543 = ( n5291 & n5541 ) | ( n5291 & ~n5542 ) | ( n5541 & ~n5542 ) ;
  assign n5544 = ( x104 & n5538 ) | ( x104 & ~n5543 ) | ( n5538 & ~n5543 ) ;
  assign n5545 = ( x105 & ~n5304 ) | ( x105 & n5544 ) | ( ~n5304 & n5544 ) ;
  assign n5546 = n152 & n4814 ;
  assign n5547 = n389 | n5546 ;
  assign n5548 = ( n389 & n5295 ) | ( n389 & n5547 ) | ( n5295 & n5547 ) ;
  assign n5549 = ( x106 & n5545 ) | ( x106 & ~n5548 ) | ( n5545 & ~n5548 ) ;
  assign n5550 = n150 | n5549 ;
  assign n5551 = ( x105 & n5544 ) | ( x105 & n5550 ) | ( n5544 & n5550 ) ;
  assign n5552 = x105 | n5544 ;
  assign n5553 = ( ~n5304 & n5551 ) | ( ~n5304 & n5552 ) | ( n5551 & n5552 ) ;
  assign n5554 = ( n5304 & n5551 ) | ( n5304 & n5552 ) | ( n5551 & n5552 ) ;
  assign n5555 = ( n5304 & n5553 ) | ( n5304 & ~n5554 ) | ( n5553 & ~n5554 ) ;
  assign n5556 = ~x20 & x64 ;
  assign n5557 = ~x21 & n5550 ;
  assign n5558 = ( x21 & ~x64 ) | ( x21 & n5550 ) | ( ~x64 & n5550 ) ;
  assign n5559 = ( n5305 & ~n5557 ) | ( n5305 & n5558 ) | ( ~n5557 & n5558 ) ;
  assign n5560 = ( x65 & n5556 ) | ( x65 & ~n5559 ) | ( n5556 & ~n5559 ) ;
  assign n5561 = ( x65 & n5305 ) | ( x65 & n5550 ) | ( n5305 & n5550 ) ;
  assign n5562 = x65 | n5305 ;
  assign n5563 = ( ~n5309 & n5561 ) | ( ~n5309 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = ( n5309 & n5561 ) | ( n5309 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5565 = ( n5309 & n5563 ) | ( n5309 & ~n5564 ) | ( n5563 & ~n5564 ) ;
  assign n5566 = ( x66 & n5560 ) | ( x66 & ~n5565 ) | ( n5560 & ~n5565 ) ;
  assign n5567 = ( x66 & n5310 ) | ( x66 & n5550 ) | ( n5310 & n5550 ) ;
  assign n5568 = x66 | n5310 ;
  assign n5569 = ( ~n5315 & n5567 ) | ( ~n5315 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5570 = ( n5315 & n5567 ) | ( n5315 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5571 = ( n5315 & n5569 ) | ( n5315 & ~n5570 ) | ( n5569 & ~n5570 ) ;
  assign n5572 = ( x67 & n5566 ) | ( x67 & ~n5571 ) | ( n5566 & ~n5571 ) ;
  assign n5573 = ( x67 & n5316 ) | ( x67 & ~n5550 ) | ( n5316 & ~n5550 ) ;
  assign n5574 = x67 & n5316 ;
  assign n5575 = ( ~n5321 & n5573 ) | ( ~n5321 & n5574 ) | ( n5573 & n5574 ) ;
  assign n5576 = ( n5321 & n5573 ) | ( n5321 & n5574 ) | ( n5573 & n5574 ) ;
  assign n5577 = ( n5321 & n5575 ) | ( n5321 & ~n5576 ) | ( n5575 & ~n5576 ) ;
  assign n5578 = ( x68 & n5572 ) | ( x68 & ~n5577 ) | ( n5572 & ~n5577 ) ;
  assign n5579 = ( x68 & n5322 ) | ( x68 & ~n5550 ) | ( n5322 & ~n5550 ) ;
  assign n5580 = x68 & n5322 ;
  assign n5581 = ( ~n5327 & n5579 ) | ( ~n5327 & n5580 ) | ( n5579 & n5580 ) ;
  assign n5582 = ( n5327 & n5579 ) | ( n5327 & n5580 ) | ( n5579 & n5580 ) ;
  assign n5583 = ( n5327 & n5581 ) | ( n5327 & ~n5582 ) | ( n5581 & ~n5582 ) ;
  assign n5584 = ( x69 & n5578 ) | ( x69 & ~n5583 ) | ( n5578 & ~n5583 ) ;
  assign n5585 = ( x69 & n5328 ) | ( x69 & ~n5550 ) | ( n5328 & ~n5550 ) ;
  assign n5586 = x69 & n5328 ;
  assign n5587 = ( ~n5333 & n5585 ) | ( ~n5333 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5588 = ( n5333 & n5585 ) | ( n5333 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5589 = ( n5333 & n5587 ) | ( n5333 & ~n5588 ) | ( n5587 & ~n5588 ) ;
  assign n5590 = ( x70 & n5584 ) | ( x70 & ~n5589 ) | ( n5584 & ~n5589 ) ;
  assign n5591 = ( x70 & n5334 ) | ( x70 & ~n5550 ) | ( n5334 & ~n5550 ) ;
  assign n5592 = x70 & n5334 ;
  assign n5593 = ( ~n5339 & n5591 ) | ( ~n5339 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5594 = ( n5339 & n5591 ) | ( n5339 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5595 = ( n5339 & n5593 ) | ( n5339 & ~n5594 ) | ( n5593 & ~n5594 ) ;
  assign n5596 = ( x71 & n5590 ) | ( x71 & ~n5595 ) | ( n5590 & ~n5595 ) ;
  assign n5597 = ( x71 & n5340 ) | ( x71 & ~n5550 ) | ( n5340 & ~n5550 ) ;
  assign n5598 = x71 & n5340 ;
  assign n5599 = ( ~n5345 & n5597 ) | ( ~n5345 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5600 = ( n5345 & n5597 ) | ( n5345 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5601 = ( n5345 & n5599 ) | ( n5345 & ~n5600 ) | ( n5599 & ~n5600 ) ;
  assign n5602 = ( x72 & n5596 ) | ( x72 & ~n5601 ) | ( n5596 & ~n5601 ) ;
  assign n5603 = ( x72 & n5346 ) | ( x72 & ~n5550 ) | ( n5346 & ~n5550 ) ;
  assign n5604 = x72 & n5346 ;
  assign n5605 = ( ~n5351 & n5603 ) | ( ~n5351 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5606 = ( n5351 & n5603 ) | ( n5351 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5607 = ( n5351 & n5605 ) | ( n5351 & ~n5606 ) | ( n5605 & ~n5606 ) ;
  assign n5608 = ( x73 & n5602 ) | ( x73 & ~n5607 ) | ( n5602 & ~n5607 ) ;
  assign n5609 = ( x73 & n5352 ) | ( x73 & ~n5550 ) | ( n5352 & ~n5550 ) ;
  assign n5610 = x73 & n5352 ;
  assign n5611 = ( ~n5357 & n5609 ) | ( ~n5357 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5612 = ( n5357 & n5609 ) | ( n5357 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5613 = ( n5357 & n5611 ) | ( n5357 & ~n5612 ) | ( n5611 & ~n5612 ) ;
  assign n5614 = ( x74 & n5608 ) | ( x74 & ~n5613 ) | ( n5608 & ~n5613 ) ;
  assign n5615 = ( x74 & n5358 ) | ( x74 & ~n5550 ) | ( n5358 & ~n5550 ) ;
  assign n5616 = x74 & n5358 ;
  assign n5617 = ( ~n5363 & n5615 ) | ( ~n5363 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5618 = ( n5363 & n5615 ) | ( n5363 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5619 = ( n5363 & n5617 ) | ( n5363 & ~n5618 ) | ( n5617 & ~n5618 ) ;
  assign n5620 = ( x75 & n5614 ) | ( x75 & ~n5619 ) | ( n5614 & ~n5619 ) ;
  assign n5621 = ( x75 & n5364 ) | ( x75 & ~n5550 ) | ( n5364 & ~n5550 ) ;
  assign n5622 = x75 & n5364 ;
  assign n5623 = ( ~n5369 & n5621 ) | ( ~n5369 & n5622 ) | ( n5621 & n5622 ) ;
  assign n5624 = ( n5369 & n5621 ) | ( n5369 & n5622 ) | ( n5621 & n5622 ) ;
  assign n5625 = ( n5369 & n5623 ) | ( n5369 & ~n5624 ) | ( n5623 & ~n5624 ) ;
  assign n5626 = ( x76 & n5620 ) | ( x76 & ~n5625 ) | ( n5620 & ~n5625 ) ;
  assign n5627 = ( x76 & n5370 ) | ( x76 & ~n5550 ) | ( n5370 & ~n5550 ) ;
  assign n5628 = x76 & n5370 ;
  assign n5629 = ( ~n5375 & n5627 ) | ( ~n5375 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5630 = ( n5375 & n5627 ) | ( n5375 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5631 = ( n5375 & n5629 ) | ( n5375 & ~n5630 ) | ( n5629 & ~n5630 ) ;
  assign n5632 = ( x77 & n5626 ) | ( x77 & ~n5631 ) | ( n5626 & ~n5631 ) ;
  assign n5633 = ( x77 & n5376 ) | ( x77 & ~n5550 ) | ( n5376 & ~n5550 ) ;
  assign n5634 = x77 & n5376 ;
  assign n5635 = ( ~n5381 & n5633 ) | ( ~n5381 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5636 = ( n5381 & n5633 ) | ( n5381 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5637 = ( n5381 & n5635 ) | ( n5381 & ~n5636 ) | ( n5635 & ~n5636 ) ;
  assign n5638 = ( x78 & n5632 ) | ( x78 & ~n5637 ) | ( n5632 & ~n5637 ) ;
  assign n5639 = ( x78 & n5382 ) | ( x78 & ~n5550 ) | ( n5382 & ~n5550 ) ;
  assign n5640 = x78 & n5382 ;
  assign n5641 = ( ~n5387 & n5639 ) | ( ~n5387 & n5640 ) | ( n5639 & n5640 ) ;
  assign n5642 = ( n5387 & n5639 ) | ( n5387 & n5640 ) | ( n5639 & n5640 ) ;
  assign n5643 = ( n5387 & n5641 ) | ( n5387 & ~n5642 ) | ( n5641 & ~n5642 ) ;
  assign n5644 = ( x79 & n5638 ) | ( x79 & ~n5643 ) | ( n5638 & ~n5643 ) ;
  assign n5645 = ( x79 & n5388 ) | ( x79 & ~n5550 ) | ( n5388 & ~n5550 ) ;
  assign n5646 = x79 & n5388 ;
  assign n5647 = ( ~n5393 & n5645 ) | ( ~n5393 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5648 = ( n5393 & n5645 ) | ( n5393 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5649 = ( n5393 & n5647 ) | ( n5393 & ~n5648 ) | ( n5647 & ~n5648 ) ;
  assign n5650 = ( x80 & n5644 ) | ( x80 & ~n5649 ) | ( n5644 & ~n5649 ) ;
  assign n5651 = ( x80 & n5394 ) | ( x80 & ~n5550 ) | ( n5394 & ~n5550 ) ;
  assign n5652 = x80 & n5394 ;
  assign n5653 = ( ~n5399 & n5651 ) | ( ~n5399 & n5652 ) | ( n5651 & n5652 ) ;
  assign n5654 = ( n5399 & n5651 ) | ( n5399 & n5652 ) | ( n5651 & n5652 ) ;
  assign n5655 = ( n5399 & n5653 ) | ( n5399 & ~n5654 ) | ( n5653 & ~n5654 ) ;
  assign n5656 = ( x81 & n5650 ) | ( x81 & ~n5655 ) | ( n5650 & ~n5655 ) ;
  assign n5657 = ( x81 & n5400 ) | ( x81 & ~n5550 ) | ( n5400 & ~n5550 ) ;
  assign n5658 = x81 & n5400 ;
  assign n5659 = ( ~n5405 & n5657 ) | ( ~n5405 & n5658 ) | ( n5657 & n5658 ) ;
  assign n5660 = ( n5405 & n5657 ) | ( n5405 & n5658 ) | ( n5657 & n5658 ) ;
  assign n5661 = ( n5405 & n5659 ) | ( n5405 & ~n5660 ) | ( n5659 & ~n5660 ) ;
  assign n5662 = ( x82 & n5656 ) | ( x82 & ~n5661 ) | ( n5656 & ~n5661 ) ;
  assign n5663 = ( x82 & n5406 ) | ( x82 & ~n5550 ) | ( n5406 & ~n5550 ) ;
  assign n5664 = x82 & n5406 ;
  assign n5665 = ( ~n5411 & n5663 ) | ( ~n5411 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5666 = ( n5411 & n5663 ) | ( n5411 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5667 = ( n5411 & n5665 ) | ( n5411 & ~n5666 ) | ( n5665 & ~n5666 ) ;
  assign n5668 = ( x83 & n5662 ) | ( x83 & ~n5667 ) | ( n5662 & ~n5667 ) ;
  assign n5669 = ( x83 & n5412 ) | ( x83 & ~n5550 ) | ( n5412 & ~n5550 ) ;
  assign n5670 = x83 & n5412 ;
  assign n5671 = ( ~n5417 & n5669 ) | ( ~n5417 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = ( n5417 & n5669 ) | ( n5417 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5673 = ( n5417 & n5671 ) | ( n5417 & ~n5672 ) | ( n5671 & ~n5672 ) ;
  assign n5674 = ( x84 & n5668 ) | ( x84 & ~n5673 ) | ( n5668 & ~n5673 ) ;
  assign n5675 = ( x84 & n5418 ) | ( x84 & ~n5550 ) | ( n5418 & ~n5550 ) ;
  assign n5676 = x84 & n5418 ;
  assign n5677 = ( ~n5423 & n5675 ) | ( ~n5423 & n5676 ) | ( n5675 & n5676 ) ;
  assign n5678 = ( n5423 & n5675 ) | ( n5423 & n5676 ) | ( n5675 & n5676 ) ;
  assign n5679 = ( n5423 & n5677 ) | ( n5423 & ~n5678 ) | ( n5677 & ~n5678 ) ;
  assign n5680 = ( x85 & n5674 ) | ( x85 & ~n5679 ) | ( n5674 & ~n5679 ) ;
  assign n5681 = ( x85 & n5424 ) | ( x85 & ~n5550 ) | ( n5424 & ~n5550 ) ;
  assign n5682 = x85 & n5424 ;
  assign n5683 = ( ~n5429 & n5681 ) | ( ~n5429 & n5682 ) | ( n5681 & n5682 ) ;
  assign n5684 = ( n5429 & n5681 ) | ( n5429 & n5682 ) | ( n5681 & n5682 ) ;
  assign n5685 = ( n5429 & n5683 ) | ( n5429 & ~n5684 ) | ( n5683 & ~n5684 ) ;
  assign n5686 = ( x86 & n5680 ) | ( x86 & ~n5685 ) | ( n5680 & ~n5685 ) ;
  assign n5687 = ( x86 & n5430 ) | ( x86 & ~n5550 ) | ( n5430 & ~n5550 ) ;
  assign n5688 = x86 & n5430 ;
  assign n5689 = ( ~n5435 & n5687 ) | ( ~n5435 & n5688 ) | ( n5687 & n5688 ) ;
  assign n5690 = ( n5435 & n5687 ) | ( n5435 & n5688 ) | ( n5687 & n5688 ) ;
  assign n5691 = ( n5435 & n5689 ) | ( n5435 & ~n5690 ) | ( n5689 & ~n5690 ) ;
  assign n5692 = ( x87 & n5686 ) | ( x87 & ~n5691 ) | ( n5686 & ~n5691 ) ;
  assign n5693 = ( x87 & n5436 ) | ( x87 & ~n5550 ) | ( n5436 & ~n5550 ) ;
  assign n5694 = x87 & n5436 ;
  assign n5695 = ( ~n5441 & n5693 ) | ( ~n5441 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5696 = ( n5441 & n5693 ) | ( n5441 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5697 = ( n5441 & n5695 ) | ( n5441 & ~n5696 ) | ( n5695 & ~n5696 ) ;
  assign n5698 = ( x88 & n5692 ) | ( x88 & ~n5697 ) | ( n5692 & ~n5697 ) ;
  assign n5699 = ( x88 & n5442 ) | ( x88 & ~n5550 ) | ( n5442 & ~n5550 ) ;
  assign n5700 = x88 & n5442 ;
  assign n5701 = ( ~n5447 & n5699 ) | ( ~n5447 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5702 = ( n5447 & n5699 ) | ( n5447 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5703 = ( n5447 & n5701 ) | ( n5447 & ~n5702 ) | ( n5701 & ~n5702 ) ;
  assign n5704 = ( x89 & n5698 ) | ( x89 & ~n5703 ) | ( n5698 & ~n5703 ) ;
  assign n5705 = ( x89 & n5448 ) | ( x89 & ~n5550 ) | ( n5448 & ~n5550 ) ;
  assign n5706 = x89 & n5448 ;
  assign n5707 = ( ~n5453 & n5705 ) | ( ~n5453 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = ( n5453 & n5705 ) | ( n5453 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5709 = ( n5453 & n5707 ) | ( n5453 & ~n5708 ) | ( n5707 & ~n5708 ) ;
  assign n5710 = ( x90 & n5704 ) | ( x90 & ~n5709 ) | ( n5704 & ~n5709 ) ;
  assign n5711 = ( x90 & n5454 ) | ( x90 & ~n5550 ) | ( n5454 & ~n5550 ) ;
  assign n5712 = x90 & n5454 ;
  assign n5713 = ( ~n5459 & n5711 ) | ( ~n5459 & n5712 ) | ( n5711 & n5712 ) ;
  assign n5714 = ( n5459 & n5711 ) | ( n5459 & n5712 ) | ( n5711 & n5712 ) ;
  assign n5715 = ( n5459 & n5713 ) | ( n5459 & ~n5714 ) | ( n5713 & ~n5714 ) ;
  assign n5716 = ( x91 & n5710 ) | ( x91 & ~n5715 ) | ( n5710 & ~n5715 ) ;
  assign n5717 = ( x91 & n5460 ) | ( x91 & ~n5550 ) | ( n5460 & ~n5550 ) ;
  assign n5718 = x91 & n5460 ;
  assign n5719 = ( ~n5465 & n5717 ) | ( ~n5465 & n5718 ) | ( n5717 & n5718 ) ;
  assign n5720 = ( n5465 & n5717 ) | ( n5465 & n5718 ) | ( n5717 & n5718 ) ;
  assign n5721 = ( n5465 & n5719 ) | ( n5465 & ~n5720 ) | ( n5719 & ~n5720 ) ;
  assign n5722 = ( x92 & n5716 ) | ( x92 & ~n5721 ) | ( n5716 & ~n5721 ) ;
  assign n5723 = ( x92 & n5466 ) | ( x92 & ~n5550 ) | ( n5466 & ~n5550 ) ;
  assign n5724 = x92 & n5466 ;
  assign n5725 = ( ~n5471 & n5723 ) | ( ~n5471 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5726 = ( n5471 & n5723 ) | ( n5471 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5727 = ( n5471 & n5725 ) | ( n5471 & ~n5726 ) | ( n5725 & ~n5726 ) ;
  assign n5728 = ( x93 & n5722 ) | ( x93 & ~n5727 ) | ( n5722 & ~n5727 ) ;
  assign n5729 = ( x93 & n5472 ) | ( x93 & ~n5550 ) | ( n5472 & ~n5550 ) ;
  assign n5730 = x93 & n5472 ;
  assign n5731 = ( ~n5477 & n5729 ) | ( ~n5477 & n5730 ) | ( n5729 & n5730 ) ;
  assign n5732 = ( n5477 & n5729 ) | ( n5477 & n5730 ) | ( n5729 & n5730 ) ;
  assign n5733 = ( n5477 & n5731 ) | ( n5477 & ~n5732 ) | ( n5731 & ~n5732 ) ;
  assign n5734 = ( x94 & n5728 ) | ( x94 & ~n5733 ) | ( n5728 & ~n5733 ) ;
  assign n5735 = ( x94 & n5478 ) | ( x94 & ~n5550 ) | ( n5478 & ~n5550 ) ;
  assign n5736 = x94 & n5478 ;
  assign n5737 = ( ~n5483 & n5735 ) | ( ~n5483 & n5736 ) | ( n5735 & n5736 ) ;
  assign n5738 = ( n5483 & n5735 ) | ( n5483 & n5736 ) | ( n5735 & n5736 ) ;
  assign n5739 = ( n5483 & n5737 ) | ( n5483 & ~n5738 ) | ( n5737 & ~n5738 ) ;
  assign n5740 = ( x95 & n5734 ) | ( x95 & ~n5739 ) | ( n5734 & ~n5739 ) ;
  assign n5741 = ( x95 & n5484 ) | ( x95 & ~n5550 ) | ( n5484 & ~n5550 ) ;
  assign n5742 = x95 & n5484 ;
  assign n5743 = ( ~n5489 & n5741 ) | ( ~n5489 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5744 = ( n5489 & n5741 ) | ( n5489 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5745 = ( n5489 & n5743 ) | ( n5489 & ~n5744 ) | ( n5743 & ~n5744 ) ;
  assign n5746 = ( x96 & n5740 ) | ( x96 & ~n5745 ) | ( n5740 & ~n5745 ) ;
  assign n5747 = ( x96 & n5490 ) | ( x96 & ~n5550 ) | ( n5490 & ~n5550 ) ;
  assign n5748 = x96 & n5490 ;
  assign n5749 = ( ~n5495 & n5747 ) | ( ~n5495 & n5748 ) | ( n5747 & n5748 ) ;
  assign n5750 = ( n5495 & n5747 ) | ( n5495 & n5748 ) | ( n5747 & n5748 ) ;
  assign n5751 = ( n5495 & n5749 ) | ( n5495 & ~n5750 ) | ( n5749 & ~n5750 ) ;
  assign n5752 = ( x97 & n5746 ) | ( x97 & ~n5751 ) | ( n5746 & ~n5751 ) ;
  assign n5753 = ( x97 & n5496 ) | ( x97 & ~n5550 ) | ( n5496 & ~n5550 ) ;
  assign n5754 = x97 & n5496 ;
  assign n5755 = ( ~n5501 & n5753 ) | ( ~n5501 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5756 = ( n5501 & n5753 ) | ( n5501 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5757 = ( n5501 & n5755 ) | ( n5501 & ~n5756 ) | ( n5755 & ~n5756 ) ;
  assign n5758 = ( x98 & n5752 ) | ( x98 & ~n5757 ) | ( n5752 & ~n5757 ) ;
  assign n5759 = ( x98 & n5502 ) | ( x98 & ~n5550 ) | ( n5502 & ~n5550 ) ;
  assign n5760 = x98 & n5502 ;
  assign n5761 = ( ~n5507 & n5759 ) | ( ~n5507 & n5760 ) | ( n5759 & n5760 ) ;
  assign n5762 = ( n5507 & n5759 ) | ( n5507 & n5760 ) | ( n5759 & n5760 ) ;
  assign n5763 = ( n5507 & n5761 ) | ( n5507 & ~n5762 ) | ( n5761 & ~n5762 ) ;
  assign n5764 = ( x99 & n5758 ) | ( x99 & ~n5763 ) | ( n5758 & ~n5763 ) ;
  assign n5765 = ( x99 & n5508 ) | ( x99 & ~n5550 ) | ( n5508 & ~n5550 ) ;
  assign n5766 = x99 & n5508 ;
  assign n5767 = ( ~n5513 & n5765 ) | ( ~n5513 & n5766 ) | ( n5765 & n5766 ) ;
  assign n5768 = ( n5513 & n5765 ) | ( n5513 & n5766 ) | ( n5765 & n5766 ) ;
  assign n5769 = ( n5513 & n5767 ) | ( n5513 & ~n5768 ) | ( n5767 & ~n5768 ) ;
  assign n5770 = ( x100 & n5764 ) | ( x100 & ~n5769 ) | ( n5764 & ~n5769 ) ;
  assign n5771 = ( x100 & n5514 ) | ( x100 & ~n5550 ) | ( n5514 & ~n5550 ) ;
  assign n5772 = x100 & n5514 ;
  assign n5773 = ( ~n5519 & n5771 ) | ( ~n5519 & n5772 ) | ( n5771 & n5772 ) ;
  assign n5774 = ( n5519 & n5771 ) | ( n5519 & n5772 ) | ( n5771 & n5772 ) ;
  assign n5775 = ( n5519 & n5773 ) | ( n5519 & ~n5774 ) | ( n5773 & ~n5774 ) ;
  assign n5776 = ( x101 & n5770 ) | ( x101 & ~n5775 ) | ( n5770 & ~n5775 ) ;
  assign n5777 = ( x101 & n5520 ) | ( x101 & ~n5550 ) | ( n5520 & ~n5550 ) ;
  assign n5778 = x101 & n5520 ;
  assign n5779 = ( ~n5525 & n5777 ) | ( ~n5525 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = ( n5525 & n5777 ) | ( n5525 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5781 = ( n5525 & n5779 ) | ( n5525 & ~n5780 ) | ( n5779 & ~n5780 ) ;
  assign n5782 = ( x102 & n5776 ) | ( x102 & ~n5781 ) | ( n5776 & ~n5781 ) ;
  assign n5783 = ( x102 & n5526 ) | ( x102 & ~n5550 ) | ( n5526 & ~n5550 ) ;
  assign n5784 = x102 & n5526 ;
  assign n5785 = ( ~n5531 & n5783 ) | ( ~n5531 & n5784 ) | ( n5783 & n5784 ) ;
  assign n5786 = ( n5531 & n5783 ) | ( n5531 & n5784 ) | ( n5783 & n5784 ) ;
  assign n5787 = ( n5531 & n5785 ) | ( n5531 & ~n5786 ) | ( n5785 & ~n5786 ) ;
  assign n5788 = ( x103 & n5782 ) | ( x103 & ~n5787 ) | ( n5782 & ~n5787 ) ;
  assign n5789 = ( x103 & n5532 ) | ( x103 & ~n5550 ) | ( n5532 & ~n5550 ) ;
  assign n5790 = x103 & n5532 ;
  assign n5791 = ( ~n5537 & n5789 ) | ( ~n5537 & n5790 ) | ( n5789 & n5790 ) ;
  assign n5792 = ( n5537 & n5789 ) | ( n5537 & n5790 ) | ( n5789 & n5790 ) ;
  assign n5793 = ( n5537 & n5791 ) | ( n5537 & ~n5792 ) | ( n5791 & ~n5792 ) ;
  assign n5794 = ( x104 & n5788 ) | ( x104 & ~n5793 ) | ( n5788 & ~n5793 ) ;
  assign n5795 = ( x104 & n5538 ) | ( x104 & ~n5550 ) | ( n5538 & ~n5550 ) ;
  assign n5796 = x104 & n5538 ;
  assign n5797 = ( ~n5543 & n5795 ) | ( ~n5543 & n5796 ) | ( n5795 & n5796 ) ;
  assign n5798 = ( n5543 & n5795 ) | ( n5543 & n5796 ) | ( n5795 & n5796 ) ;
  assign n5799 = ( n5543 & n5797 ) | ( n5543 & ~n5798 ) | ( n5797 & ~n5798 ) ;
  assign n5800 = ( x105 & n5794 ) | ( x105 & ~n5799 ) | ( n5794 & ~n5799 ) ;
  assign n5801 = ( x106 & ~n5555 ) | ( x106 & n5800 ) | ( ~n5555 & n5800 ) ;
  assign n5802 = ( x106 & n150 ) | ( x106 & n5545 ) | ( n150 & n5545 ) ;
  assign n5803 = x106 | n5545 ;
  assign n5804 = ( n5548 & n5802 ) | ( n5548 & ~n5803 ) | ( n5802 & ~n5803 ) ;
  assign n5805 = ( x107 & n5801 ) | ( x107 & ~n5804 ) | ( n5801 & ~n5804 ) ;
  assign n5806 = n149 | n5805 ;
  assign n5807 = ( x106 & n5800 ) | ( x106 & n5806 ) | ( n5800 & n5806 ) ;
  assign n5808 = x106 | n5800 ;
  assign n5809 = ( ~n5555 & n5807 ) | ( ~n5555 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5810 = ( n5555 & n5807 ) | ( n5555 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5811 = ( n5555 & n5809 ) | ( n5555 & ~n5810 ) | ( n5809 & ~n5810 ) ;
  assign n5812 = ~x19 & x64 ;
  assign n5813 = ~x20 & n5806 ;
  assign n5814 = ( x20 & ~x64 ) | ( x20 & n5806 ) | ( ~x64 & n5806 ) ;
  assign n5815 = ( n5556 & ~n5813 ) | ( n5556 & n5814 ) | ( ~n5813 & n5814 ) ;
  assign n5816 = ( x65 & n5812 ) | ( x65 & ~n5815 ) | ( n5812 & ~n5815 ) ;
  assign n5817 = ( x65 & n5556 ) | ( x65 & n5806 ) | ( n5556 & n5806 ) ;
  assign n5818 = x65 | n5556 ;
  assign n5819 = ( ~n5559 & n5817 ) | ( ~n5559 & n5818 ) | ( n5817 & n5818 ) ;
  assign n5820 = ( n5559 & n5817 ) | ( n5559 & n5818 ) | ( n5817 & n5818 ) ;
  assign n5821 = ( n5559 & n5819 ) | ( n5559 & ~n5820 ) | ( n5819 & ~n5820 ) ;
  assign n5822 = ( x66 & n5816 ) | ( x66 & ~n5821 ) | ( n5816 & ~n5821 ) ;
  assign n5823 = ( x66 & n5560 ) | ( x66 & n5806 ) | ( n5560 & n5806 ) ;
  assign n5824 = x66 | n5560 ;
  assign n5825 = ( ~n5565 & n5823 ) | ( ~n5565 & n5824 ) | ( n5823 & n5824 ) ;
  assign n5826 = ( n5565 & n5823 ) | ( n5565 & n5824 ) | ( n5823 & n5824 ) ;
  assign n5827 = ( n5565 & n5825 ) | ( n5565 & ~n5826 ) | ( n5825 & ~n5826 ) ;
  assign n5828 = ( x67 & n5822 ) | ( x67 & ~n5827 ) | ( n5822 & ~n5827 ) ;
  assign n5829 = ( x67 & n5566 ) | ( x67 & ~n5806 ) | ( n5566 & ~n5806 ) ;
  assign n5830 = x67 & n5566 ;
  assign n5831 = ( ~n5571 & n5829 ) | ( ~n5571 & n5830 ) | ( n5829 & n5830 ) ;
  assign n5832 = ( n5571 & n5829 ) | ( n5571 & n5830 ) | ( n5829 & n5830 ) ;
  assign n5833 = ( n5571 & n5831 ) | ( n5571 & ~n5832 ) | ( n5831 & ~n5832 ) ;
  assign n5834 = ( x68 & n5828 ) | ( x68 & ~n5833 ) | ( n5828 & ~n5833 ) ;
  assign n5835 = ( x68 & n5572 ) | ( x68 & ~n5806 ) | ( n5572 & ~n5806 ) ;
  assign n5836 = x68 & n5572 ;
  assign n5837 = ( ~n5577 & n5835 ) | ( ~n5577 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = ( n5577 & n5835 ) | ( n5577 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5839 = ( n5577 & n5837 ) | ( n5577 & ~n5838 ) | ( n5837 & ~n5838 ) ;
  assign n5840 = ( x69 & n5834 ) | ( x69 & ~n5839 ) | ( n5834 & ~n5839 ) ;
  assign n5841 = ( x69 & n5578 ) | ( x69 & ~n5806 ) | ( n5578 & ~n5806 ) ;
  assign n5842 = x69 & n5578 ;
  assign n5843 = ( ~n5583 & n5841 ) | ( ~n5583 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = ( n5583 & n5841 ) | ( n5583 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5845 = ( n5583 & n5843 ) | ( n5583 & ~n5844 ) | ( n5843 & ~n5844 ) ;
  assign n5846 = ( x70 & n5840 ) | ( x70 & ~n5845 ) | ( n5840 & ~n5845 ) ;
  assign n5847 = ( x70 & n5584 ) | ( x70 & ~n5806 ) | ( n5584 & ~n5806 ) ;
  assign n5848 = x70 & n5584 ;
  assign n5849 = ( ~n5589 & n5847 ) | ( ~n5589 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5850 = ( n5589 & n5847 ) | ( n5589 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5851 = ( n5589 & n5849 ) | ( n5589 & ~n5850 ) | ( n5849 & ~n5850 ) ;
  assign n5852 = ( x71 & n5846 ) | ( x71 & ~n5851 ) | ( n5846 & ~n5851 ) ;
  assign n5853 = ( x71 & n5590 ) | ( x71 & ~n5806 ) | ( n5590 & ~n5806 ) ;
  assign n5854 = x71 & n5590 ;
  assign n5855 = ( ~n5595 & n5853 ) | ( ~n5595 & n5854 ) | ( n5853 & n5854 ) ;
  assign n5856 = ( n5595 & n5853 ) | ( n5595 & n5854 ) | ( n5853 & n5854 ) ;
  assign n5857 = ( n5595 & n5855 ) | ( n5595 & ~n5856 ) | ( n5855 & ~n5856 ) ;
  assign n5858 = ( x72 & n5852 ) | ( x72 & ~n5857 ) | ( n5852 & ~n5857 ) ;
  assign n5859 = ( x72 & n5596 ) | ( x72 & ~n5806 ) | ( n5596 & ~n5806 ) ;
  assign n5860 = x72 & n5596 ;
  assign n5861 = ( ~n5601 & n5859 ) | ( ~n5601 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5862 = ( n5601 & n5859 ) | ( n5601 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5863 = ( n5601 & n5861 ) | ( n5601 & ~n5862 ) | ( n5861 & ~n5862 ) ;
  assign n5864 = ( x73 & n5858 ) | ( x73 & ~n5863 ) | ( n5858 & ~n5863 ) ;
  assign n5865 = ( x73 & n5602 ) | ( x73 & ~n5806 ) | ( n5602 & ~n5806 ) ;
  assign n5866 = x73 & n5602 ;
  assign n5867 = ( ~n5607 & n5865 ) | ( ~n5607 & n5866 ) | ( n5865 & n5866 ) ;
  assign n5868 = ( n5607 & n5865 ) | ( n5607 & n5866 ) | ( n5865 & n5866 ) ;
  assign n5869 = ( n5607 & n5867 ) | ( n5607 & ~n5868 ) | ( n5867 & ~n5868 ) ;
  assign n5870 = ( x74 & n5864 ) | ( x74 & ~n5869 ) | ( n5864 & ~n5869 ) ;
  assign n5871 = ( x74 & n5608 ) | ( x74 & ~n5806 ) | ( n5608 & ~n5806 ) ;
  assign n5872 = x74 & n5608 ;
  assign n5873 = ( ~n5613 & n5871 ) | ( ~n5613 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5874 = ( n5613 & n5871 ) | ( n5613 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5875 = ( n5613 & n5873 ) | ( n5613 & ~n5874 ) | ( n5873 & ~n5874 ) ;
  assign n5876 = ( x75 & n5870 ) | ( x75 & ~n5875 ) | ( n5870 & ~n5875 ) ;
  assign n5877 = ( x75 & n5614 ) | ( x75 & ~n5806 ) | ( n5614 & ~n5806 ) ;
  assign n5878 = x75 & n5614 ;
  assign n5879 = ( ~n5619 & n5877 ) | ( ~n5619 & n5878 ) | ( n5877 & n5878 ) ;
  assign n5880 = ( n5619 & n5877 ) | ( n5619 & n5878 ) | ( n5877 & n5878 ) ;
  assign n5881 = ( n5619 & n5879 ) | ( n5619 & ~n5880 ) | ( n5879 & ~n5880 ) ;
  assign n5882 = ( x76 & n5876 ) | ( x76 & ~n5881 ) | ( n5876 & ~n5881 ) ;
  assign n5883 = ( x76 & n5620 ) | ( x76 & ~n5806 ) | ( n5620 & ~n5806 ) ;
  assign n5884 = x76 & n5620 ;
  assign n5885 = ( ~n5625 & n5883 ) | ( ~n5625 & n5884 ) | ( n5883 & n5884 ) ;
  assign n5886 = ( n5625 & n5883 ) | ( n5625 & n5884 ) | ( n5883 & n5884 ) ;
  assign n5887 = ( n5625 & n5885 ) | ( n5625 & ~n5886 ) | ( n5885 & ~n5886 ) ;
  assign n5888 = ( x77 & n5882 ) | ( x77 & ~n5887 ) | ( n5882 & ~n5887 ) ;
  assign n5889 = ( x77 & n5626 ) | ( x77 & ~n5806 ) | ( n5626 & ~n5806 ) ;
  assign n5890 = x77 & n5626 ;
  assign n5891 = ( ~n5631 & n5889 ) | ( ~n5631 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5892 = ( n5631 & n5889 ) | ( n5631 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5893 = ( n5631 & n5891 ) | ( n5631 & ~n5892 ) | ( n5891 & ~n5892 ) ;
  assign n5894 = ( x78 & n5888 ) | ( x78 & ~n5893 ) | ( n5888 & ~n5893 ) ;
  assign n5895 = ( x78 & n5632 ) | ( x78 & ~n5806 ) | ( n5632 & ~n5806 ) ;
  assign n5896 = x78 & n5632 ;
  assign n5897 = ( ~n5637 & n5895 ) | ( ~n5637 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5898 = ( n5637 & n5895 ) | ( n5637 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5899 = ( n5637 & n5897 ) | ( n5637 & ~n5898 ) | ( n5897 & ~n5898 ) ;
  assign n5900 = ( x79 & n5894 ) | ( x79 & ~n5899 ) | ( n5894 & ~n5899 ) ;
  assign n5901 = ( x79 & n5638 ) | ( x79 & ~n5806 ) | ( n5638 & ~n5806 ) ;
  assign n5902 = x79 & n5638 ;
  assign n5903 = ( ~n5643 & n5901 ) | ( ~n5643 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5904 = ( n5643 & n5901 ) | ( n5643 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5905 = ( n5643 & n5903 ) | ( n5643 & ~n5904 ) | ( n5903 & ~n5904 ) ;
  assign n5906 = ( x80 & n5900 ) | ( x80 & ~n5905 ) | ( n5900 & ~n5905 ) ;
  assign n5907 = ( x80 & n5644 ) | ( x80 & ~n5806 ) | ( n5644 & ~n5806 ) ;
  assign n5908 = x80 & n5644 ;
  assign n5909 = ( ~n5649 & n5907 ) | ( ~n5649 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5910 = ( n5649 & n5907 ) | ( n5649 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5911 = ( n5649 & n5909 ) | ( n5649 & ~n5910 ) | ( n5909 & ~n5910 ) ;
  assign n5912 = ( x81 & n5906 ) | ( x81 & ~n5911 ) | ( n5906 & ~n5911 ) ;
  assign n5913 = ( x81 & n5650 ) | ( x81 & ~n5806 ) | ( n5650 & ~n5806 ) ;
  assign n5914 = x81 & n5650 ;
  assign n5915 = ( ~n5655 & n5913 ) | ( ~n5655 & n5914 ) | ( n5913 & n5914 ) ;
  assign n5916 = ( n5655 & n5913 ) | ( n5655 & n5914 ) | ( n5913 & n5914 ) ;
  assign n5917 = ( n5655 & n5915 ) | ( n5655 & ~n5916 ) | ( n5915 & ~n5916 ) ;
  assign n5918 = ( x82 & n5912 ) | ( x82 & ~n5917 ) | ( n5912 & ~n5917 ) ;
  assign n5919 = ( x82 & n5656 ) | ( x82 & ~n5806 ) | ( n5656 & ~n5806 ) ;
  assign n5920 = x82 & n5656 ;
  assign n5921 = ( ~n5661 & n5919 ) | ( ~n5661 & n5920 ) | ( n5919 & n5920 ) ;
  assign n5922 = ( n5661 & n5919 ) | ( n5661 & n5920 ) | ( n5919 & n5920 ) ;
  assign n5923 = ( n5661 & n5921 ) | ( n5661 & ~n5922 ) | ( n5921 & ~n5922 ) ;
  assign n5924 = ( x83 & n5918 ) | ( x83 & ~n5923 ) | ( n5918 & ~n5923 ) ;
  assign n5925 = ( x83 & n5662 ) | ( x83 & ~n5806 ) | ( n5662 & ~n5806 ) ;
  assign n5926 = x83 & n5662 ;
  assign n5927 = ( ~n5667 & n5925 ) | ( ~n5667 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5928 = ( n5667 & n5925 ) | ( n5667 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5929 = ( n5667 & n5927 ) | ( n5667 & ~n5928 ) | ( n5927 & ~n5928 ) ;
  assign n5930 = ( x84 & n5924 ) | ( x84 & ~n5929 ) | ( n5924 & ~n5929 ) ;
  assign n5931 = ( x84 & n5668 ) | ( x84 & ~n5806 ) | ( n5668 & ~n5806 ) ;
  assign n5932 = x84 & n5668 ;
  assign n5933 = ( ~n5673 & n5931 ) | ( ~n5673 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5934 = ( n5673 & n5931 ) | ( n5673 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5935 = ( n5673 & n5933 ) | ( n5673 & ~n5934 ) | ( n5933 & ~n5934 ) ;
  assign n5936 = ( x85 & n5930 ) | ( x85 & ~n5935 ) | ( n5930 & ~n5935 ) ;
  assign n5937 = ( x85 & n5674 ) | ( x85 & ~n5806 ) | ( n5674 & ~n5806 ) ;
  assign n5938 = x85 & n5674 ;
  assign n5939 = ( ~n5679 & n5937 ) | ( ~n5679 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5940 = ( n5679 & n5937 ) | ( n5679 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5941 = ( n5679 & n5939 ) | ( n5679 & ~n5940 ) | ( n5939 & ~n5940 ) ;
  assign n5942 = ( x86 & n5936 ) | ( x86 & ~n5941 ) | ( n5936 & ~n5941 ) ;
  assign n5943 = ( x86 & n5680 ) | ( x86 & ~n5806 ) | ( n5680 & ~n5806 ) ;
  assign n5944 = x86 & n5680 ;
  assign n5945 = ( ~n5685 & n5943 ) | ( ~n5685 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5946 = ( n5685 & n5943 ) | ( n5685 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5947 = ( n5685 & n5945 ) | ( n5685 & ~n5946 ) | ( n5945 & ~n5946 ) ;
  assign n5948 = ( x87 & n5942 ) | ( x87 & ~n5947 ) | ( n5942 & ~n5947 ) ;
  assign n5949 = ( x87 & n5686 ) | ( x87 & ~n5806 ) | ( n5686 & ~n5806 ) ;
  assign n5950 = x87 & n5686 ;
  assign n5951 = ( ~n5691 & n5949 ) | ( ~n5691 & n5950 ) | ( n5949 & n5950 ) ;
  assign n5952 = ( n5691 & n5949 ) | ( n5691 & n5950 ) | ( n5949 & n5950 ) ;
  assign n5953 = ( n5691 & n5951 ) | ( n5691 & ~n5952 ) | ( n5951 & ~n5952 ) ;
  assign n5954 = ( x88 & n5948 ) | ( x88 & ~n5953 ) | ( n5948 & ~n5953 ) ;
  assign n5955 = ( x88 & n5692 ) | ( x88 & ~n5806 ) | ( n5692 & ~n5806 ) ;
  assign n5956 = x88 & n5692 ;
  assign n5957 = ( ~n5697 & n5955 ) | ( ~n5697 & n5956 ) | ( n5955 & n5956 ) ;
  assign n5958 = ( n5697 & n5955 ) | ( n5697 & n5956 ) | ( n5955 & n5956 ) ;
  assign n5959 = ( n5697 & n5957 ) | ( n5697 & ~n5958 ) | ( n5957 & ~n5958 ) ;
  assign n5960 = ( x89 & n5954 ) | ( x89 & ~n5959 ) | ( n5954 & ~n5959 ) ;
  assign n5961 = ( x89 & n5698 ) | ( x89 & ~n5806 ) | ( n5698 & ~n5806 ) ;
  assign n5962 = x89 & n5698 ;
  assign n5963 = ( ~n5703 & n5961 ) | ( ~n5703 & n5962 ) | ( n5961 & n5962 ) ;
  assign n5964 = ( n5703 & n5961 ) | ( n5703 & n5962 ) | ( n5961 & n5962 ) ;
  assign n5965 = ( n5703 & n5963 ) | ( n5703 & ~n5964 ) | ( n5963 & ~n5964 ) ;
  assign n5966 = ( x90 & n5960 ) | ( x90 & ~n5965 ) | ( n5960 & ~n5965 ) ;
  assign n5967 = ( x90 & n5704 ) | ( x90 & ~n5806 ) | ( n5704 & ~n5806 ) ;
  assign n5968 = x90 & n5704 ;
  assign n5969 = ( ~n5709 & n5967 ) | ( ~n5709 & n5968 ) | ( n5967 & n5968 ) ;
  assign n5970 = ( n5709 & n5967 ) | ( n5709 & n5968 ) | ( n5967 & n5968 ) ;
  assign n5971 = ( n5709 & n5969 ) | ( n5709 & ~n5970 ) | ( n5969 & ~n5970 ) ;
  assign n5972 = ( x91 & n5966 ) | ( x91 & ~n5971 ) | ( n5966 & ~n5971 ) ;
  assign n5973 = ( x91 & n5710 ) | ( x91 & ~n5806 ) | ( n5710 & ~n5806 ) ;
  assign n5974 = x91 & n5710 ;
  assign n5975 = ( ~n5715 & n5973 ) | ( ~n5715 & n5974 ) | ( n5973 & n5974 ) ;
  assign n5976 = ( n5715 & n5973 ) | ( n5715 & n5974 ) | ( n5973 & n5974 ) ;
  assign n5977 = ( n5715 & n5975 ) | ( n5715 & ~n5976 ) | ( n5975 & ~n5976 ) ;
  assign n5978 = ( x92 & n5972 ) | ( x92 & ~n5977 ) | ( n5972 & ~n5977 ) ;
  assign n5979 = ( x92 & n5716 ) | ( x92 & ~n5806 ) | ( n5716 & ~n5806 ) ;
  assign n5980 = x92 & n5716 ;
  assign n5981 = ( ~n5721 & n5979 ) | ( ~n5721 & n5980 ) | ( n5979 & n5980 ) ;
  assign n5982 = ( n5721 & n5979 ) | ( n5721 & n5980 ) | ( n5979 & n5980 ) ;
  assign n5983 = ( n5721 & n5981 ) | ( n5721 & ~n5982 ) | ( n5981 & ~n5982 ) ;
  assign n5984 = ( x93 & n5978 ) | ( x93 & ~n5983 ) | ( n5978 & ~n5983 ) ;
  assign n5985 = ( x93 & n5722 ) | ( x93 & ~n5806 ) | ( n5722 & ~n5806 ) ;
  assign n5986 = x93 & n5722 ;
  assign n5987 = ( ~n5727 & n5985 ) | ( ~n5727 & n5986 ) | ( n5985 & n5986 ) ;
  assign n5988 = ( n5727 & n5985 ) | ( n5727 & n5986 ) | ( n5985 & n5986 ) ;
  assign n5989 = ( n5727 & n5987 ) | ( n5727 & ~n5988 ) | ( n5987 & ~n5988 ) ;
  assign n5990 = ( x94 & n5984 ) | ( x94 & ~n5989 ) | ( n5984 & ~n5989 ) ;
  assign n5991 = ( x94 & n5728 ) | ( x94 & ~n5806 ) | ( n5728 & ~n5806 ) ;
  assign n5992 = x94 & n5728 ;
  assign n5993 = ( ~n5733 & n5991 ) | ( ~n5733 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5994 = ( n5733 & n5991 ) | ( n5733 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5995 = ( n5733 & n5993 ) | ( n5733 & ~n5994 ) | ( n5993 & ~n5994 ) ;
  assign n5996 = ( x95 & n5990 ) | ( x95 & ~n5995 ) | ( n5990 & ~n5995 ) ;
  assign n5997 = ( x95 & n5734 ) | ( x95 & ~n5806 ) | ( n5734 & ~n5806 ) ;
  assign n5998 = x95 & n5734 ;
  assign n5999 = ( ~n5739 & n5997 ) | ( ~n5739 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = ( n5739 & n5997 ) | ( n5739 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6001 = ( n5739 & n5999 ) | ( n5739 & ~n6000 ) | ( n5999 & ~n6000 ) ;
  assign n6002 = ( x96 & n5996 ) | ( x96 & ~n6001 ) | ( n5996 & ~n6001 ) ;
  assign n6003 = ( x96 & n5740 ) | ( x96 & ~n5806 ) | ( n5740 & ~n5806 ) ;
  assign n6004 = x96 & n5740 ;
  assign n6005 = ( ~n5745 & n6003 ) | ( ~n5745 & n6004 ) | ( n6003 & n6004 ) ;
  assign n6006 = ( n5745 & n6003 ) | ( n5745 & n6004 ) | ( n6003 & n6004 ) ;
  assign n6007 = ( n5745 & n6005 ) | ( n5745 & ~n6006 ) | ( n6005 & ~n6006 ) ;
  assign n6008 = ( x97 & n6002 ) | ( x97 & ~n6007 ) | ( n6002 & ~n6007 ) ;
  assign n6009 = ( x97 & n5746 ) | ( x97 & ~n5806 ) | ( n5746 & ~n5806 ) ;
  assign n6010 = x97 & n5746 ;
  assign n6011 = ( ~n5751 & n6009 ) | ( ~n5751 & n6010 ) | ( n6009 & n6010 ) ;
  assign n6012 = ( n5751 & n6009 ) | ( n5751 & n6010 ) | ( n6009 & n6010 ) ;
  assign n6013 = ( n5751 & n6011 ) | ( n5751 & ~n6012 ) | ( n6011 & ~n6012 ) ;
  assign n6014 = ( x98 & n6008 ) | ( x98 & ~n6013 ) | ( n6008 & ~n6013 ) ;
  assign n6015 = ( x98 & n5752 ) | ( x98 & ~n5806 ) | ( n5752 & ~n5806 ) ;
  assign n6016 = x98 & n5752 ;
  assign n6017 = ( ~n5757 & n6015 ) | ( ~n5757 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6018 = ( n5757 & n6015 ) | ( n5757 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6019 = ( n5757 & n6017 ) | ( n5757 & ~n6018 ) | ( n6017 & ~n6018 ) ;
  assign n6020 = ( x99 & n6014 ) | ( x99 & ~n6019 ) | ( n6014 & ~n6019 ) ;
  assign n6021 = ( x99 & n5758 ) | ( x99 & ~n5806 ) | ( n5758 & ~n5806 ) ;
  assign n6022 = x99 & n5758 ;
  assign n6023 = ( ~n5763 & n6021 ) | ( ~n5763 & n6022 ) | ( n6021 & n6022 ) ;
  assign n6024 = ( n5763 & n6021 ) | ( n5763 & n6022 ) | ( n6021 & n6022 ) ;
  assign n6025 = ( n5763 & n6023 ) | ( n5763 & ~n6024 ) | ( n6023 & ~n6024 ) ;
  assign n6026 = ( x100 & n6020 ) | ( x100 & ~n6025 ) | ( n6020 & ~n6025 ) ;
  assign n6027 = ( x100 & n5764 ) | ( x100 & ~n5806 ) | ( n5764 & ~n5806 ) ;
  assign n6028 = x100 & n5764 ;
  assign n6029 = ( ~n5769 & n6027 ) | ( ~n5769 & n6028 ) | ( n6027 & n6028 ) ;
  assign n6030 = ( n5769 & n6027 ) | ( n5769 & n6028 ) | ( n6027 & n6028 ) ;
  assign n6031 = ( n5769 & n6029 ) | ( n5769 & ~n6030 ) | ( n6029 & ~n6030 ) ;
  assign n6032 = ( x101 & n6026 ) | ( x101 & ~n6031 ) | ( n6026 & ~n6031 ) ;
  assign n6033 = ( x101 & n5770 ) | ( x101 & ~n5806 ) | ( n5770 & ~n5806 ) ;
  assign n6034 = x101 & n5770 ;
  assign n6035 = ( ~n5775 & n6033 ) | ( ~n5775 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6036 = ( n5775 & n6033 ) | ( n5775 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6037 = ( n5775 & n6035 ) | ( n5775 & ~n6036 ) | ( n6035 & ~n6036 ) ;
  assign n6038 = ( x102 & n6032 ) | ( x102 & ~n6037 ) | ( n6032 & ~n6037 ) ;
  assign n6039 = ( x102 & n5776 ) | ( x102 & ~n5806 ) | ( n5776 & ~n5806 ) ;
  assign n6040 = x102 & n5776 ;
  assign n6041 = ( ~n5781 & n6039 ) | ( ~n5781 & n6040 ) | ( n6039 & n6040 ) ;
  assign n6042 = ( n5781 & n6039 ) | ( n5781 & n6040 ) | ( n6039 & n6040 ) ;
  assign n6043 = ( n5781 & n6041 ) | ( n5781 & ~n6042 ) | ( n6041 & ~n6042 ) ;
  assign n6044 = ( x103 & n6038 ) | ( x103 & ~n6043 ) | ( n6038 & ~n6043 ) ;
  assign n6045 = ( x103 & n5782 ) | ( x103 & ~n5806 ) | ( n5782 & ~n5806 ) ;
  assign n6046 = x103 & n5782 ;
  assign n6047 = ( ~n5787 & n6045 ) | ( ~n5787 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6048 = ( n5787 & n6045 ) | ( n5787 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6049 = ( n5787 & n6047 ) | ( n5787 & ~n6048 ) | ( n6047 & ~n6048 ) ;
  assign n6050 = ( x104 & n6044 ) | ( x104 & ~n6049 ) | ( n6044 & ~n6049 ) ;
  assign n6051 = ( x104 & n5788 ) | ( x104 & ~n5806 ) | ( n5788 & ~n5806 ) ;
  assign n6052 = x104 & n5788 ;
  assign n6053 = ( ~n5793 & n6051 ) | ( ~n5793 & n6052 ) | ( n6051 & n6052 ) ;
  assign n6054 = ( n5793 & n6051 ) | ( n5793 & n6052 ) | ( n6051 & n6052 ) ;
  assign n6055 = ( n5793 & n6053 ) | ( n5793 & ~n6054 ) | ( n6053 & ~n6054 ) ;
  assign n6056 = ( x105 & n6050 ) | ( x105 & ~n6055 ) | ( n6050 & ~n6055 ) ;
  assign n6057 = ( x105 & n5794 ) | ( x105 & ~n5806 ) | ( n5794 & ~n5806 ) ;
  assign n6058 = x105 & n5794 ;
  assign n6059 = ( ~n5799 & n6057 ) | ( ~n5799 & n6058 ) | ( n6057 & n6058 ) ;
  assign n6060 = ( n5799 & n6057 ) | ( n5799 & n6058 ) | ( n6057 & n6058 ) ;
  assign n6061 = ( n5799 & n6059 ) | ( n5799 & ~n6060 ) | ( n6059 & ~n6060 ) ;
  assign n6062 = ( x106 & n6056 ) | ( x106 & ~n6061 ) | ( n6056 & ~n6061 ) ;
  assign n6063 = ( x107 & ~n5811 ) | ( x107 & n6062 ) | ( ~n5811 & n6062 ) ;
  assign n6064 = ( x107 & ~n149 ) | ( x107 & n5801 ) | ( ~n149 & n5801 ) ;
  assign n6065 = x107 & n5801 ;
  assign n6066 = ( n5804 & ~n6064 ) | ( n5804 & n6065 ) | ( ~n6064 & n6065 ) ;
  assign n6067 = ( x108 & n6063 ) | ( x108 & ~n6066 ) | ( n6063 & ~n6066 ) ;
  assign n6068 = n148 | n6067 ;
  assign n6069 = ( x107 & n6062 ) | ( x107 & n6068 ) | ( n6062 & n6068 ) ;
  assign n6070 = x107 | n6062 ;
  assign n6071 = ( ~n5811 & n6069 ) | ( ~n5811 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6072 = ( n5811 & n6069 ) | ( n5811 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6073 = ( n5811 & n6071 ) | ( n5811 & ~n6072 ) | ( n6071 & ~n6072 ) ;
  assign n6074 = ~x18 & x64 ;
  assign n6075 = ~x19 & n6068 ;
  assign n6076 = ( x19 & ~x64 ) | ( x19 & n6068 ) | ( ~x64 & n6068 ) ;
  assign n6077 = ( n5812 & ~n6075 ) | ( n5812 & n6076 ) | ( ~n6075 & n6076 ) ;
  assign n6078 = ( x65 & n6074 ) | ( x65 & ~n6077 ) | ( n6074 & ~n6077 ) ;
  assign n6079 = ( x65 & n5812 ) | ( x65 & n6068 ) | ( n5812 & n6068 ) ;
  assign n6080 = x65 | n5812 ;
  assign n6081 = ( ~n5815 & n6079 ) | ( ~n5815 & n6080 ) | ( n6079 & n6080 ) ;
  assign n6082 = ( n5815 & n6079 ) | ( n5815 & n6080 ) | ( n6079 & n6080 ) ;
  assign n6083 = ( n5815 & n6081 ) | ( n5815 & ~n6082 ) | ( n6081 & ~n6082 ) ;
  assign n6084 = ( x66 & n6078 ) | ( x66 & ~n6083 ) | ( n6078 & ~n6083 ) ;
  assign n6085 = ( x66 & n5816 ) | ( x66 & n6068 ) | ( n5816 & n6068 ) ;
  assign n6086 = x66 | n5816 ;
  assign n6087 = ( ~n5821 & n6085 ) | ( ~n5821 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6088 = ( n5821 & n6085 ) | ( n5821 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6089 = ( n5821 & n6087 ) | ( n5821 & ~n6088 ) | ( n6087 & ~n6088 ) ;
  assign n6090 = ( x67 & n6084 ) | ( x67 & ~n6089 ) | ( n6084 & ~n6089 ) ;
  assign n6091 = ( x67 & n5822 ) | ( x67 & ~n6068 ) | ( n5822 & ~n6068 ) ;
  assign n6092 = x67 & n5822 ;
  assign n6093 = ( ~n5827 & n6091 ) | ( ~n5827 & n6092 ) | ( n6091 & n6092 ) ;
  assign n6094 = ( n5827 & n6091 ) | ( n5827 & n6092 ) | ( n6091 & n6092 ) ;
  assign n6095 = ( n5827 & n6093 ) | ( n5827 & ~n6094 ) | ( n6093 & ~n6094 ) ;
  assign n6096 = ( x68 & n6090 ) | ( x68 & ~n6095 ) | ( n6090 & ~n6095 ) ;
  assign n6097 = ( x68 & n5828 ) | ( x68 & ~n6068 ) | ( n5828 & ~n6068 ) ;
  assign n6098 = x68 & n5828 ;
  assign n6099 = ( ~n5833 & n6097 ) | ( ~n5833 & n6098 ) | ( n6097 & n6098 ) ;
  assign n6100 = ( n5833 & n6097 ) | ( n5833 & n6098 ) | ( n6097 & n6098 ) ;
  assign n6101 = ( n5833 & n6099 ) | ( n5833 & ~n6100 ) | ( n6099 & ~n6100 ) ;
  assign n6102 = ( x69 & n6096 ) | ( x69 & ~n6101 ) | ( n6096 & ~n6101 ) ;
  assign n6103 = ( x69 & n5834 ) | ( x69 & ~n6068 ) | ( n5834 & ~n6068 ) ;
  assign n6104 = x69 & n5834 ;
  assign n6105 = ( ~n5839 & n6103 ) | ( ~n5839 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6106 = ( n5839 & n6103 ) | ( n5839 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6107 = ( n5839 & n6105 ) | ( n5839 & ~n6106 ) | ( n6105 & ~n6106 ) ;
  assign n6108 = ( x70 & n6102 ) | ( x70 & ~n6107 ) | ( n6102 & ~n6107 ) ;
  assign n6109 = ( x70 & n5840 ) | ( x70 & ~n6068 ) | ( n5840 & ~n6068 ) ;
  assign n6110 = x70 & n5840 ;
  assign n6111 = ( ~n5845 & n6109 ) | ( ~n5845 & n6110 ) | ( n6109 & n6110 ) ;
  assign n6112 = ( n5845 & n6109 ) | ( n5845 & n6110 ) | ( n6109 & n6110 ) ;
  assign n6113 = ( n5845 & n6111 ) | ( n5845 & ~n6112 ) | ( n6111 & ~n6112 ) ;
  assign n6114 = ( x71 & n6108 ) | ( x71 & ~n6113 ) | ( n6108 & ~n6113 ) ;
  assign n6115 = ( x71 & n5846 ) | ( x71 & ~n6068 ) | ( n5846 & ~n6068 ) ;
  assign n6116 = x71 & n5846 ;
  assign n6117 = ( ~n5851 & n6115 ) | ( ~n5851 & n6116 ) | ( n6115 & n6116 ) ;
  assign n6118 = ( n5851 & n6115 ) | ( n5851 & n6116 ) | ( n6115 & n6116 ) ;
  assign n6119 = ( n5851 & n6117 ) | ( n5851 & ~n6118 ) | ( n6117 & ~n6118 ) ;
  assign n6120 = ( x72 & n6114 ) | ( x72 & ~n6119 ) | ( n6114 & ~n6119 ) ;
  assign n6121 = ( x72 & n5852 ) | ( x72 & ~n6068 ) | ( n5852 & ~n6068 ) ;
  assign n6122 = x72 & n5852 ;
  assign n6123 = ( ~n5857 & n6121 ) | ( ~n5857 & n6122 ) | ( n6121 & n6122 ) ;
  assign n6124 = ( n5857 & n6121 ) | ( n5857 & n6122 ) | ( n6121 & n6122 ) ;
  assign n6125 = ( n5857 & n6123 ) | ( n5857 & ~n6124 ) | ( n6123 & ~n6124 ) ;
  assign n6126 = ( x73 & n6120 ) | ( x73 & ~n6125 ) | ( n6120 & ~n6125 ) ;
  assign n6127 = ( x73 & n5858 ) | ( x73 & ~n6068 ) | ( n5858 & ~n6068 ) ;
  assign n6128 = x73 & n5858 ;
  assign n6129 = ( ~n5863 & n6127 ) | ( ~n5863 & n6128 ) | ( n6127 & n6128 ) ;
  assign n6130 = ( n5863 & n6127 ) | ( n5863 & n6128 ) | ( n6127 & n6128 ) ;
  assign n6131 = ( n5863 & n6129 ) | ( n5863 & ~n6130 ) | ( n6129 & ~n6130 ) ;
  assign n6132 = ( x74 & n6126 ) | ( x74 & ~n6131 ) | ( n6126 & ~n6131 ) ;
  assign n6133 = ( x74 & n5864 ) | ( x74 & ~n6068 ) | ( n5864 & ~n6068 ) ;
  assign n6134 = x74 & n5864 ;
  assign n6135 = ( ~n5869 & n6133 ) | ( ~n5869 & n6134 ) | ( n6133 & n6134 ) ;
  assign n6136 = ( n5869 & n6133 ) | ( n5869 & n6134 ) | ( n6133 & n6134 ) ;
  assign n6137 = ( n5869 & n6135 ) | ( n5869 & ~n6136 ) | ( n6135 & ~n6136 ) ;
  assign n6138 = ( x75 & n6132 ) | ( x75 & ~n6137 ) | ( n6132 & ~n6137 ) ;
  assign n6139 = ( x75 & n5870 ) | ( x75 & ~n6068 ) | ( n5870 & ~n6068 ) ;
  assign n6140 = x75 & n5870 ;
  assign n6141 = ( ~n5875 & n6139 ) | ( ~n5875 & n6140 ) | ( n6139 & n6140 ) ;
  assign n6142 = ( n5875 & n6139 ) | ( n5875 & n6140 ) | ( n6139 & n6140 ) ;
  assign n6143 = ( n5875 & n6141 ) | ( n5875 & ~n6142 ) | ( n6141 & ~n6142 ) ;
  assign n6144 = ( x76 & n6138 ) | ( x76 & ~n6143 ) | ( n6138 & ~n6143 ) ;
  assign n6145 = ( x76 & n5876 ) | ( x76 & ~n6068 ) | ( n5876 & ~n6068 ) ;
  assign n6146 = x76 & n5876 ;
  assign n6147 = ( ~n5881 & n6145 ) | ( ~n5881 & n6146 ) | ( n6145 & n6146 ) ;
  assign n6148 = ( n5881 & n6145 ) | ( n5881 & n6146 ) | ( n6145 & n6146 ) ;
  assign n6149 = ( n5881 & n6147 ) | ( n5881 & ~n6148 ) | ( n6147 & ~n6148 ) ;
  assign n6150 = ( x77 & n6144 ) | ( x77 & ~n6149 ) | ( n6144 & ~n6149 ) ;
  assign n6151 = ( x77 & n5882 ) | ( x77 & ~n6068 ) | ( n5882 & ~n6068 ) ;
  assign n6152 = x77 & n5882 ;
  assign n6153 = ( ~n5887 & n6151 ) | ( ~n5887 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6154 = ( n5887 & n6151 ) | ( n5887 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6155 = ( n5887 & n6153 ) | ( n5887 & ~n6154 ) | ( n6153 & ~n6154 ) ;
  assign n6156 = ( x78 & n6150 ) | ( x78 & ~n6155 ) | ( n6150 & ~n6155 ) ;
  assign n6157 = ( x78 & n5888 ) | ( x78 & ~n6068 ) | ( n5888 & ~n6068 ) ;
  assign n6158 = x78 & n5888 ;
  assign n6159 = ( ~n5893 & n6157 ) | ( ~n5893 & n6158 ) | ( n6157 & n6158 ) ;
  assign n6160 = ( n5893 & n6157 ) | ( n5893 & n6158 ) | ( n6157 & n6158 ) ;
  assign n6161 = ( n5893 & n6159 ) | ( n5893 & ~n6160 ) | ( n6159 & ~n6160 ) ;
  assign n6162 = ( x79 & n6156 ) | ( x79 & ~n6161 ) | ( n6156 & ~n6161 ) ;
  assign n6163 = ( x79 & n5894 ) | ( x79 & ~n6068 ) | ( n5894 & ~n6068 ) ;
  assign n6164 = x79 & n5894 ;
  assign n6165 = ( ~n5899 & n6163 ) | ( ~n5899 & n6164 ) | ( n6163 & n6164 ) ;
  assign n6166 = ( n5899 & n6163 ) | ( n5899 & n6164 ) | ( n6163 & n6164 ) ;
  assign n6167 = ( n5899 & n6165 ) | ( n5899 & ~n6166 ) | ( n6165 & ~n6166 ) ;
  assign n6168 = ( x80 & n6162 ) | ( x80 & ~n6167 ) | ( n6162 & ~n6167 ) ;
  assign n6169 = ( x80 & n5900 ) | ( x80 & ~n6068 ) | ( n5900 & ~n6068 ) ;
  assign n6170 = x80 & n5900 ;
  assign n6171 = ( ~n5905 & n6169 ) | ( ~n5905 & n6170 ) | ( n6169 & n6170 ) ;
  assign n6172 = ( n5905 & n6169 ) | ( n5905 & n6170 ) | ( n6169 & n6170 ) ;
  assign n6173 = ( n5905 & n6171 ) | ( n5905 & ~n6172 ) | ( n6171 & ~n6172 ) ;
  assign n6174 = ( x81 & n6168 ) | ( x81 & ~n6173 ) | ( n6168 & ~n6173 ) ;
  assign n6175 = ( x81 & n5906 ) | ( x81 & ~n6068 ) | ( n5906 & ~n6068 ) ;
  assign n6176 = x81 & n5906 ;
  assign n6177 = ( ~n5911 & n6175 ) | ( ~n5911 & n6176 ) | ( n6175 & n6176 ) ;
  assign n6178 = ( n5911 & n6175 ) | ( n5911 & n6176 ) | ( n6175 & n6176 ) ;
  assign n6179 = ( n5911 & n6177 ) | ( n5911 & ~n6178 ) | ( n6177 & ~n6178 ) ;
  assign n6180 = ( x82 & n6174 ) | ( x82 & ~n6179 ) | ( n6174 & ~n6179 ) ;
  assign n6181 = ( x82 & n5912 ) | ( x82 & ~n6068 ) | ( n5912 & ~n6068 ) ;
  assign n6182 = x82 & n5912 ;
  assign n6183 = ( ~n5917 & n6181 ) | ( ~n5917 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6184 = ( n5917 & n6181 ) | ( n5917 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6185 = ( n5917 & n6183 ) | ( n5917 & ~n6184 ) | ( n6183 & ~n6184 ) ;
  assign n6186 = ( x83 & n6180 ) | ( x83 & ~n6185 ) | ( n6180 & ~n6185 ) ;
  assign n6187 = ( x83 & n5918 ) | ( x83 & ~n6068 ) | ( n5918 & ~n6068 ) ;
  assign n6188 = x83 & n5918 ;
  assign n6189 = ( ~n5923 & n6187 ) | ( ~n5923 & n6188 ) | ( n6187 & n6188 ) ;
  assign n6190 = ( n5923 & n6187 ) | ( n5923 & n6188 ) | ( n6187 & n6188 ) ;
  assign n6191 = ( n5923 & n6189 ) | ( n5923 & ~n6190 ) | ( n6189 & ~n6190 ) ;
  assign n6192 = ( x84 & n6186 ) | ( x84 & ~n6191 ) | ( n6186 & ~n6191 ) ;
  assign n6193 = ( x84 & n5924 ) | ( x84 & ~n6068 ) | ( n5924 & ~n6068 ) ;
  assign n6194 = x84 & n5924 ;
  assign n6195 = ( ~n5929 & n6193 ) | ( ~n5929 & n6194 ) | ( n6193 & n6194 ) ;
  assign n6196 = ( n5929 & n6193 ) | ( n5929 & n6194 ) | ( n6193 & n6194 ) ;
  assign n6197 = ( n5929 & n6195 ) | ( n5929 & ~n6196 ) | ( n6195 & ~n6196 ) ;
  assign n6198 = ( x85 & n6192 ) | ( x85 & ~n6197 ) | ( n6192 & ~n6197 ) ;
  assign n6199 = ( x85 & n5930 ) | ( x85 & ~n6068 ) | ( n5930 & ~n6068 ) ;
  assign n6200 = x85 & n5930 ;
  assign n6201 = ( ~n5935 & n6199 ) | ( ~n5935 & n6200 ) | ( n6199 & n6200 ) ;
  assign n6202 = ( n5935 & n6199 ) | ( n5935 & n6200 ) | ( n6199 & n6200 ) ;
  assign n6203 = ( n5935 & n6201 ) | ( n5935 & ~n6202 ) | ( n6201 & ~n6202 ) ;
  assign n6204 = ( x86 & n6198 ) | ( x86 & ~n6203 ) | ( n6198 & ~n6203 ) ;
  assign n6205 = ( x86 & n5936 ) | ( x86 & ~n6068 ) | ( n5936 & ~n6068 ) ;
  assign n6206 = x86 & n5936 ;
  assign n6207 = ( ~n5941 & n6205 ) | ( ~n5941 & n6206 ) | ( n6205 & n6206 ) ;
  assign n6208 = ( n5941 & n6205 ) | ( n5941 & n6206 ) | ( n6205 & n6206 ) ;
  assign n6209 = ( n5941 & n6207 ) | ( n5941 & ~n6208 ) | ( n6207 & ~n6208 ) ;
  assign n6210 = ( x87 & n6204 ) | ( x87 & ~n6209 ) | ( n6204 & ~n6209 ) ;
  assign n6211 = ( x87 & n5942 ) | ( x87 & ~n6068 ) | ( n5942 & ~n6068 ) ;
  assign n6212 = x87 & n5942 ;
  assign n6213 = ( ~n5947 & n6211 ) | ( ~n5947 & n6212 ) | ( n6211 & n6212 ) ;
  assign n6214 = ( n5947 & n6211 ) | ( n5947 & n6212 ) | ( n6211 & n6212 ) ;
  assign n6215 = ( n5947 & n6213 ) | ( n5947 & ~n6214 ) | ( n6213 & ~n6214 ) ;
  assign n6216 = ( x88 & n6210 ) | ( x88 & ~n6215 ) | ( n6210 & ~n6215 ) ;
  assign n6217 = ( x88 & n5948 ) | ( x88 & ~n6068 ) | ( n5948 & ~n6068 ) ;
  assign n6218 = x88 & n5948 ;
  assign n6219 = ( ~n5953 & n6217 ) | ( ~n5953 & n6218 ) | ( n6217 & n6218 ) ;
  assign n6220 = ( n5953 & n6217 ) | ( n5953 & n6218 ) | ( n6217 & n6218 ) ;
  assign n6221 = ( n5953 & n6219 ) | ( n5953 & ~n6220 ) | ( n6219 & ~n6220 ) ;
  assign n6222 = ( x89 & n6216 ) | ( x89 & ~n6221 ) | ( n6216 & ~n6221 ) ;
  assign n6223 = ( x89 & n5954 ) | ( x89 & ~n6068 ) | ( n5954 & ~n6068 ) ;
  assign n6224 = x89 & n5954 ;
  assign n6225 = ( ~n5959 & n6223 ) | ( ~n5959 & n6224 ) | ( n6223 & n6224 ) ;
  assign n6226 = ( n5959 & n6223 ) | ( n5959 & n6224 ) | ( n6223 & n6224 ) ;
  assign n6227 = ( n5959 & n6225 ) | ( n5959 & ~n6226 ) | ( n6225 & ~n6226 ) ;
  assign n6228 = ( x90 & n6222 ) | ( x90 & ~n6227 ) | ( n6222 & ~n6227 ) ;
  assign n6229 = ( x90 & n5960 ) | ( x90 & ~n6068 ) | ( n5960 & ~n6068 ) ;
  assign n6230 = x90 & n5960 ;
  assign n6231 = ( ~n5965 & n6229 ) | ( ~n5965 & n6230 ) | ( n6229 & n6230 ) ;
  assign n6232 = ( n5965 & n6229 ) | ( n5965 & n6230 ) | ( n6229 & n6230 ) ;
  assign n6233 = ( n5965 & n6231 ) | ( n5965 & ~n6232 ) | ( n6231 & ~n6232 ) ;
  assign n6234 = ( x91 & n6228 ) | ( x91 & ~n6233 ) | ( n6228 & ~n6233 ) ;
  assign n6235 = ( x91 & n5966 ) | ( x91 & ~n6068 ) | ( n5966 & ~n6068 ) ;
  assign n6236 = x91 & n5966 ;
  assign n6237 = ( ~n5971 & n6235 ) | ( ~n5971 & n6236 ) | ( n6235 & n6236 ) ;
  assign n6238 = ( n5971 & n6235 ) | ( n5971 & n6236 ) | ( n6235 & n6236 ) ;
  assign n6239 = ( n5971 & n6237 ) | ( n5971 & ~n6238 ) | ( n6237 & ~n6238 ) ;
  assign n6240 = ( x92 & n6234 ) | ( x92 & ~n6239 ) | ( n6234 & ~n6239 ) ;
  assign n6241 = ( x92 & n5972 ) | ( x92 & ~n6068 ) | ( n5972 & ~n6068 ) ;
  assign n6242 = x92 & n5972 ;
  assign n6243 = ( ~n5977 & n6241 ) | ( ~n5977 & n6242 ) | ( n6241 & n6242 ) ;
  assign n6244 = ( n5977 & n6241 ) | ( n5977 & n6242 ) | ( n6241 & n6242 ) ;
  assign n6245 = ( n5977 & n6243 ) | ( n5977 & ~n6244 ) | ( n6243 & ~n6244 ) ;
  assign n6246 = ( x93 & n6240 ) | ( x93 & ~n6245 ) | ( n6240 & ~n6245 ) ;
  assign n6247 = ( x93 & n5978 ) | ( x93 & ~n6068 ) | ( n5978 & ~n6068 ) ;
  assign n6248 = x93 & n5978 ;
  assign n6249 = ( ~n5983 & n6247 ) | ( ~n5983 & n6248 ) | ( n6247 & n6248 ) ;
  assign n6250 = ( n5983 & n6247 ) | ( n5983 & n6248 ) | ( n6247 & n6248 ) ;
  assign n6251 = ( n5983 & n6249 ) | ( n5983 & ~n6250 ) | ( n6249 & ~n6250 ) ;
  assign n6252 = ( x94 & n6246 ) | ( x94 & ~n6251 ) | ( n6246 & ~n6251 ) ;
  assign n6253 = ( x94 & n5984 ) | ( x94 & ~n6068 ) | ( n5984 & ~n6068 ) ;
  assign n6254 = x94 & n5984 ;
  assign n6255 = ( ~n5989 & n6253 ) | ( ~n5989 & n6254 ) | ( n6253 & n6254 ) ;
  assign n6256 = ( n5989 & n6253 ) | ( n5989 & n6254 ) | ( n6253 & n6254 ) ;
  assign n6257 = ( n5989 & n6255 ) | ( n5989 & ~n6256 ) | ( n6255 & ~n6256 ) ;
  assign n6258 = ( x95 & n6252 ) | ( x95 & ~n6257 ) | ( n6252 & ~n6257 ) ;
  assign n6259 = ( x95 & n5990 ) | ( x95 & ~n6068 ) | ( n5990 & ~n6068 ) ;
  assign n6260 = x95 & n5990 ;
  assign n6261 = ( ~n5995 & n6259 ) | ( ~n5995 & n6260 ) | ( n6259 & n6260 ) ;
  assign n6262 = ( n5995 & n6259 ) | ( n5995 & n6260 ) | ( n6259 & n6260 ) ;
  assign n6263 = ( n5995 & n6261 ) | ( n5995 & ~n6262 ) | ( n6261 & ~n6262 ) ;
  assign n6264 = ( x96 & n6258 ) | ( x96 & ~n6263 ) | ( n6258 & ~n6263 ) ;
  assign n6265 = ( x96 & n5996 ) | ( x96 & ~n6068 ) | ( n5996 & ~n6068 ) ;
  assign n6266 = x96 & n5996 ;
  assign n6267 = ( ~n6001 & n6265 ) | ( ~n6001 & n6266 ) | ( n6265 & n6266 ) ;
  assign n6268 = ( n6001 & n6265 ) | ( n6001 & n6266 ) | ( n6265 & n6266 ) ;
  assign n6269 = ( n6001 & n6267 ) | ( n6001 & ~n6268 ) | ( n6267 & ~n6268 ) ;
  assign n6270 = ( x97 & n6264 ) | ( x97 & ~n6269 ) | ( n6264 & ~n6269 ) ;
  assign n6271 = ( x97 & n6002 ) | ( x97 & ~n6068 ) | ( n6002 & ~n6068 ) ;
  assign n6272 = x97 & n6002 ;
  assign n6273 = ( ~n6007 & n6271 ) | ( ~n6007 & n6272 ) | ( n6271 & n6272 ) ;
  assign n6274 = ( n6007 & n6271 ) | ( n6007 & n6272 ) | ( n6271 & n6272 ) ;
  assign n6275 = ( n6007 & n6273 ) | ( n6007 & ~n6274 ) | ( n6273 & ~n6274 ) ;
  assign n6276 = ( x98 & n6270 ) | ( x98 & ~n6275 ) | ( n6270 & ~n6275 ) ;
  assign n6277 = ( x98 & n6008 ) | ( x98 & ~n6068 ) | ( n6008 & ~n6068 ) ;
  assign n6278 = x98 & n6008 ;
  assign n6279 = ( ~n6013 & n6277 ) | ( ~n6013 & n6278 ) | ( n6277 & n6278 ) ;
  assign n6280 = ( n6013 & n6277 ) | ( n6013 & n6278 ) | ( n6277 & n6278 ) ;
  assign n6281 = ( n6013 & n6279 ) | ( n6013 & ~n6280 ) | ( n6279 & ~n6280 ) ;
  assign n6282 = ( x99 & n6276 ) | ( x99 & ~n6281 ) | ( n6276 & ~n6281 ) ;
  assign n6283 = ( x99 & n6014 ) | ( x99 & ~n6068 ) | ( n6014 & ~n6068 ) ;
  assign n6284 = x99 & n6014 ;
  assign n6285 = ( ~n6019 & n6283 ) | ( ~n6019 & n6284 ) | ( n6283 & n6284 ) ;
  assign n6286 = ( n6019 & n6283 ) | ( n6019 & n6284 ) | ( n6283 & n6284 ) ;
  assign n6287 = ( n6019 & n6285 ) | ( n6019 & ~n6286 ) | ( n6285 & ~n6286 ) ;
  assign n6288 = ( x100 & n6282 ) | ( x100 & ~n6287 ) | ( n6282 & ~n6287 ) ;
  assign n6289 = ( x100 & n6020 ) | ( x100 & ~n6068 ) | ( n6020 & ~n6068 ) ;
  assign n6290 = x100 & n6020 ;
  assign n6291 = ( ~n6025 & n6289 ) | ( ~n6025 & n6290 ) | ( n6289 & n6290 ) ;
  assign n6292 = ( n6025 & n6289 ) | ( n6025 & n6290 ) | ( n6289 & n6290 ) ;
  assign n6293 = ( n6025 & n6291 ) | ( n6025 & ~n6292 ) | ( n6291 & ~n6292 ) ;
  assign n6294 = ( x101 & n6288 ) | ( x101 & ~n6293 ) | ( n6288 & ~n6293 ) ;
  assign n6295 = ( x101 & n6026 ) | ( x101 & ~n6068 ) | ( n6026 & ~n6068 ) ;
  assign n6296 = x101 & n6026 ;
  assign n6297 = ( ~n6031 & n6295 ) | ( ~n6031 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6298 = ( n6031 & n6295 ) | ( n6031 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6299 = ( n6031 & n6297 ) | ( n6031 & ~n6298 ) | ( n6297 & ~n6298 ) ;
  assign n6300 = ( x102 & n6294 ) | ( x102 & ~n6299 ) | ( n6294 & ~n6299 ) ;
  assign n6301 = ( x102 & n6032 ) | ( x102 & ~n6068 ) | ( n6032 & ~n6068 ) ;
  assign n6302 = x102 & n6032 ;
  assign n6303 = ( ~n6037 & n6301 ) | ( ~n6037 & n6302 ) | ( n6301 & n6302 ) ;
  assign n6304 = ( n6037 & n6301 ) | ( n6037 & n6302 ) | ( n6301 & n6302 ) ;
  assign n6305 = ( n6037 & n6303 ) | ( n6037 & ~n6304 ) | ( n6303 & ~n6304 ) ;
  assign n6306 = ( x103 & n6300 ) | ( x103 & ~n6305 ) | ( n6300 & ~n6305 ) ;
  assign n6307 = ( x103 & n6038 ) | ( x103 & ~n6068 ) | ( n6038 & ~n6068 ) ;
  assign n6308 = x103 & n6038 ;
  assign n6309 = ( ~n6043 & n6307 ) | ( ~n6043 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = ( n6043 & n6307 ) | ( n6043 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6311 = ( n6043 & n6309 ) | ( n6043 & ~n6310 ) | ( n6309 & ~n6310 ) ;
  assign n6312 = ( x104 & n6306 ) | ( x104 & ~n6311 ) | ( n6306 & ~n6311 ) ;
  assign n6313 = ( x104 & n6044 ) | ( x104 & ~n6068 ) | ( n6044 & ~n6068 ) ;
  assign n6314 = x104 & n6044 ;
  assign n6315 = ( ~n6049 & n6313 ) | ( ~n6049 & n6314 ) | ( n6313 & n6314 ) ;
  assign n6316 = ( n6049 & n6313 ) | ( n6049 & n6314 ) | ( n6313 & n6314 ) ;
  assign n6317 = ( n6049 & n6315 ) | ( n6049 & ~n6316 ) | ( n6315 & ~n6316 ) ;
  assign n6318 = ( x105 & n6312 ) | ( x105 & ~n6317 ) | ( n6312 & ~n6317 ) ;
  assign n6319 = ( x105 & n6050 ) | ( x105 & ~n6068 ) | ( n6050 & ~n6068 ) ;
  assign n6320 = x105 & n6050 ;
  assign n6321 = ( ~n6055 & n6319 ) | ( ~n6055 & n6320 ) | ( n6319 & n6320 ) ;
  assign n6322 = ( n6055 & n6319 ) | ( n6055 & n6320 ) | ( n6319 & n6320 ) ;
  assign n6323 = ( n6055 & n6321 ) | ( n6055 & ~n6322 ) | ( n6321 & ~n6322 ) ;
  assign n6324 = ( x106 & n6318 ) | ( x106 & ~n6323 ) | ( n6318 & ~n6323 ) ;
  assign n6325 = ( x106 & n6056 ) | ( x106 & ~n6068 ) | ( n6056 & ~n6068 ) ;
  assign n6326 = x106 & n6056 ;
  assign n6327 = ( ~n6061 & n6325 ) | ( ~n6061 & n6326 ) | ( n6325 & n6326 ) ;
  assign n6328 = ( n6061 & n6325 ) | ( n6061 & n6326 ) | ( n6325 & n6326 ) ;
  assign n6329 = ( n6061 & n6327 ) | ( n6061 & ~n6328 ) | ( n6327 & ~n6328 ) ;
  assign n6330 = ( x107 & n6324 ) | ( x107 & ~n6329 ) | ( n6324 & ~n6329 ) ;
  assign n6331 = ( x108 & ~n148 ) | ( x108 & n6063 ) | ( ~n148 & n6063 ) ;
  assign n6332 = x108 & n6063 ;
  assign n6333 = ( n6066 & ~n6331 ) | ( n6066 & n6332 ) | ( ~n6331 & n6332 ) ;
  assign n6334 = ( x108 & ~n6073 ) | ( x108 & n6330 ) | ( ~n6073 & n6330 ) ;
  assign n6335 = ( x109 & ~n6333 ) | ( x109 & n6334 ) | ( ~n6333 & n6334 ) ;
  assign n6336 = n147 | n6335 ;
  assign n6337 = ( x108 & n6330 ) | ( x108 & n6336 ) | ( n6330 & n6336 ) ;
  assign n6338 = x108 | n6330 ;
  assign n6339 = ( ~n6073 & n6337 ) | ( ~n6073 & n6338 ) | ( n6337 & n6338 ) ;
  assign n6340 = ( n6073 & n6337 ) | ( n6073 & n6338 ) | ( n6337 & n6338 ) ;
  assign n6341 = ( n6073 & n6339 ) | ( n6073 & ~n6340 ) | ( n6339 & ~n6340 ) ;
  assign n6342 = ~x17 & x64 ;
  assign n6343 = ~x18 & n6336 ;
  assign n6344 = ( x18 & ~x64 ) | ( x18 & n6336 ) | ( ~x64 & n6336 ) ;
  assign n6345 = ( n6074 & ~n6343 ) | ( n6074 & n6344 ) | ( ~n6343 & n6344 ) ;
  assign n6346 = ( x65 & n6342 ) | ( x65 & ~n6345 ) | ( n6342 & ~n6345 ) ;
  assign n6347 = ( x65 & n6074 ) | ( x65 & n6336 ) | ( n6074 & n6336 ) ;
  assign n6348 = x65 | n6074 ;
  assign n6349 = ( ~n6077 & n6347 ) | ( ~n6077 & n6348 ) | ( n6347 & n6348 ) ;
  assign n6350 = ( n6077 & n6347 ) | ( n6077 & n6348 ) | ( n6347 & n6348 ) ;
  assign n6351 = ( n6077 & n6349 ) | ( n6077 & ~n6350 ) | ( n6349 & ~n6350 ) ;
  assign n6352 = ( x66 & n6346 ) | ( x66 & ~n6351 ) | ( n6346 & ~n6351 ) ;
  assign n6353 = ( x66 & n6078 ) | ( x66 & n6336 ) | ( n6078 & n6336 ) ;
  assign n6354 = x66 | n6078 ;
  assign n6355 = ( ~n6083 & n6353 ) | ( ~n6083 & n6354 ) | ( n6353 & n6354 ) ;
  assign n6356 = ( n6083 & n6353 ) | ( n6083 & n6354 ) | ( n6353 & n6354 ) ;
  assign n6357 = ( n6083 & n6355 ) | ( n6083 & ~n6356 ) | ( n6355 & ~n6356 ) ;
  assign n6358 = ( x67 & n6352 ) | ( x67 & ~n6357 ) | ( n6352 & ~n6357 ) ;
  assign n6359 = ( x67 & n6084 ) | ( x67 & ~n6336 ) | ( n6084 & ~n6336 ) ;
  assign n6360 = x67 & n6084 ;
  assign n6361 = ( ~n6089 & n6359 ) | ( ~n6089 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6362 = ( n6089 & n6359 ) | ( n6089 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6363 = ( n6089 & n6361 ) | ( n6089 & ~n6362 ) | ( n6361 & ~n6362 ) ;
  assign n6364 = ( x68 & n6358 ) | ( x68 & ~n6363 ) | ( n6358 & ~n6363 ) ;
  assign n6365 = ( x68 & n6090 ) | ( x68 & ~n6336 ) | ( n6090 & ~n6336 ) ;
  assign n6366 = x68 & n6090 ;
  assign n6367 = ( ~n6095 & n6365 ) | ( ~n6095 & n6366 ) | ( n6365 & n6366 ) ;
  assign n6368 = ( n6095 & n6365 ) | ( n6095 & n6366 ) | ( n6365 & n6366 ) ;
  assign n6369 = ( n6095 & n6367 ) | ( n6095 & ~n6368 ) | ( n6367 & ~n6368 ) ;
  assign n6370 = ( x69 & n6364 ) | ( x69 & ~n6369 ) | ( n6364 & ~n6369 ) ;
  assign n6371 = ( x69 & n6096 ) | ( x69 & ~n6336 ) | ( n6096 & ~n6336 ) ;
  assign n6372 = x69 & n6096 ;
  assign n6373 = ( ~n6101 & n6371 ) | ( ~n6101 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6374 = ( n6101 & n6371 ) | ( n6101 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6375 = ( n6101 & n6373 ) | ( n6101 & ~n6374 ) | ( n6373 & ~n6374 ) ;
  assign n6376 = ( x70 & n6370 ) | ( x70 & ~n6375 ) | ( n6370 & ~n6375 ) ;
  assign n6377 = ( x70 & n6102 ) | ( x70 & ~n6336 ) | ( n6102 & ~n6336 ) ;
  assign n6378 = x70 & n6102 ;
  assign n6379 = ( ~n6107 & n6377 ) | ( ~n6107 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6380 = ( n6107 & n6377 ) | ( n6107 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6381 = ( n6107 & n6379 ) | ( n6107 & ~n6380 ) | ( n6379 & ~n6380 ) ;
  assign n6382 = ( x71 & n6376 ) | ( x71 & ~n6381 ) | ( n6376 & ~n6381 ) ;
  assign n6383 = ( x71 & n6108 ) | ( x71 & ~n6336 ) | ( n6108 & ~n6336 ) ;
  assign n6384 = x71 & n6108 ;
  assign n6385 = ( ~n6113 & n6383 ) | ( ~n6113 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6386 = ( n6113 & n6383 ) | ( n6113 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6387 = ( n6113 & n6385 ) | ( n6113 & ~n6386 ) | ( n6385 & ~n6386 ) ;
  assign n6388 = ( x72 & n6382 ) | ( x72 & ~n6387 ) | ( n6382 & ~n6387 ) ;
  assign n6389 = ( x72 & n6114 ) | ( x72 & ~n6336 ) | ( n6114 & ~n6336 ) ;
  assign n6390 = x72 & n6114 ;
  assign n6391 = ( ~n6119 & n6389 ) | ( ~n6119 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6392 = ( n6119 & n6389 ) | ( n6119 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6393 = ( n6119 & n6391 ) | ( n6119 & ~n6392 ) | ( n6391 & ~n6392 ) ;
  assign n6394 = ( x73 & n6388 ) | ( x73 & ~n6393 ) | ( n6388 & ~n6393 ) ;
  assign n6395 = ( x73 & n6120 ) | ( x73 & ~n6336 ) | ( n6120 & ~n6336 ) ;
  assign n6396 = x73 & n6120 ;
  assign n6397 = ( ~n6125 & n6395 ) | ( ~n6125 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = ( n6125 & n6395 ) | ( n6125 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6399 = ( n6125 & n6397 ) | ( n6125 & ~n6398 ) | ( n6397 & ~n6398 ) ;
  assign n6400 = ( x74 & n6394 ) | ( x74 & ~n6399 ) | ( n6394 & ~n6399 ) ;
  assign n6401 = ( x74 & n6126 ) | ( x74 & ~n6336 ) | ( n6126 & ~n6336 ) ;
  assign n6402 = x74 & n6126 ;
  assign n6403 = ( ~n6131 & n6401 ) | ( ~n6131 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6404 = ( n6131 & n6401 ) | ( n6131 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6405 = ( n6131 & n6403 ) | ( n6131 & ~n6404 ) | ( n6403 & ~n6404 ) ;
  assign n6406 = ( x75 & n6400 ) | ( x75 & ~n6405 ) | ( n6400 & ~n6405 ) ;
  assign n6407 = ( x75 & n6132 ) | ( x75 & ~n6336 ) | ( n6132 & ~n6336 ) ;
  assign n6408 = x75 & n6132 ;
  assign n6409 = ( ~n6137 & n6407 ) | ( ~n6137 & n6408 ) | ( n6407 & n6408 ) ;
  assign n6410 = ( n6137 & n6407 ) | ( n6137 & n6408 ) | ( n6407 & n6408 ) ;
  assign n6411 = ( n6137 & n6409 ) | ( n6137 & ~n6410 ) | ( n6409 & ~n6410 ) ;
  assign n6412 = ( x76 & n6406 ) | ( x76 & ~n6411 ) | ( n6406 & ~n6411 ) ;
  assign n6413 = ( x76 & n6138 ) | ( x76 & ~n6336 ) | ( n6138 & ~n6336 ) ;
  assign n6414 = x76 & n6138 ;
  assign n6415 = ( ~n6143 & n6413 ) | ( ~n6143 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6416 = ( n6143 & n6413 ) | ( n6143 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6417 = ( n6143 & n6415 ) | ( n6143 & ~n6416 ) | ( n6415 & ~n6416 ) ;
  assign n6418 = ( x77 & n6412 ) | ( x77 & ~n6417 ) | ( n6412 & ~n6417 ) ;
  assign n6419 = ( x77 & n6144 ) | ( x77 & ~n6336 ) | ( n6144 & ~n6336 ) ;
  assign n6420 = x77 & n6144 ;
  assign n6421 = ( ~n6149 & n6419 ) | ( ~n6149 & n6420 ) | ( n6419 & n6420 ) ;
  assign n6422 = ( n6149 & n6419 ) | ( n6149 & n6420 ) | ( n6419 & n6420 ) ;
  assign n6423 = ( n6149 & n6421 ) | ( n6149 & ~n6422 ) | ( n6421 & ~n6422 ) ;
  assign n6424 = ( x78 & n6418 ) | ( x78 & ~n6423 ) | ( n6418 & ~n6423 ) ;
  assign n6425 = ( x78 & n6150 ) | ( x78 & ~n6336 ) | ( n6150 & ~n6336 ) ;
  assign n6426 = x78 & n6150 ;
  assign n6427 = ( ~n6155 & n6425 ) | ( ~n6155 & n6426 ) | ( n6425 & n6426 ) ;
  assign n6428 = ( n6155 & n6425 ) | ( n6155 & n6426 ) | ( n6425 & n6426 ) ;
  assign n6429 = ( n6155 & n6427 ) | ( n6155 & ~n6428 ) | ( n6427 & ~n6428 ) ;
  assign n6430 = ( x79 & n6424 ) | ( x79 & ~n6429 ) | ( n6424 & ~n6429 ) ;
  assign n6431 = ( x79 & n6156 ) | ( x79 & ~n6336 ) | ( n6156 & ~n6336 ) ;
  assign n6432 = x79 & n6156 ;
  assign n6433 = ( ~n6161 & n6431 ) | ( ~n6161 & n6432 ) | ( n6431 & n6432 ) ;
  assign n6434 = ( n6161 & n6431 ) | ( n6161 & n6432 ) | ( n6431 & n6432 ) ;
  assign n6435 = ( n6161 & n6433 ) | ( n6161 & ~n6434 ) | ( n6433 & ~n6434 ) ;
  assign n6436 = ( x80 & n6430 ) | ( x80 & ~n6435 ) | ( n6430 & ~n6435 ) ;
  assign n6437 = ( x80 & n6162 ) | ( x80 & ~n6336 ) | ( n6162 & ~n6336 ) ;
  assign n6438 = x80 & n6162 ;
  assign n6439 = ( ~n6167 & n6437 ) | ( ~n6167 & n6438 ) | ( n6437 & n6438 ) ;
  assign n6440 = ( n6167 & n6437 ) | ( n6167 & n6438 ) | ( n6437 & n6438 ) ;
  assign n6441 = ( n6167 & n6439 ) | ( n6167 & ~n6440 ) | ( n6439 & ~n6440 ) ;
  assign n6442 = ( x81 & n6436 ) | ( x81 & ~n6441 ) | ( n6436 & ~n6441 ) ;
  assign n6443 = ( x81 & n6168 ) | ( x81 & ~n6336 ) | ( n6168 & ~n6336 ) ;
  assign n6444 = x81 & n6168 ;
  assign n6445 = ( ~n6173 & n6443 ) | ( ~n6173 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6446 = ( n6173 & n6443 ) | ( n6173 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6447 = ( n6173 & n6445 ) | ( n6173 & ~n6446 ) | ( n6445 & ~n6446 ) ;
  assign n6448 = ( x82 & n6442 ) | ( x82 & ~n6447 ) | ( n6442 & ~n6447 ) ;
  assign n6449 = ( x82 & n6174 ) | ( x82 & ~n6336 ) | ( n6174 & ~n6336 ) ;
  assign n6450 = x82 & n6174 ;
  assign n6451 = ( ~n6179 & n6449 ) | ( ~n6179 & n6450 ) | ( n6449 & n6450 ) ;
  assign n6452 = ( n6179 & n6449 ) | ( n6179 & n6450 ) | ( n6449 & n6450 ) ;
  assign n6453 = ( n6179 & n6451 ) | ( n6179 & ~n6452 ) | ( n6451 & ~n6452 ) ;
  assign n6454 = ( x83 & n6448 ) | ( x83 & ~n6453 ) | ( n6448 & ~n6453 ) ;
  assign n6455 = ( x83 & n6180 ) | ( x83 & ~n6336 ) | ( n6180 & ~n6336 ) ;
  assign n6456 = x83 & n6180 ;
  assign n6457 = ( ~n6185 & n6455 ) | ( ~n6185 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = ( n6185 & n6455 ) | ( n6185 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6459 = ( n6185 & n6457 ) | ( n6185 & ~n6458 ) | ( n6457 & ~n6458 ) ;
  assign n6460 = ( x84 & n6454 ) | ( x84 & ~n6459 ) | ( n6454 & ~n6459 ) ;
  assign n6461 = ( x84 & n6186 ) | ( x84 & ~n6336 ) | ( n6186 & ~n6336 ) ;
  assign n6462 = x84 & n6186 ;
  assign n6463 = ( ~n6191 & n6461 ) | ( ~n6191 & n6462 ) | ( n6461 & n6462 ) ;
  assign n6464 = ( n6191 & n6461 ) | ( n6191 & n6462 ) | ( n6461 & n6462 ) ;
  assign n6465 = ( n6191 & n6463 ) | ( n6191 & ~n6464 ) | ( n6463 & ~n6464 ) ;
  assign n6466 = ( x85 & n6460 ) | ( x85 & ~n6465 ) | ( n6460 & ~n6465 ) ;
  assign n6467 = ( x85 & n6192 ) | ( x85 & ~n6336 ) | ( n6192 & ~n6336 ) ;
  assign n6468 = x85 & n6192 ;
  assign n6469 = ( ~n6197 & n6467 ) | ( ~n6197 & n6468 ) | ( n6467 & n6468 ) ;
  assign n6470 = ( n6197 & n6467 ) | ( n6197 & n6468 ) | ( n6467 & n6468 ) ;
  assign n6471 = ( n6197 & n6469 ) | ( n6197 & ~n6470 ) | ( n6469 & ~n6470 ) ;
  assign n6472 = ( x86 & n6466 ) | ( x86 & ~n6471 ) | ( n6466 & ~n6471 ) ;
  assign n6473 = ( x86 & n6198 ) | ( x86 & ~n6336 ) | ( n6198 & ~n6336 ) ;
  assign n6474 = x86 & n6198 ;
  assign n6475 = ( ~n6203 & n6473 ) | ( ~n6203 & n6474 ) | ( n6473 & n6474 ) ;
  assign n6476 = ( n6203 & n6473 ) | ( n6203 & n6474 ) | ( n6473 & n6474 ) ;
  assign n6477 = ( n6203 & n6475 ) | ( n6203 & ~n6476 ) | ( n6475 & ~n6476 ) ;
  assign n6478 = ( x87 & n6472 ) | ( x87 & ~n6477 ) | ( n6472 & ~n6477 ) ;
  assign n6479 = ( x87 & n6204 ) | ( x87 & ~n6336 ) | ( n6204 & ~n6336 ) ;
  assign n6480 = x87 & n6204 ;
  assign n6481 = ( ~n6209 & n6479 ) | ( ~n6209 & n6480 ) | ( n6479 & n6480 ) ;
  assign n6482 = ( n6209 & n6479 ) | ( n6209 & n6480 ) | ( n6479 & n6480 ) ;
  assign n6483 = ( n6209 & n6481 ) | ( n6209 & ~n6482 ) | ( n6481 & ~n6482 ) ;
  assign n6484 = ( x88 & n6478 ) | ( x88 & ~n6483 ) | ( n6478 & ~n6483 ) ;
  assign n6485 = ( x88 & n6210 ) | ( x88 & ~n6336 ) | ( n6210 & ~n6336 ) ;
  assign n6486 = x88 & n6210 ;
  assign n6487 = ( ~n6215 & n6485 ) | ( ~n6215 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6488 = ( n6215 & n6485 ) | ( n6215 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6489 = ( n6215 & n6487 ) | ( n6215 & ~n6488 ) | ( n6487 & ~n6488 ) ;
  assign n6490 = ( x89 & n6484 ) | ( x89 & ~n6489 ) | ( n6484 & ~n6489 ) ;
  assign n6491 = ( x89 & n6216 ) | ( x89 & ~n6336 ) | ( n6216 & ~n6336 ) ;
  assign n6492 = x89 & n6216 ;
  assign n6493 = ( ~n6221 & n6491 ) | ( ~n6221 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6494 = ( n6221 & n6491 ) | ( n6221 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6495 = ( n6221 & n6493 ) | ( n6221 & ~n6494 ) | ( n6493 & ~n6494 ) ;
  assign n6496 = ( x90 & n6490 ) | ( x90 & ~n6495 ) | ( n6490 & ~n6495 ) ;
  assign n6497 = ( x90 & n6222 ) | ( x90 & ~n6336 ) | ( n6222 & ~n6336 ) ;
  assign n6498 = x90 & n6222 ;
  assign n6499 = ( ~n6227 & n6497 ) | ( ~n6227 & n6498 ) | ( n6497 & n6498 ) ;
  assign n6500 = ( n6227 & n6497 ) | ( n6227 & n6498 ) | ( n6497 & n6498 ) ;
  assign n6501 = ( n6227 & n6499 ) | ( n6227 & ~n6500 ) | ( n6499 & ~n6500 ) ;
  assign n6502 = ( x91 & n6496 ) | ( x91 & ~n6501 ) | ( n6496 & ~n6501 ) ;
  assign n6503 = ( x91 & n6228 ) | ( x91 & ~n6336 ) | ( n6228 & ~n6336 ) ;
  assign n6504 = x91 & n6228 ;
  assign n6505 = ( ~n6233 & n6503 ) | ( ~n6233 & n6504 ) | ( n6503 & n6504 ) ;
  assign n6506 = ( n6233 & n6503 ) | ( n6233 & n6504 ) | ( n6503 & n6504 ) ;
  assign n6507 = ( n6233 & n6505 ) | ( n6233 & ~n6506 ) | ( n6505 & ~n6506 ) ;
  assign n6508 = ( x92 & n6502 ) | ( x92 & ~n6507 ) | ( n6502 & ~n6507 ) ;
  assign n6509 = ( x92 & n6234 ) | ( x92 & ~n6336 ) | ( n6234 & ~n6336 ) ;
  assign n6510 = x92 & n6234 ;
  assign n6511 = ( ~n6239 & n6509 ) | ( ~n6239 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6512 = ( n6239 & n6509 ) | ( n6239 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6513 = ( n6239 & n6511 ) | ( n6239 & ~n6512 ) | ( n6511 & ~n6512 ) ;
  assign n6514 = ( x93 & n6508 ) | ( x93 & ~n6513 ) | ( n6508 & ~n6513 ) ;
  assign n6515 = ( x93 & n6240 ) | ( x93 & ~n6336 ) | ( n6240 & ~n6336 ) ;
  assign n6516 = x93 & n6240 ;
  assign n6517 = ( ~n6245 & n6515 ) | ( ~n6245 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6518 = ( n6245 & n6515 ) | ( n6245 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6519 = ( n6245 & n6517 ) | ( n6245 & ~n6518 ) | ( n6517 & ~n6518 ) ;
  assign n6520 = ( x94 & n6514 ) | ( x94 & ~n6519 ) | ( n6514 & ~n6519 ) ;
  assign n6521 = ( x94 & n6246 ) | ( x94 & ~n6336 ) | ( n6246 & ~n6336 ) ;
  assign n6522 = x94 & n6246 ;
  assign n6523 = ( ~n6251 & n6521 ) | ( ~n6251 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6524 = ( n6251 & n6521 ) | ( n6251 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6525 = ( n6251 & n6523 ) | ( n6251 & ~n6524 ) | ( n6523 & ~n6524 ) ;
  assign n6526 = ( x95 & n6520 ) | ( x95 & ~n6525 ) | ( n6520 & ~n6525 ) ;
  assign n6527 = ( x95 & n6252 ) | ( x95 & ~n6336 ) | ( n6252 & ~n6336 ) ;
  assign n6528 = x95 & n6252 ;
  assign n6529 = ( ~n6257 & n6527 ) | ( ~n6257 & n6528 ) | ( n6527 & n6528 ) ;
  assign n6530 = ( n6257 & n6527 ) | ( n6257 & n6528 ) | ( n6527 & n6528 ) ;
  assign n6531 = ( n6257 & n6529 ) | ( n6257 & ~n6530 ) | ( n6529 & ~n6530 ) ;
  assign n6532 = ( x96 & n6526 ) | ( x96 & ~n6531 ) | ( n6526 & ~n6531 ) ;
  assign n6533 = ( x96 & n6258 ) | ( x96 & ~n6336 ) | ( n6258 & ~n6336 ) ;
  assign n6534 = x96 & n6258 ;
  assign n6535 = ( ~n6263 & n6533 ) | ( ~n6263 & n6534 ) | ( n6533 & n6534 ) ;
  assign n6536 = ( n6263 & n6533 ) | ( n6263 & n6534 ) | ( n6533 & n6534 ) ;
  assign n6537 = ( n6263 & n6535 ) | ( n6263 & ~n6536 ) | ( n6535 & ~n6536 ) ;
  assign n6538 = ( x97 & n6532 ) | ( x97 & ~n6537 ) | ( n6532 & ~n6537 ) ;
  assign n6539 = ( x97 & n6264 ) | ( x97 & ~n6336 ) | ( n6264 & ~n6336 ) ;
  assign n6540 = x97 & n6264 ;
  assign n6541 = ( ~n6269 & n6539 ) | ( ~n6269 & n6540 ) | ( n6539 & n6540 ) ;
  assign n6542 = ( n6269 & n6539 ) | ( n6269 & n6540 ) | ( n6539 & n6540 ) ;
  assign n6543 = ( n6269 & n6541 ) | ( n6269 & ~n6542 ) | ( n6541 & ~n6542 ) ;
  assign n6544 = ( x98 & n6538 ) | ( x98 & ~n6543 ) | ( n6538 & ~n6543 ) ;
  assign n6545 = ( x98 & n6270 ) | ( x98 & ~n6336 ) | ( n6270 & ~n6336 ) ;
  assign n6546 = x98 & n6270 ;
  assign n6547 = ( ~n6275 & n6545 ) | ( ~n6275 & n6546 ) | ( n6545 & n6546 ) ;
  assign n6548 = ( n6275 & n6545 ) | ( n6275 & n6546 ) | ( n6545 & n6546 ) ;
  assign n6549 = ( n6275 & n6547 ) | ( n6275 & ~n6548 ) | ( n6547 & ~n6548 ) ;
  assign n6550 = ( x99 & n6544 ) | ( x99 & ~n6549 ) | ( n6544 & ~n6549 ) ;
  assign n6551 = ( x99 & n6276 ) | ( x99 & ~n6336 ) | ( n6276 & ~n6336 ) ;
  assign n6552 = x99 & n6276 ;
  assign n6553 = ( ~n6281 & n6551 ) | ( ~n6281 & n6552 ) | ( n6551 & n6552 ) ;
  assign n6554 = ( n6281 & n6551 ) | ( n6281 & n6552 ) | ( n6551 & n6552 ) ;
  assign n6555 = ( n6281 & n6553 ) | ( n6281 & ~n6554 ) | ( n6553 & ~n6554 ) ;
  assign n6556 = ( x100 & n6550 ) | ( x100 & ~n6555 ) | ( n6550 & ~n6555 ) ;
  assign n6557 = ( x100 & n6282 ) | ( x100 & ~n6336 ) | ( n6282 & ~n6336 ) ;
  assign n6558 = x100 & n6282 ;
  assign n6559 = ( ~n6287 & n6557 ) | ( ~n6287 & n6558 ) | ( n6557 & n6558 ) ;
  assign n6560 = ( n6287 & n6557 ) | ( n6287 & n6558 ) | ( n6557 & n6558 ) ;
  assign n6561 = ( n6287 & n6559 ) | ( n6287 & ~n6560 ) | ( n6559 & ~n6560 ) ;
  assign n6562 = ( x101 & n6556 ) | ( x101 & ~n6561 ) | ( n6556 & ~n6561 ) ;
  assign n6563 = ( x101 & n6288 ) | ( x101 & ~n6336 ) | ( n6288 & ~n6336 ) ;
  assign n6564 = x101 & n6288 ;
  assign n6565 = ( ~n6293 & n6563 ) | ( ~n6293 & n6564 ) | ( n6563 & n6564 ) ;
  assign n6566 = ( n6293 & n6563 ) | ( n6293 & n6564 ) | ( n6563 & n6564 ) ;
  assign n6567 = ( n6293 & n6565 ) | ( n6293 & ~n6566 ) | ( n6565 & ~n6566 ) ;
  assign n6568 = ( x102 & n6562 ) | ( x102 & ~n6567 ) | ( n6562 & ~n6567 ) ;
  assign n6569 = ( x102 & n6294 ) | ( x102 & ~n6336 ) | ( n6294 & ~n6336 ) ;
  assign n6570 = x102 & n6294 ;
  assign n6571 = ( ~n6299 & n6569 ) | ( ~n6299 & n6570 ) | ( n6569 & n6570 ) ;
  assign n6572 = ( n6299 & n6569 ) | ( n6299 & n6570 ) | ( n6569 & n6570 ) ;
  assign n6573 = ( n6299 & n6571 ) | ( n6299 & ~n6572 ) | ( n6571 & ~n6572 ) ;
  assign n6574 = ( x103 & n6568 ) | ( x103 & ~n6573 ) | ( n6568 & ~n6573 ) ;
  assign n6575 = ( x103 & n6300 ) | ( x103 & ~n6336 ) | ( n6300 & ~n6336 ) ;
  assign n6576 = x103 & n6300 ;
  assign n6577 = ( ~n6305 & n6575 ) | ( ~n6305 & n6576 ) | ( n6575 & n6576 ) ;
  assign n6578 = ( n6305 & n6575 ) | ( n6305 & n6576 ) | ( n6575 & n6576 ) ;
  assign n6579 = ( n6305 & n6577 ) | ( n6305 & ~n6578 ) | ( n6577 & ~n6578 ) ;
  assign n6580 = ( x104 & n6574 ) | ( x104 & ~n6579 ) | ( n6574 & ~n6579 ) ;
  assign n6581 = ( x104 & n6306 ) | ( x104 & ~n6336 ) | ( n6306 & ~n6336 ) ;
  assign n6582 = x104 & n6306 ;
  assign n6583 = ( ~n6311 & n6581 ) | ( ~n6311 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6584 = ( n6311 & n6581 ) | ( n6311 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6585 = ( n6311 & n6583 ) | ( n6311 & ~n6584 ) | ( n6583 & ~n6584 ) ;
  assign n6586 = ( x105 & n6580 ) | ( x105 & ~n6585 ) | ( n6580 & ~n6585 ) ;
  assign n6587 = ( x105 & n6312 ) | ( x105 & ~n6336 ) | ( n6312 & ~n6336 ) ;
  assign n6588 = x105 & n6312 ;
  assign n6589 = ( ~n6317 & n6587 ) | ( ~n6317 & n6588 ) | ( n6587 & n6588 ) ;
  assign n6590 = ( n6317 & n6587 ) | ( n6317 & n6588 ) | ( n6587 & n6588 ) ;
  assign n6591 = ( n6317 & n6589 ) | ( n6317 & ~n6590 ) | ( n6589 & ~n6590 ) ;
  assign n6592 = ( x106 & n6586 ) | ( x106 & ~n6591 ) | ( n6586 & ~n6591 ) ;
  assign n6593 = ( x106 & n6318 ) | ( x106 & ~n6336 ) | ( n6318 & ~n6336 ) ;
  assign n6594 = x106 & n6318 ;
  assign n6595 = ( ~n6323 & n6593 ) | ( ~n6323 & n6594 ) | ( n6593 & n6594 ) ;
  assign n6596 = ( n6323 & n6593 ) | ( n6323 & n6594 ) | ( n6593 & n6594 ) ;
  assign n6597 = ( n6323 & n6595 ) | ( n6323 & ~n6596 ) | ( n6595 & ~n6596 ) ;
  assign n6598 = ( x107 & n6592 ) | ( x107 & ~n6597 ) | ( n6592 & ~n6597 ) ;
  assign n6599 = ( x107 & n6324 ) | ( x107 & ~n6336 ) | ( n6324 & ~n6336 ) ;
  assign n6600 = x107 & n6324 ;
  assign n6601 = ( ~n6329 & n6599 ) | ( ~n6329 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6602 = ( n6329 & n6599 ) | ( n6329 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6603 = ( n6329 & n6601 ) | ( n6329 & ~n6602 ) | ( n6601 & ~n6602 ) ;
  assign n6604 = ( x108 & n6598 ) | ( x108 & ~n6603 ) | ( n6598 & ~n6603 ) ;
  assign n6605 = ( x109 & ~n6341 ) | ( x109 & n6604 ) | ( ~n6341 & n6604 ) ;
  assign n6606 = ( n146 & n147 ) | ( n146 & ~n6333 ) | ( n147 & ~n6333 ) ;
  assign n6607 = ( ~x109 & n147 ) | ( ~x109 & n6334 ) | ( n147 & n6334 ) ;
  assign n6608 = ( ~x109 & n6333 ) | ( ~x109 & n6334 ) | ( n6333 & n6334 ) ;
  assign n6609 = ~n6607 & n6608 ;
  assign n6610 = ( n6605 & n6606 ) | ( n6605 & ~n6609 ) | ( n6606 & ~n6609 ) ;
  assign n6611 = ( x109 & n6604 ) | ( x109 & n6610 ) | ( n6604 & n6610 ) ;
  assign n6612 = x109 | n6604 ;
  assign n6613 = ( ~n6341 & n6611 ) | ( ~n6341 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = ( n6341 & n6611 ) | ( n6341 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6615 = ( n6341 & n6613 ) | ( n6341 & ~n6614 ) | ( n6613 & ~n6614 ) ;
  assign n6616 = ~x16 & x64 ;
  assign n6617 = ~x17 & n6610 ;
  assign n6618 = ( x17 & ~x64 ) | ( x17 & n6610 ) | ( ~x64 & n6610 ) ;
  assign n6619 = ( n6342 & ~n6617 ) | ( n6342 & n6618 ) | ( ~n6617 & n6618 ) ;
  assign n6620 = ( x65 & n6616 ) | ( x65 & ~n6619 ) | ( n6616 & ~n6619 ) ;
  assign n6621 = ( x65 & n6342 ) | ( x65 & n6610 ) | ( n6342 & n6610 ) ;
  assign n6622 = x65 | n6342 ;
  assign n6623 = ( ~n6345 & n6621 ) | ( ~n6345 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6624 = ( n6345 & n6621 ) | ( n6345 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6625 = ( n6345 & n6623 ) | ( n6345 & ~n6624 ) | ( n6623 & ~n6624 ) ;
  assign n6626 = ( x66 & n6620 ) | ( x66 & ~n6625 ) | ( n6620 & ~n6625 ) ;
  assign n6627 = ( x66 & n6346 ) | ( x66 & n6610 ) | ( n6346 & n6610 ) ;
  assign n6628 = x66 | n6346 ;
  assign n6629 = ( ~n6351 & n6627 ) | ( ~n6351 & n6628 ) | ( n6627 & n6628 ) ;
  assign n6630 = ( n6351 & n6627 ) | ( n6351 & n6628 ) | ( n6627 & n6628 ) ;
  assign n6631 = ( n6351 & n6629 ) | ( n6351 & ~n6630 ) | ( n6629 & ~n6630 ) ;
  assign n6632 = ( x67 & n6626 ) | ( x67 & ~n6631 ) | ( n6626 & ~n6631 ) ;
  assign n6633 = ( x67 & n6352 ) | ( x67 & ~n6610 ) | ( n6352 & ~n6610 ) ;
  assign n6634 = x67 & n6352 ;
  assign n6635 = ( ~n6357 & n6633 ) | ( ~n6357 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6636 = ( n6357 & n6633 ) | ( n6357 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6637 = ( n6357 & n6635 ) | ( n6357 & ~n6636 ) | ( n6635 & ~n6636 ) ;
  assign n6638 = ( x68 & n6632 ) | ( x68 & ~n6637 ) | ( n6632 & ~n6637 ) ;
  assign n6639 = ( x68 & n6358 ) | ( x68 & ~n6610 ) | ( n6358 & ~n6610 ) ;
  assign n6640 = x68 & n6358 ;
  assign n6641 = ( ~n6363 & n6639 ) | ( ~n6363 & n6640 ) | ( n6639 & n6640 ) ;
  assign n6642 = ( n6363 & n6639 ) | ( n6363 & n6640 ) | ( n6639 & n6640 ) ;
  assign n6643 = ( n6363 & n6641 ) | ( n6363 & ~n6642 ) | ( n6641 & ~n6642 ) ;
  assign n6644 = ( x69 & n6638 ) | ( x69 & ~n6643 ) | ( n6638 & ~n6643 ) ;
  assign n6645 = ( x69 & n6364 ) | ( x69 & ~n6610 ) | ( n6364 & ~n6610 ) ;
  assign n6646 = x69 & n6364 ;
  assign n6647 = ( ~n6369 & n6645 ) | ( ~n6369 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6648 = ( n6369 & n6645 ) | ( n6369 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6649 = ( n6369 & n6647 ) | ( n6369 & ~n6648 ) | ( n6647 & ~n6648 ) ;
  assign n6650 = ( x70 & n6644 ) | ( x70 & ~n6649 ) | ( n6644 & ~n6649 ) ;
  assign n6651 = ( x70 & n6370 ) | ( x70 & ~n6610 ) | ( n6370 & ~n6610 ) ;
  assign n6652 = x70 & n6370 ;
  assign n6653 = ( ~n6375 & n6651 ) | ( ~n6375 & n6652 ) | ( n6651 & n6652 ) ;
  assign n6654 = ( n6375 & n6651 ) | ( n6375 & n6652 ) | ( n6651 & n6652 ) ;
  assign n6655 = ( n6375 & n6653 ) | ( n6375 & ~n6654 ) | ( n6653 & ~n6654 ) ;
  assign n6656 = ( x71 & n6650 ) | ( x71 & ~n6655 ) | ( n6650 & ~n6655 ) ;
  assign n6657 = ( x71 & n6376 ) | ( x71 & ~n6610 ) | ( n6376 & ~n6610 ) ;
  assign n6658 = x71 & n6376 ;
  assign n6659 = ( ~n6381 & n6657 ) | ( ~n6381 & n6658 ) | ( n6657 & n6658 ) ;
  assign n6660 = ( n6381 & n6657 ) | ( n6381 & n6658 ) | ( n6657 & n6658 ) ;
  assign n6661 = ( n6381 & n6659 ) | ( n6381 & ~n6660 ) | ( n6659 & ~n6660 ) ;
  assign n6662 = ( x72 & n6656 ) | ( x72 & ~n6661 ) | ( n6656 & ~n6661 ) ;
  assign n6663 = ( x72 & n6382 ) | ( x72 & ~n6610 ) | ( n6382 & ~n6610 ) ;
  assign n6664 = x72 & n6382 ;
  assign n6665 = ( ~n6387 & n6663 ) | ( ~n6387 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = ( n6387 & n6663 ) | ( n6387 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6667 = ( n6387 & n6665 ) | ( n6387 & ~n6666 ) | ( n6665 & ~n6666 ) ;
  assign n6668 = ( x73 & n6662 ) | ( x73 & ~n6667 ) | ( n6662 & ~n6667 ) ;
  assign n6669 = ( x73 & n6388 ) | ( x73 & ~n6610 ) | ( n6388 & ~n6610 ) ;
  assign n6670 = x73 & n6388 ;
  assign n6671 = ( ~n6393 & n6669 ) | ( ~n6393 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6672 = ( n6393 & n6669 ) | ( n6393 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6673 = ( n6393 & n6671 ) | ( n6393 & ~n6672 ) | ( n6671 & ~n6672 ) ;
  assign n6674 = ( x74 & n6668 ) | ( x74 & ~n6673 ) | ( n6668 & ~n6673 ) ;
  assign n6675 = ( x74 & n6394 ) | ( x74 & ~n6610 ) | ( n6394 & ~n6610 ) ;
  assign n6676 = x74 & n6394 ;
  assign n6677 = ( ~n6399 & n6675 ) | ( ~n6399 & n6676 ) | ( n6675 & n6676 ) ;
  assign n6678 = ( n6399 & n6675 ) | ( n6399 & n6676 ) | ( n6675 & n6676 ) ;
  assign n6679 = ( n6399 & n6677 ) | ( n6399 & ~n6678 ) | ( n6677 & ~n6678 ) ;
  assign n6680 = ( x75 & n6674 ) | ( x75 & ~n6679 ) | ( n6674 & ~n6679 ) ;
  assign n6681 = ( x75 & n6400 ) | ( x75 & ~n6610 ) | ( n6400 & ~n6610 ) ;
  assign n6682 = x75 & n6400 ;
  assign n6683 = ( ~n6405 & n6681 ) | ( ~n6405 & n6682 ) | ( n6681 & n6682 ) ;
  assign n6684 = ( n6405 & n6681 ) | ( n6405 & n6682 ) | ( n6681 & n6682 ) ;
  assign n6685 = ( n6405 & n6683 ) | ( n6405 & ~n6684 ) | ( n6683 & ~n6684 ) ;
  assign n6686 = ( x76 & n6680 ) | ( x76 & ~n6685 ) | ( n6680 & ~n6685 ) ;
  assign n6687 = ( x76 & n6406 ) | ( x76 & ~n6610 ) | ( n6406 & ~n6610 ) ;
  assign n6688 = x76 & n6406 ;
  assign n6689 = ( ~n6411 & n6687 ) | ( ~n6411 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6690 = ( n6411 & n6687 ) | ( n6411 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6691 = ( n6411 & n6689 ) | ( n6411 & ~n6690 ) | ( n6689 & ~n6690 ) ;
  assign n6692 = ( x77 & n6686 ) | ( x77 & ~n6691 ) | ( n6686 & ~n6691 ) ;
  assign n6693 = ( x77 & n6412 ) | ( x77 & ~n6610 ) | ( n6412 & ~n6610 ) ;
  assign n6694 = x77 & n6412 ;
  assign n6695 = ( ~n6417 & n6693 ) | ( ~n6417 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6696 = ( n6417 & n6693 ) | ( n6417 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6697 = ( n6417 & n6695 ) | ( n6417 & ~n6696 ) | ( n6695 & ~n6696 ) ;
  assign n6698 = ( x78 & n6692 ) | ( x78 & ~n6697 ) | ( n6692 & ~n6697 ) ;
  assign n6699 = ( x78 & n6418 ) | ( x78 & ~n6610 ) | ( n6418 & ~n6610 ) ;
  assign n6700 = x78 & n6418 ;
  assign n6701 = ( ~n6423 & n6699 ) | ( ~n6423 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6702 = ( n6423 & n6699 ) | ( n6423 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6703 = ( n6423 & n6701 ) | ( n6423 & ~n6702 ) | ( n6701 & ~n6702 ) ;
  assign n6704 = ( x79 & n6698 ) | ( x79 & ~n6703 ) | ( n6698 & ~n6703 ) ;
  assign n6705 = ( x79 & n6424 ) | ( x79 & ~n6610 ) | ( n6424 & ~n6610 ) ;
  assign n6706 = x79 & n6424 ;
  assign n6707 = ( ~n6429 & n6705 ) | ( ~n6429 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6708 = ( n6429 & n6705 ) | ( n6429 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6709 = ( n6429 & n6707 ) | ( n6429 & ~n6708 ) | ( n6707 & ~n6708 ) ;
  assign n6710 = ( x80 & n6704 ) | ( x80 & ~n6709 ) | ( n6704 & ~n6709 ) ;
  assign n6711 = ( x80 & n6430 ) | ( x80 & ~n6610 ) | ( n6430 & ~n6610 ) ;
  assign n6712 = x80 & n6430 ;
  assign n6713 = ( ~n6435 & n6711 ) | ( ~n6435 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6714 = ( n6435 & n6711 ) | ( n6435 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6715 = ( n6435 & n6713 ) | ( n6435 & ~n6714 ) | ( n6713 & ~n6714 ) ;
  assign n6716 = ( x81 & n6710 ) | ( x81 & ~n6715 ) | ( n6710 & ~n6715 ) ;
  assign n6717 = ( x81 & n6436 ) | ( x81 & ~n6610 ) | ( n6436 & ~n6610 ) ;
  assign n6718 = x81 & n6436 ;
  assign n6719 = ( ~n6441 & n6717 ) | ( ~n6441 & n6718 ) | ( n6717 & n6718 ) ;
  assign n6720 = ( n6441 & n6717 ) | ( n6441 & n6718 ) | ( n6717 & n6718 ) ;
  assign n6721 = ( n6441 & n6719 ) | ( n6441 & ~n6720 ) | ( n6719 & ~n6720 ) ;
  assign n6722 = ( x82 & n6716 ) | ( x82 & ~n6721 ) | ( n6716 & ~n6721 ) ;
  assign n6723 = ( x82 & n6442 ) | ( x82 & ~n6610 ) | ( n6442 & ~n6610 ) ;
  assign n6724 = x82 & n6442 ;
  assign n6725 = ( ~n6447 & n6723 ) | ( ~n6447 & n6724 ) | ( n6723 & n6724 ) ;
  assign n6726 = ( n6447 & n6723 ) | ( n6447 & n6724 ) | ( n6723 & n6724 ) ;
  assign n6727 = ( n6447 & n6725 ) | ( n6447 & ~n6726 ) | ( n6725 & ~n6726 ) ;
  assign n6728 = ( x83 & n6722 ) | ( x83 & ~n6727 ) | ( n6722 & ~n6727 ) ;
  assign n6729 = ( x83 & n6448 ) | ( x83 & ~n6610 ) | ( n6448 & ~n6610 ) ;
  assign n6730 = x83 & n6448 ;
  assign n6731 = ( ~n6453 & n6729 ) | ( ~n6453 & n6730 ) | ( n6729 & n6730 ) ;
  assign n6732 = ( n6453 & n6729 ) | ( n6453 & n6730 ) | ( n6729 & n6730 ) ;
  assign n6733 = ( n6453 & n6731 ) | ( n6453 & ~n6732 ) | ( n6731 & ~n6732 ) ;
  assign n6734 = ( x84 & n6728 ) | ( x84 & ~n6733 ) | ( n6728 & ~n6733 ) ;
  assign n6735 = ( x84 & n6454 ) | ( x84 & ~n6610 ) | ( n6454 & ~n6610 ) ;
  assign n6736 = x84 & n6454 ;
  assign n6737 = ( ~n6459 & n6735 ) | ( ~n6459 & n6736 ) | ( n6735 & n6736 ) ;
  assign n6738 = ( n6459 & n6735 ) | ( n6459 & n6736 ) | ( n6735 & n6736 ) ;
  assign n6739 = ( n6459 & n6737 ) | ( n6459 & ~n6738 ) | ( n6737 & ~n6738 ) ;
  assign n6740 = ( x85 & n6734 ) | ( x85 & ~n6739 ) | ( n6734 & ~n6739 ) ;
  assign n6741 = ( x85 & n6460 ) | ( x85 & ~n6610 ) | ( n6460 & ~n6610 ) ;
  assign n6742 = x85 & n6460 ;
  assign n6743 = ( ~n6465 & n6741 ) | ( ~n6465 & n6742 ) | ( n6741 & n6742 ) ;
  assign n6744 = ( n6465 & n6741 ) | ( n6465 & n6742 ) | ( n6741 & n6742 ) ;
  assign n6745 = ( n6465 & n6743 ) | ( n6465 & ~n6744 ) | ( n6743 & ~n6744 ) ;
  assign n6746 = ( x86 & n6740 ) | ( x86 & ~n6745 ) | ( n6740 & ~n6745 ) ;
  assign n6747 = ( x86 & n6466 ) | ( x86 & ~n6610 ) | ( n6466 & ~n6610 ) ;
  assign n6748 = x86 & n6466 ;
  assign n6749 = ( ~n6471 & n6747 ) | ( ~n6471 & n6748 ) | ( n6747 & n6748 ) ;
  assign n6750 = ( n6471 & n6747 ) | ( n6471 & n6748 ) | ( n6747 & n6748 ) ;
  assign n6751 = ( n6471 & n6749 ) | ( n6471 & ~n6750 ) | ( n6749 & ~n6750 ) ;
  assign n6752 = ( x87 & n6746 ) | ( x87 & ~n6751 ) | ( n6746 & ~n6751 ) ;
  assign n6753 = ( x87 & n6472 ) | ( x87 & ~n6610 ) | ( n6472 & ~n6610 ) ;
  assign n6754 = x87 & n6472 ;
  assign n6755 = ( ~n6477 & n6753 ) | ( ~n6477 & n6754 ) | ( n6753 & n6754 ) ;
  assign n6756 = ( n6477 & n6753 ) | ( n6477 & n6754 ) | ( n6753 & n6754 ) ;
  assign n6757 = ( n6477 & n6755 ) | ( n6477 & ~n6756 ) | ( n6755 & ~n6756 ) ;
  assign n6758 = ( x88 & n6752 ) | ( x88 & ~n6757 ) | ( n6752 & ~n6757 ) ;
  assign n6759 = ( x88 & n6478 ) | ( x88 & ~n6610 ) | ( n6478 & ~n6610 ) ;
  assign n6760 = x88 & n6478 ;
  assign n6761 = ( ~n6483 & n6759 ) | ( ~n6483 & n6760 ) | ( n6759 & n6760 ) ;
  assign n6762 = ( n6483 & n6759 ) | ( n6483 & n6760 ) | ( n6759 & n6760 ) ;
  assign n6763 = ( n6483 & n6761 ) | ( n6483 & ~n6762 ) | ( n6761 & ~n6762 ) ;
  assign n6764 = ( x89 & n6758 ) | ( x89 & ~n6763 ) | ( n6758 & ~n6763 ) ;
  assign n6765 = ( x89 & n6484 ) | ( x89 & ~n6610 ) | ( n6484 & ~n6610 ) ;
  assign n6766 = x89 & n6484 ;
  assign n6767 = ( ~n6489 & n6765 ) | ( ~n6489 & n6766 ) | ( n6765 & n6766 ) ;
  assign n6768 = ( n6489 & n6765 ) | ( n6489 & n6766 ) | ( n6765 & n6766 ) ;
  assign n6769 = ( n6489 & n6767 ) | ( n6489 & ~n6768 ) | ( n6767 & ~n6768 ) ;
  assign n6770 = ( x90 & n6764 ) | ( x90 & ~n6769 ) | ( n6764 & ~n6769 ) ;
  assign n6771 = ( x90 & n6490 ) | ( x90 & ~n6610 ) | ( n6490 & ~n6610 ) ;
  assign n6772 = x90 & n6490 ;
  assign n6773 = ( ~n6495 & n6771 ) | ( ~n6495 & n6772 ) | ( n6771 & n6772 ) ;
  assign n6774 = ( n6495 & n6771 ) | ( n6495 & n6772 ) | ( n6771 & n6772 ) ;
  assign n6775 = ( n6495 & n6773 ) | ( n6495 & ~n6774 ) | ( n6773 & ~n6774 ) ;
  assign n6776 = ( x91 & n6770 ) | ( x91 & ~n6775 ) | ( n6770 & ~n6775 ) ;
  assign n6777 = ( x91 & n6496 ) | ( x91 & ~n6610 ) | ( n6496 & ~n6610 ) ;
  assign n6778 = x91 & n6496 ;
  assign n6779 = ( ~n6501 & n6777 ) | ( ~n6501 & n6778 ) | ( n6777 & n6778 ) ;
  assign n6780 = ( n6501 & n6777 ) | ( n6501 & n6778 ) | ( n6777 & n6778 ) ;
  assign n6781 = ( n6501 & n6779 ) | ( n6501 & ~n6780 ) | ( n6779 & ~n6780 ) ;
  assign n6782 = ( x92 & n6776 ) | ( x92 & ~n6781 ) | ( n6776 & ~n6781 ) ;
  assign n6783 = ( x92 & n6502 ) | ( x92 & ~n6610 ) | ( n6502 & ~n6610 ) ;
  assign n6784 = x92 & n6502 ;
  assign n6785 = ( ~n6507 & n6783 ) | ( ~n6507 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6786 = ( n6507 & n6783 ) | ( n6507 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6787 = ( n6507 & n6785 ) | ( n6507 & ~n6786 ) | ( n6785 & ~n6786 ) ;
  assign n6788 = ( x93 & n6782 ) | ( x93 & ~n6787 ) | ( n6782 & ~n6787 ) ;
  assign n6789 = ( x93 & n6508 ) | ( x93 & ~n6610 ) | ( n6508 & ~n6610 ) ;
  assign n6790 = x93 & n6508 ;
  assign n6791 = ( ~n6513 & n6789 ) | ( ~n6513 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6792 = ( n6513 & n6789 ) | ( n6513 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6793 = ( n6513 & n6791 ) | ( n6513 & ~n6792 ) | ( n6791 & ~n6792 ) ;
  assign n6794 = ( x94 & n6788 ) | ( x94 & ~n6793 ) | ( n6788 & ~n6793 ) ;
  assign n6795 = ( x94 & n6514 ) | ( x94 & ~n6610 ) | ( n6514 & ~n6610 ) ;
  assign n6796 = x94 & n6514 ;
  assign n6797 = ( ~n6519 & n6795 ) | ( ~n6519 & n6796 ) | ( n6795 & n6796 ) ;
  assign n6798 = ( n6519 & n6795 ) | ( n6519 & n6796 ) | ( n6795 & n6796 ) ;
  assign n6799 = ( n6519 & n6797 ) | ( n6519 & ~n6798 ) | ( n6797 & ~n6798 ) ;
  assign n6800 = ( x95 & n6794 ) | ( x95 & ~n6799 ) | ( n6794 & ~n6799 ) ;
  assign n6801 = ( x95 & n6520 ) | ( x95 & ~n6610 ) | ( n6520 & ~n6610 ) ;
  assign n6802 = x95 & n6520 ;
  assign n6803 = ( ~n6525 & n6801 ) | ( ~n6525 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6804 = ( n6525 & n6801 ) | ( n6525 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6805 = ( n6525 & n6803 ) | ( n6525 & ~n6804 ) | ( n6803 & ~n6804 ) ;
  assign n6806 = ( x96 & n6800 ) | ( x96 & ~n6805 ) | ( n6800 & ~n6805 ) ;
  assign n6807 = ( x96 & n6526 ) | ( x96 & ~n6610 ) | ( n6526 & ~n6610 ) ;
  assign n6808 = x96 & n6526 ;
  assign n6809 = ( ~n6531 & n6807 ) | ( ~n6531 & n6808 ) | ( n6807 & n6808 ) ;
  assign n6810 = ( n6531 & n6807 ) | ( n6531 & n6808 ) | ( n6807 & n6808 ) ;
  assign n6811 = ( n6531 & n6809 ) | ( n6531 & ~n6810 ) | ( n6809 & ~n6810 ) ;
  assign n6812 = ( x97 & n6806 ) | ( x97 & ~n6811 ) | ( n6806 & ~n6811 ) ;
  assign n6813 = ( x97 & n6532 ) | ( x97 & ~n6610 ) | ( n6532 & ~n6610 ) ;
  assign n6814 = x97 & n6532 ;
  assign n6815 = ( ~n6537 & n6813 ) | ( ~n6537 & n6814 ) | ( n6813 & n6814 ) ;
  assign n6816 = ( n6537 & n6813 ) | ( n6537 & n6814 ) | ( n6813 & n6814 ) ;
  assign n6817 = ( n6537 & n6815 ) | ( n6537 & ~n6816 ) | ( n6815 & ~n6816 ) ;
  assign n6818 = ( x98 & n6812 ) | ( x98 & ~n6817 ) | ( n6812 & ~n6817 ) ;
  assign n6819 = ( x98 & n6538 ) | ( x98 & ~n6610 ) | ( n6538 & ~n6610 ) ;
  assign n6820 = x98 & n6538 ;
  assign n6821 = ( ~n6543 & n6819 ) | ( ~n6543 & n6820 ) | ( n6819 & n6820 ) ;
  assign n6822 = ( n6543 & n6819 ) | ( n6543 & n6820 ) | ( n6819 & n6820 ) ;
  assign n6823 = ( n6543 & n6821 ) | ( n6543 & ~n6822 ) | ( n6821 & ~n6822 ) ;
  assign n6824 = ( x99 & n6818 ) | ( x99 & ~n6823 ) | ( n6818 & ~n6823 ) ;
  assign n6825 = ( x99 & n6544 ) | ( x99 & ~n6610 ) | ( n6544 & ~n6610 ) ;
  assign n6826 = x99 & n6544 ;
  assign n6827 = ( ~n6549 & n6825 ) | ( ~n6549 & n6826 ) | ( n6825 & n6826 ) ;
  assign n6828 = ( n6549 & n6825 ) | ( n6549 & n6826 ) | ( n6825 & n6826 ) ;
  assign n6829 = ( n6549 & n6827 ) | ( n6549 & ~n6828 ) | ( n6827 & ~n6828 ) ;
  assign n6830 = ( x100 & n6824 ) | ( x100 & ~n6829 ) | ( n6824 & ~n6829 ) ;
  assign n6831 = ( x100 & n6550 ) | ( x100 & ~n6610 ) | ( n6550 & ~n6610 ) ;
  assign n6832 = x100 & n6550 ;
  assign n6833 = ( ~n6555 & n6831 ) | ( ~n6555 & n6832 ) | ( n6831 & n6832 ) ;
  assign n6834 = ( n6555 & n6831 ) | ( n6555 & n6832 ) | ( n6831 & n6832 ) ;
  assign n6835 = ( n6555 & n6833 ) | ( n6555 & ~n6834 ) | ( n6833 & ~n6834 ) ;
  assign n6836 = ( x101 & n6830 ) | ( x101 & ~n6835 ) | ( n6830 & ~n6835 ) ;
  assign n6837 = ( x101 & n6556 ) | ( x101 & ~n6610 ) | ( n6556 & ~n6610 ) ;
  assign n6838 = x101 & n6556 ;
  assign n6839 = ( ~n6561 & n6837 ) | ( ~n6561 & n6838 ) | ( n6837 & n6838 ) ;
  assign n6840 = ( n6561 & n6837 ) | ( n6561 & n6838 ) | ( n6837 & n6838 ) ;
  assign n6841 = ( n6561 & n6839 ) | ( n6561 & ~n6840 ) | ( n6839 & ~n6840 ) ;
  assign n6842 = ( x102 & n6836 ) | ( x102 & ~n6841 ) | ( n6836 & ~n6841 ) ;
  assign n6843 = ( x102 & n6562 ) | ( x102 & ~n6610 ) | ( n6562 & ~n6610 ) ;
  assign n6844 = x102 & n6562 ;
  assign n6845 = ( ~n6567 & n6843 ) | ( ~n6567 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6846 = ( n6567 & n6843 ) | ( n6567 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6847 = ( n6567 & n6845 ) | ( n6567 & ~n6846 ) | ( n6845 & ~n6846 ) ;
  assign n6848 = ( x103 & n6842 ) | ( x103 & ~n6847 ) | ( n6842 & ~n6847 ) ;
  assign n6849 = ( x103 & n6568 ) | ( x103 & ~n6610 ) | ( n6568 & ~n6610 ) ;
  assign n6850 = x103 & n6568 ;
  assign n6851 = ( ~n6573 & n6849 ) | ( ~n6573 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6852 = ( n6573 & n6849 ) | ( n6573 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6853 = ( n6573 & n6851 ) | ( n6573 & ~n6852 ) | ( n6851 & ~n6852 ) ;
  assign n6854 = ( x104 & n6848 ) | ( x104 & ~n6853 ) | ( n6848 & ~n6853 ) ;
  assign n6855 = ( x104 & n6574 ) | ( x104 & ~n6610 ) | ( n6574 & ~n6610 ) ;
  assign n6856 = x104 & n6574 ;
  assign n6857 = ( ~n6579 & n6855 ) | ( ~n6579 & n6856 ) | ( n6855 & n6856 ) ;
  assign n6858 = ( n6579 & n6855 ) | ( n6579 & n6856 ) | ( n6855 & n6856 ) ;
  assign n6859 = ( n6579 & n6857 ) | ( n6579 & ~n6858 ) | ( n6857 & ~n6858 ) ;
  assign n6860 = ( x105 & n6854 ) | ( x105 & ~n6859 ) | ( n6854 & ~n6859 ) ;
  assign n6861 = ( x105 & n6580 ) | ( x105 & ~n6610 ) | ( n6580 & ~n6610 ) ;
  assign n6862 = x105 & n6580 ;
  assign n6863 = ( ~n6585 & n6861 ) | ( ~n6585 & n6862 ) | ( n6861 & n6862 ) ;
  assign n6864 = ( n6585 & n6861 ) | ( n6585 & n6862 ) | ( n6861 & n6862 ) ;
  assign n6865 = ( n6585 & n6863 ) | ( n6585 & ~n6864 ) | ( n6863 & ~n6864 ) ;
  assign n6866 = ( x106 & n6860 ) | ( x106 & ~n6865 ) | ( n6860 & ~n6865 ) ;
  assign n6867 = ( x106 & n6586 ) | ( x106 & ~n6610 ) | ( n6586 & ~n6610 ) ;
  assign n6868 = x106 & n6586 ;
  assign n6869 = ( ~n6591 & n6867 ) | ( ~n6591 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6870 = ( n6591 & n6867 ) | ( n6591 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6871 = ( n6591 & n6869 ) | ( n6591 & ~n6870 ) | ( n6869 & ~n6870 ) ;
  assign n6872 = ( x107 & n6866 ) | ( x107 & ~n6871 ) | ( n6866 & ~n6871 ) ;
  assign n6873 = ( x107 & n6592 ) | ( x107 & ~n6610 ) | ( n6592 & ~n6610 ) ;
  assign n6874 = x107 & n6592 ;
  assign n6875 = ( ~n6597 & n6873 ) | ( ~n6597 & n6874 ) | ( n6873 & n6874 ) ;
  assign n6876 = ( n6597 & n6873 ) | ( n6597 & n6874 ) | ( n6873 & n6874 ) ;
  assign n6877 = ( n6597 & n6875 ) | ( n6597 & ~n6876 ) | ( n6875 & ~n6876 ) ;
  assign n6878 = ( x108 & n6872 ) | ( x108 & ~n6877 ) | ( n6872 & ~n6877 ) ;
  assign n6879 = ( x108 & n6598 ) | ( x108 & ~n6610 ) | ( n6598 & ~n6610 ) ;
  assign n6880 = x108 & n6598 ;
  assign n6881 = ( ~n6603 & n6879 ) | ( ~n6603 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6882 = ( n6603 & n6879 ) | ( n6603 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6883 = ( n6603 & n6881 ) | ( n6603 & ~n6882 ) | ( n6881 & ~n6882 ) ;
  assign n6884 = ( x109 & n6878 ) | ( x109 & ~n6883 ) | ( n6878 & ~n6883 ) ;
  assign n6885 = ( x110 & ~n6615 ) | ( x110 & n6884 ) | ( ~n6615 & n6884 ) ;
  assign n6886 = n145 | n6885 ;
  assign n6887 = n146 | n389 ;
  assign n6888 = ( n389 & n6333 ) | ( n389 & n6887 ) | ( n6333 & n6887 ) ;
  assign n6889 = x110 & n6333 ;
  assign n6890 = n6605 & n6889 ;
  assign n6891 = n6888 | n6890 ;
  assign n6892 = ( n146 & n6886 ) | ( n146 & ~n6891 ) | ( n6886 & ~n6891 ) ;
  assign n6893 = ( x110 & n6884 ) | ( x110 & n6892 ) | ( n6884 & n6892 ) ;
  assign n6894 = x110 | n6884 ;
  assign n6895 = ( ~n6615 & n6893 ) | ( ~n6615 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6896 = ( n6615 & n6893 ) | ( n6615 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6897 = ( n6615 & n6895 ) | ( n6615 & ~n6896 ) | ( n6895 & ~n6896 ) ;
  assign n6898 = ~x15 & x64 ;
  assign n6899 = ~x16 & n6892 ;
  assign n6900 = ( x16 & ~x64 ) | ( x16 & n6892 ) | ( ~x64 & n6892 ) ;
  assign n6901 = ( n6616 & ~n6899 ) | ( n6616 & n6900 ) | ( ~n6899 & n6900 ) ;
  assign n6902 = ( x65 & n6898 ) | ( x65 & ~n6901 ) | ( n6898 & ~n6901 ) ;
  assign n6903 = ( x65 & n6616 ) | ( x65 & n6892 ) | ( n6616 & n6892 ) ;
  assign n6904 = x65 | n6616 ;
  assign n6905 = ( ~n6619 & n6903 ) | ( ~n6619 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6906 = ( n6619 & n6903 ) | ( n6619 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6907 = ( n6619 & n6905 ) | ( n6619 & ~n6906 ) | ( n6905 & ~n6906 ) ;
  assign n6908 = ( x66 & n6902 ) | ( x66 & ~n6907 ) | ( n6902 & ~n6907 ) ;
  assign n6909 = ( x66 & n6620 ) | ( x66 & n6892 ) | ( n6620 & n6892 ) ;
  assign n6910 = x66 | n6620 ;
  assign n6911 = ( ~n6625 & n6909 ) | ( ~n6625 & n6910 ) | ( n6909 & n6910 ) ;
  assign n6912 = ( n6625 & n6909 ) | ( n6625 & n6910 ) | ( n6909 & n6910 ) ;
  assign n6913 = ( n6625 & n6911 ) | ( n6625 & ~n6912 ) | ( n6911 & ~n6912 ) ;
  assign n6914 = ( x67 & n6908 ) | ( x67 & ~n6913 ) | ( n6908 & ~n6913 ) ;
  assign n6915 = ( x67 & n6626 ) | ( x67 & ~n6892 ) | ( n6626 & ~n6892 ) ;
  assign n6916 = x67 & n6626 ;
  assign n6917 = ( ~n6631 & n6915 ) | ( ~n6631 & n6916 ) | ( n6915 & n6916 ) ;
  assign n6918 = ( n6631 & n6915 ) | ( n6631 & n6916 ) | ( n6915 & n6916 ) ;
  assign n6919 = ( n6631 & n6917 ) | ( n6631 & ~n6918 ) | ( n6917 & ~n6918 ) ;
  assign n6920 = ( x68 & n6914 ) | ( x68 & ~n6919 ) | ( n6914 & ~n6919 ) ;
  assign n6921 = ( x68 & n6632 ) | ( x68 & ~n6892 ) | ( n6632 & ~n6892 ) ;
  assign n6922 = x68 & n6632 ;
  assign n6923 = ( ~n6637 & n6921 ) | ( ~n6637 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6924 = ( n6637 & n6921 ) | ( n6637 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6925 = ( n6637 & n6923 ) | ( n6637 & ~n6924 ) | ( n6923 & ~n6924 ) ;
  assign n6926 = ( x69 & n6920 ) | ( x69 & ~n6925 ) | ( n6920 & ~n6925 ) ;
  assign n6927 = ( x69 & n6638 ) | ( x69 & ~n6892 ) | ( n6638 & ~n6892 ) ;
  assign n6928 = x69 & n6638 ;
  assign n6929 = ( ~n6643 & n6927 ) | ( ~n6643 & n6928 ) | ( n6927 & n6928 ) ;
  assign n6930 = ( n6643 & n6927 ) | ( n6643 & n6928 ) | ( n6927 & n6928 ) ;
  assign n6931 = ( n6643 & n6929 ) | ( n6643 & ~n6930 ) | ( n6929 & ~n6930 ) ;
  assign n6932 = ( x70 & n6926 ) | ( x70 & ~n6931 ) | ( n6926 & ~n6931 ) ;
  assign n6933 = ( x70 & n6644 ) | ( x70 & ~n6892 ) | ( n6644 & ~n6892 ) ;
  assign n6934 = x70 & n6644 ;
  assign n6935 = ( ~n6649 & n6933 ) | ( ~n6649 & n6934 ) | ( n6933 & n6934 ) ;
  assign n6936 = ( n6649 & n6933 ) | ( n6649 & n6934 ) | ( n6933 & n6934 ) ;
  assign n6937 = ( n6649 & n6935 ) | ( n6649 & ~n6936 ) | ( n6935 & ~n6936 ) ;
  assign n6938 = ( x71 & n6932 ) | ( x71 & ~n6937 ) | ( n6932 & ~n6937 ) ;
  assign n6939 = ( x71 & n6650 ) | ( x71 & ~n6892 ) | ( n6650 & ~n6892 ) ;
  assign n6940 = x71 & n6650 ;
  assign n6941 = ( ~n6655 & n6939 ) | ( ~n6655 & n6940 ) | ( n6939 & n6940 ) ;
  assign n6942 = ( n6655 & n6939 ) | ( n6655 & n6940 ) | ( n6939 & n6940 ) ;
  assign n6943 = ( n6655 & n6941 ) | ( n6655 & ~n6942 ) | ( n6941 & ~n6942 ) ;
  assign n6944 = ( x72 & n6938 ) | ( x72 & ~n6943 ) | ( n6938 & ~n6943 ) ;
  assign n6945 = ( x72 & n6656 ) | ( x72 & ~n6892 ) | ( n6656 & ~n6892 ) ;
  assign n6946 = x72 & n6656 ;
  assign n6947 = ( ~n6661 & n6945 ) | ( ~n6661 & n6946 ) | ( n6945 & n6946 ) ;
  assign n6948 = ( n6661 & n6945 ) | ( n6661 & n6946 ) | ( n6945 & n6946 ) ;
  assign n6949 = ( n6661 & n6947 ) | ( n6661 & ~n6948 ) | ( n6947 & ~n6948 ) ;
  assign n6950 = ( x73 & n6944 ) | ( x73 & ~n6949 ) | ( n6944 & ~n6949 ) ;
  assign n6951 = ( x73 & n6662 ) | ( x73 & ~n6892 ) | ( n6662 & ~n6892 ) ;
  assign n6952 = x73 & n6662 ;
  assign n6953 = ( ~n6667 & n6951 ) | ( ~n6667 & n6952 ) | ( n6951 & n6952 ) ;
  assign n6954 = ( n6667 & n6951 ) | ( n6667 & n6952 ) | ( n6951 & n6952 ) ;
  assign n6955 = ( n6667 & n6953 ) | ( n6667 & ~n6954 ) | ( n6953 & ~n6954 ) ;
  assign n6956 = ( x74 & n6950 ) | ( x74 & ~n6955 ) | ( n6950 & ~n6955 ) ;
  assign n6957 = ( x74 & n6668 ) | ( x74 & ~n6892 ) | ( n6668 & ~n6892 ) ;
  assign n6958 = x74 & n6668 ;
  assign n6959 = ( ~n6673 & n6957 ) | ( ~n6673 & n6958 ) | ( n6957 & n6958 ) ;
  assign n6960 = ( n6673 & n6957 ) | ( n6673 & n6958 ) | ( n6957 & n6958 ) ;
  assign n6961 = ( n6673 & n6959 ) | ( n6673 & ~n6960 ) | ( n6959 & ~n6960 ) ;
  assign n6962 = ( x75 & n6956 ) | ( x75 & ~n6961 ) | ( n6956 & ~n6961 ) ;
  assign n6963 = ( x75 & n6674 ) | ( x75 & ~n6892 ) | ( n6674 & ~n6892 ) ;
  assign n6964 = x75 & n6674 ;
  assign n6965 = ( ~n6679 & n6963 ) | ( ~n6679 & n6964 ) | ( n6963 & n6964 ) ;
  assign n6966 = ( n6679 & n6963 ) | ( n6679 & n6964 ) | ( n6963 & n6964 ) ;
  assign n6967 = ( n6679 & n6965 ) | ( n6679 & ~n6966 ) | ( n6965 & ~n6966 ) ;
  assign n6968 = ( x76 & n6962 ) | ( x76 & ~n6967 ) | ( n6962 & ~n6967 ) ;
  assign n6969 = ( x76 & n6680 ) | ( x76 & ~n6892 ) | ( n6680 & ~n6892 ) ;
  assign n6970 = x76 & n6680 ;
  assign n6971 = ( ~n6685 & n6969 ) | ( ~n6685 & n6970 ) | ( n6969 & n6970 ) ;
  assign n6972 = ( n6685 & n6969 ) | ( n6685 & n6970 ) | ( n6969 & n6970 ) ;
  assign n6973 = ( n6685 & n6971 ) | ( n6685 & ~n6972 ) | ( n6971 & ~n6972 ) ;
  assign n6974 = ( x77 & n6968 ) | ( x77 & ~n6973 ) | ( n6968 & ~n6973 ) ;
  assign n6975 = ( x77 & n6686 ) | ( x77 & ~n6892 ) | ( n6686 & ~n6892 ) ;
  assign n6976 = x77 & n6686 ;
  assign n6977 = ( ~n6691 & n6975 ) | ( ~n6691 & n6976 ) | ( n6975 & n6976 ) ;
  assign n6978 = ( n6691 & n6975 ) | ( n6691 & n6976 ) | ( n6975 & n6976 ) ;
  assign n6979 = ( n6691 & n6977 ) | ( n6691 & ~n6978 ) | ( n6977 & ~n6978 ) ;
  assign n6980 = ( x78 & n6974 ) | ( x78 & ~n6979 ) | ( n6974 & ~n6979 ) ;
  assign n6981 = ( x78 & n6692 ) | ( x78 & ~n6892 ) | ( n6692 & ~n6892 ) ;
  assign n6982 = x78 & n6692 ;
  assign n6983 = ( ~n6697 & n6981 ) | ( ~n6697 & n6982 ) | ( n6981 & n6982 ) ;
  assign n6984 = ( n6697 & n6981 ) | ( n6697 & n6982 ) | ( n6981 & n6982 ) ;
  assign n6985 = ( n6697 & n6983 ) | ( n6697 & ~n6984 ) | ( n6983 & ~n6984 ) ;
  assign n6986 = ( x79 & n6980 ) | ( x79 & ~n6985 ) | ( n6980 & ~n6985 ) ;
  assign n6987 = ( x79 & n6698 ) | ( x79 & ~n6892 ) | ( n6698 & ~n6892 ) ;
  assign n6988 = x79 & n6698 ;
  assign n6989 = ( ~n6703 & n6987 ) | ( ~n6703 & n6988 ) | ( n6987 & n6988 ) ;
  assign n6990 = ( n6703 & n6987 ) | ( n6703 & n6988 ) | ( n6987 & n6988 ) ;
  assign n6991 = ( n6703 & n6989 ) | ( n6703 & ~n6990 ) | ( n6989 & ~n6990 ) ;
  assign n6992 = ( x80 & n6986 ) | ( x80 & ~n6991 ) | ( n6986 & ~n6991 ) ;
  assign n6993 = ( x80 & n6704 ) | ( x80 & ~n6892 ) | ( n6704 & ~n6892 ) ;
  assign n6994 = x80 & n6704 ;
  assign n6995 = ( ~n6709 & n6993 ) | ( ~n6709 & n6994 ) | ( n6993 & n6994 ) ;
  assign n6996 = ( n6709 & n6993 ) | ( n6709 & n6994 ) | ( n6993 & n6994 ) ;
  assign n6997 = ( n6709 & n6995 ) | ( n6709 & ~n6996 ) | ( n6995 & ~n6996 ) ;
  assign n6998 = ( x81 & n6992 ) | ( x81 & ~n6997 ) | ( n6992 & ~n6997 ) ;
  assign n6999 = ( x81 & n6710 ) | ( x81 & ~n6892 ) | ( n6710 & ~n6892 ) ;
  assign n7000 = x81 & n6710 ;
  assign n7001 = ( ~n6715 & n6999 ) | ( ~n6715 & n7000 ) | ( n6999 & n7000 ) ;
  assign n7002 = ( n6715 & n6999 ) | ( n6715 & n7000 ) | ( n6999 & n7000 ) ;
  assign n7003 = ( n6715 & n7001 ) | ( n6715 & ~n7002 ) | ( n7001 & ~n7002 ) ;
  assign n7004 = ( x82 & n6998 ) | ( x82 & ~n7003 ) | ( n6998 & ~n7003 ) ;
  assign n7005 = ( x82 & n6716 ) | ( x82 & ~n6892 ) | ( n6716 & ~n6892 ) ;
  assign n7006 = x82 & n6716 ;
  assign n7007 = ( ~n6721 & n7005 ) | ( ~n6721 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7008 = ( n6721 & n7005 ) | ( n6721 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7009 = ( n6721 & n7007 ) | ( n6721 & ~n7008 ) | ( n7007 & ~n7008 ) ;
  assign n7010 = ( x83 & n7004 ) | ( x83 & ~n7009 ) | ( n7004 & ~n7009 ) ;
  assign n7011 = ( x83 & n6722 ) | ( x83 & ~n6892 ) | ( n6722 & ~n6892 ) ;
  assign n7012 = x83 & n6722 ;
  assign n7013 = ( ~n6727 & n7011 ) | ( ~n6727 & n7012 ) | ( n7011 & n7012 ) ;
  assign n7014 = ( n6727 & n7011 ) | ( n6727 & n7012 ) | ( n7011 & n7012 ) ;
  assign n7015 = ( n6727 & n7013 ) | ( n6727 & ~n7014 ) | ( n7013 & ~n7014 ) ;
  assign n7016 = ( x84 & n7010 ) | ( x84 & ~n7015 ) | ( n7010 & ~n7015 ) ;
  assign n7017 = ( x84 & n6728 ) | ( x84 & ~n6892 ) | ( n6728 & ~n6892 ) ;
  assign n7018 = x84 & n6728 ;
  assign n7019 = ( ~n6733 & n7017 ) | ( ~n6733 & n7018 ) | ( n7017 & n7018 ) ;
  assign n7020 = ( n6733 & n7017 ) | ( n6733 & n7018 ) | ( n7017 & n7018 ) ;
  assign n7021 = ( n6733 & n7019 ) | ( n6733 & ~n7020 ) | ( n7019 & ~n7020 ) ;
  assign n7022 = ( x85 & n7016 ) | ( x85 & ~n7021 ) | ( n7016 & ~n7021 ) ;
  assign n7023 = ( x85 & n6734 ) | ( x85 & ~n6892 ) | ( n6734 & ~n6892 ) ;
  assign n7024 = x85 & n6734 ;
  assign n7025 = ( ~n6739 & n7023 ) | ( ~n6739 & n7024 ) | ( n7023 & n7024 ) ;
  assign n7026 = ( n6739 & n7023 ) | ( n6739 & n7024 ) | ( n7023 & n7024 ) ;
  assign n7027 = ( n6739 & n7025 ) | ( n6739 & ~n7026 ) | ( n7025 & ~n7026 ) ;
  assign n7028 = ( x86 & n7022 ) | ( x86 & ~n7027 ) | ( n7022 & ~n7027 ) ;
  assign n7029 = ( x86 & n6740 ) | ( x86 & ~n6892 ) | ( n6740 & ~n6892 ) ;
  assign n7030 = x86 & n6740 ;
  assign n7031 = ( ~n6745 & n7029 ) | ( ~n6745 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7032 = ( n6745 & n7029 ) | ( n6745 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7033 = ( n6745 & n7031 ) | ( n6745 & ~n7032 ) | ( n7031 & ~n7032 ) ;
  assign n7034 = ( x87 & n7028 ) | ( x87 & ~n7033 ) | ( n7028 & ~n7033 ) ;
  assign n7035 = ( x87 & n6746 ) | ( x87 & ~n6892 ) | ( n6746 & ~n6892 ) ;
  assign n7036 = x87 & n6746 ;
  assign n7037 = ( ~n6751 & n7035 ) | ( ~n6751 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7038 = ( n6751 & n7035 ) | ( n6751 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7039 = ( n6751 & n7037 ) | ( n6751 & ~n7038 ) | ( n7037 & ~n7038 ) ;
  assign n7040 = ( x88 & n7034 ) | ( x88 & ~n7039 ) | ( n7034 & ~n7039 ) ;
  assign n7041 = ( x88 & n6752 ) | ( x88 & ~n6892 ) | ( n6752 & ~n6892 ) ;
  assign n7042 = x88 & n6752 ;
  assign n7043 = ( ~n6757 & n7041 ) | ( ~n6757 & n7042 ) | ( n7041 & n7042 ) ;
  assign n7044 = ( n6757 & n7041 ) | ( n6757 & n7042 ) | ( n7041 & n7042 ) ;
  assign n7045 = ( n6757 & n7043 ) | ( n6757 & ~n7044 ) | ( n7043 & ~n7044 ) ;
  assign n7046 = ( x89 & n7040 ) | ( x89 & ~n7045 ) | ( n7040 & ~n7045 ) ;
  assign n7047 = ( x89 & n6758 ) | ( x89 & ~n6892 ) | ( n6758 & ~n6892 ) ;
  assign n7048 = x89 & n6758 ;
  assign n7049 = ( ~n6763 & n7047 ) | ( ~n6763 & n7048 ) | ( n7047 & n7048 ) ;
  assign n7050 = ( n6763 & n7047 ) | ( n6763 & n7048 ) | ( n7047 & n7048 ) ;
  assign n7051 = ( n6763 & n7049 ) | ( n6763 & ~n7050 ) | ( n7049 & ~n7050 ) ;
  assign n7052 = ( x90 & n7046 ) | ( x90 & ~n7051 ) | ( n7046 & ~n7051 ) ;
  assign n7053 = ( x90 & n6764 ) | ( x90 & ~n6892 ) | ( n6764 & ~n6892 ) ;
  assign n7054 = x90 & n6764 ;
  assign n7055 = ( ~n6769 & n7053 ) | ( ~n6769 & n7054 ) | ( n7053 & n7054 ) ;
  assign n7056 = ( n6769 & n7053 ) | ( n6769 & n7054 ) | ( n7053 & n7054 ) ;
  assign n7057 = ( n6769 & n7055 ) | ( n6769 & ~n7056 ) | ( n7055 & ~n7056 ) ;
  assign n7058 = ( x91 & n7052 ) | ( x91 & ~n7057 ) | ( n7052 & ~n7057 ) ;
  assign n7059 = ( x91 & n6770 ) | ( x91 & ~n6892 ) | ( n6770 & ~n6892 ) ;
  assign n7060 = x91 & n6770 ;
  assign n7061 = ( ~n6775 & n7059 ) | ( ~n6775 & n7060 ) | ( n7059 & n7060 ) ;
  assign n7062 = ( n6775 & n7059 ) | ( n6775 & n7060 ) | ( n7059 & n7060 ) ;
  assign n7063 = ( n6775 & n7061 ) | ( n6775 & ~n7062 ) | ( n7061 & ~n7062 ) ;
  assign n7064 = ( x92 & n7058 ) | ( x92 & ~n7063 ) | ( n7058 & ~n7063 ) ;
  assign n7065 = ( x92 & n6776 ) | ( x92 & ~n6892 ) | ( n6776 & ~n6892 ) ;
  assign n7066 = x92 & n6776 ;
  assign n7067 = ( ~n6781 & n7065 ) | ( ~n6781 & n7066 ) | ( n7065 & n7066 ) ;
  assign n7068 = ( n6781 & n7065 ) | ( n6781 & n7066 ) | ( n7065 & n7066 ) ;
  assign n7069 = ( n6781 & n7067 ) | ( n6781 & ~n7068 ) | ( n7067 & ~n7068 ) ;
  assign n7070 = ( x93 & n7064 ) | ( x93 & ~n7069 ) | ( n7064 & ~n7069 ) ;
  assign n7071 = ( x93 & n6782 ) | ( x93 & ~n6892 ) | ( n6782 & ~n6892 ) ;
  assign n7072 = x93 & n6782 ;
  assign n7073 = ( ~n6787 & n7071 ) | ( ~n6787 & n7072 ) | ( n7071 & n7072 ) ;
  assign n7074 = ( n6787 & n7071 ) | ( n6787 & n7072 ) | ( n7071 & n7072 ) ;
  assign n7075 = ( n6787 & n7073 ) | ( n6787 & ~n7074 ) | ( n7073 & ~n7074 ) ;
  assign n7076 = ( x94 & n7070 ) | ( x94 & ~n7075 ) | ( n7070 & ~n7075 ) ;
  assign n7077 = ( x94 & n6788 ) | ( x94 & ~n6892 ) | ( n6788 & ~n6892 ) ;
  assign n7078 = x94 & n6788 ;
  assign n7079 = ( ~n6793 & n7077 ) | ( ~n6793 & n7078 ) | ( n7077 & n7078 ) ;
  assign n7080 = ( n6793 & n7077 ) | ( n6793 & n7078 ) | ( n7077 & n7078 ) ;
  assign n7081 = ( n6793 & n7079 ) | ( n6793 & ~n7080 ) | ( n7079 & ~n7080 ) ;
  assign n7082 = ( x95 & n7076 ) | ( x95 & ~n7081 ) | ( n7076 & ~n7081 ) ;
  assign n7083 = ( x95 & n6794 ) | ( x95 & ~n6892 ) | ( n6794 & ~n6892 ) ;
  assign n7084 = x95 & n6794 ;
  assign n7085 = ( ~n6799 & n7083 ) | ( ~n6799 & n7084 ) | ( n7083 & n7084 ) ;
  assign n7086 = ( n6799 & n7083 ) | ( n6799 & n7084 ) | ( n7083 & n7084 ) ;
  assign n7087 = ( n6799 & n7085 ) | ( n6799 & ~n7086 ) | ( n7085 & ~n7086 ) ;
  assign n7088 = ( x96 & n7082 ) | ( x96 & ~n7087 ) | ( n7082 & ~n7087 ) ;
  assign n7089 = ( x96 & n6800 ) | ( x96 & ~n6892 ) | ( n6800 & ~n6892 ) ;
  assign n7090 = x96 & n6800 ;
  assign n7091 = ( ~n6805 & n7089 ) | ( ~n6805 & n7090 ) | ( n7089 & n7090 ) ;
  assign n7092 = ( n6805 & n7089 ) | ( n6805 & n7090 ) | ( n7089 & n7090 ) ;
  assign n7093 = ( n6805 & n7091 ) | ( n6805 & ~n7092 ) | ( n7091 & ~n7092 ) ;
  assign n7094 = ( x97 & n7088 ) | ( x97 & ~n7093 ) | ( n7088 & ~n7093 ) ;
  assign n7095 = ( x97 & n6806 ) | ( x97 & ~n6892 ) | ( n6806 & ~n6892 ) ;
  assign n7096 = x97 & n6806 ;
  assign n7097 = ( ~n6811 & n7095 ) | ( ~n6811 & n7096 ) | ( n7095 & n7096 ) ;
  assign n7098 = ( n6811 & n7095 ) | ( n6811 & n7096 ) | ( n7095 & n7096 ) ;
  assign n7099 = ( n6811 & n7097 ) | ( n6811 & ~n7098 ) | ( n7097 & ~n7098 ) ;
  assign n7100 = ( x98 & n7094 ) | ( x98 & ~n7099 ) | ( n7094 & ~n7099 ) ;
  assign n7101 = ( x98 & n6812 ) | ( x98 & ~n6892 ) | ( n6812 & ~n6892 ) ;
  assign n7102 = x98 & n6812 ;
  assign n7103 = ( ~n6817 & n7101 ) | ( ~n6817 & n7102 ) | ( n7101 & n7102 ) ;
  assign n7104 = ( n6817 & n7101 ) | ( n6817 & n7102 ) | ( n7101 & n7102 ) ;
  assign n7105 = ( n6817 & n7103 ) | ( n6817 & ~n7104 ) | ( n7103 & ~n7104 ) ;
  assign n7106 = ( x99 & n7100 ) | ( x99 & ~n7105 ) | ( n7100 & ~n7105 ) ;
  assign n7107 = ( x99 & n6818 ) | ( x99 & ~n6892 ) | ( n6818 & ~n6892 ) ;
  assign n7108 = x99 & n6818 ;
  assign n7109 = ( ~n6823 & n7107 ) | ( ~n6823 & n7108 ) | ( n7107 & n7108 ) ;
  assign n7110 = ( n6823 & n7107 ) | ( n6823 & n7108 ) | ( n7107 & n7108 ) ;
  assign n7111 = ( n6823 & n7109 ) | ( n6823 & ~n7110 ) | ( n7109 & ~n7110 ) ;
  assign n7112 = ( x100 & n7106 ) | ( x100 & ~n7111 ) | ( n7106 & ~n7111 ) ;
  assign n7113 = ( x100 & n6824 ) | ( x100 & ~n6892 ) | ( n6824 & ~n6892 ) ;
  assign n7114 = x100 & n6824 ;
  assign n7115 = ( ~n6829 & n7113 ) | ( ~n6829 & n7114 ) | ( n7113 & n7114 ) ;
  assign n7116 = ( n6829 & n7113 ) | ( n6829 & n7114 ) | ( n7113 & n7114 ) ;
  assign n7117 = ( n6829 & n7115 ) | ( n6829 & ~n7116 ) | ( n7115 & ~n7116 ) ;
  assign n7118 = ( x101 & n7112 ) | ( x101 & ~n7117 ) | ( n7112 & ~n7117 ) ;
  assign n7119 = ( x101 & n6830 ) | ( x101 & ~n6892 ) | ( n6830 & ~n6892 ) ;
  assign n7120 = x101 & n6830 ;
  assign n7121 = ( ~n6835 & n7119 ) | ( ~n6835 & n7120 ) | ( n7119 & n7120 ) ;
  assign n7122 = ( n6835 & n7119 ) | ( n6835 & n7120 ) | ( n7119 & n7120 ) ;
  assign n7123 = ( n6835 & n7121 ) | ( n6835 & ~n7122 ) | ( n7121 & ~n7122 ) ;
  assign n7124 = ( x102 & n7118 ) | ( x102 & ~n7123 ) | ( n7118 & ~n7123 ) ;
  assign n7125 = ( x102 & n6836 ) | ( x102 & ~n6892 ) | ( n6836 & ~n6892 ) ;
  assign n7126 = x102 & n6836 ;
  assign n7127 = ( ~n6841 & n7125 ) | ( ~n6841 & n7126 ) | ( n7125 & n7126 ) ;
  assign n7128 = ( n6841 & n7125 ) | ( n6841 & n7126 ) | ( n7125 & n7126 ) ;
  assign n7129 = ( n6841 & n7127 ) | ( n6841 & ~n7128 ) | ( n7127 & ~n7128 ) ;
  assign n7130 = ( x103 & n7124 ) | ( x103 & ~n7129 ) | ( n7124 & ~n7129 ) ;
  assign n7131 = ( x103 & n6842 ) | ( x103 & ~n6892 ) | ( n6842 & ~n6892 ) ;
  assign n7132 = x103 & n6842 ;
  assign n7133 = ( ~n6847 & n7131 ) | ( ~n6847 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7134 = ( n6847 & n7131 ) | ( n6847 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7135 = ( n6847 & n7133 ) | ( n6847 & ~n7134 ) | ( n7133 & ~n7134 ) ;
  assign n7136 = ( x104 & n7130 ) | ( x104 & ~n7135 ) | ( n7130 & ~n7135 ) ;
  assign n7137 = ( x104 & n6848 ) | ( x104 & ~n6892 ) | ( n6848 & ~n6892 ) ;
  assign n7138 = x104 & n6848 ;
  assign n7139 = ( ~n6853 & n7137 ) | ( ~n6853 & n7138 ) | ( n7137 & n7138 ) ;
  assign n7140 = ( n6853 & n7137 ) | ( n6853 & n7138 ) | ( n7137 & n7138 ) ;
  assign n7141 = ( n6853 & n7139 ) | ( n6853 & ~n7140 ) | ( n7139 & ~n7140 ) ;
  assign n7142 = ( x105 & n7136 ) | ( x105 & ~n7141 ) | ( n7136 & ~n7141 ) ;
  assign n7143 = ( x105 & n6854 ) | ( x105 & ~n6892 ) | ( n6854 & ~n6892 ) ;
  assign n7144 = x105 & n6854 ;
  assign n7145 = ( ~n6859 & n7143 ) | ( ~n6859 & n7144 ) | ( n7143 & n7144 ) ;
  assign n7146 = ( n6859 & n7143 ) | ( n6859 & n7144 ) | ( n7143 & n7144 ) ;
  assign n7147 = ( n6859 & n7145 ) | ( n6859 & ~n7146 ) | ( n7145 & ~n7146 ) ;
  assign n7148 = ( x106 & n7142 ) | ( x106 & ~n7147 ) | ( n7142 & ~n7147 ) ;
  assign n7149 = ( x106 & n6860 ) | ( x106 & ~n6892 ) | ( n6860 & ~n6892 ) ;
  assign n7150 = x106 & n6860 ;
  assign n7151 = ( ~n6865 & n7149 ) | ( ~n6865 & n7150 ) | ( n7149 & n7150 ) ;
  assign n7152 = ( n6865 & n7149 ) | ( n6865 & n7150 ) | ( n7149 & n7150 ) ;
  assign n7153 = ( n6865 & n7151 ) | ( n6865 & ~n7152 ) | ( n7151 & ~n7152 ) ;
  assign n7154 = ( x107 & n7148 ) | ( x107 & ~n7153 ) | ( n7148 & ~n7153 ) ;
  assign n7155 = ( x107 & n6866 ) | ( x107 & ~n6892 ) | ( n6866 & ~n6892 ) ;
  assign n7156 = x107 & n6866 ;
  assign n7157 = ( ~n6871 & n7155 ) | ( ~n6871 & n7156 ) | ( n7155 & n7156 ) ;
  assign n7158 = ( n6871 & n7155 ) | ( n6871 & n7156 ) | ( n7155 & n7156 ) ;
  assign n7159 = ( n6871 & n7157 ) | ( n6871 & ~n7158 ) | ( n7157 & ~n7158 ) ;
  assign n7160 = ( x108 & n7154 ) | ( x108 & ~n7159 ) | ( n7154 & ~n7159 ) ;
  assign n7161 = ( x108 & n6872 ) | ( x108 & ~n6892 ) | ( n6872 & ~n6892 ) ;
  assign n7162 = x108 & n6872 ;
  assign n7163 = ( ~n6877 & n7161 ) | ( ~n6877 & n7162 ) | ( n7161 & n7162 ) ;
  assign n7164 = ( n6877 & n7161 ) | ( n6877 & n7162 ) | ( n7161 & n7162 ) ;
  assign n7165 = ( n6877 & n7163 ) | ( n6877 & ~n7164 ) | ( n7163 & ~n7164 ) ;
  assign n7166 = ( x109 & n7160 ) | ( x109 & ~n7165 ) | ( n7160 & ~n7165 ) ;
  assign n7167 = ( x109 & n6878 ) | ( x109 & ~n6892 ) | ( n6878 & ~n6892 ) ;
  assign n7168 = x109 & n6878 ;
  assign n7169 = ( ~n6883 & n7167 ) | ( ~n6883 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7170 = ( n6883 & n7167 ) | ( n6883 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7171 = ( n6883 & n7169 ) | ( n6883 & ~n7170 ) | ( n7169 & ~n7170 ) ;
  assign n7172 = ( x110 & n7166 ) | ( x110 & ~n7171 ) | ( n7166 & ~n7171 ) ;
  assign n7173 = ~x111 & n6888 ;
  assign n7174 = ( n6886 & n6888 ) | ( n6886 & n7173 ) | ( n6888 & n7173 ) ;
  assign n7175 = ( x111 & ~n6897 ) | ( x111 & n7172 ) | ( ~n6897 & n7172 ) ;
  assign n7176 = ( x112 & ~n7174 ) | ( x112 & n7175 ) | ( ~n7174 & n7175 ) ;
  assign n7177 = n144 | n7176 ;
  assign n7178 = ( x111 & n7172 ) | ( x111 & n7177 ) | ( n7172 & n7177 ) ;
  assign n7179 = x111 | n7172 ;
  assign n7180 = ( ~n6897 & n7178 ) | ( ~n6897 & n7179 ) | ( n7178 & n7179 ) ;
  assign n7181 = ( n6897 & n7178 ) | ( n6897 & n7179 ) | ( n7178 & n7179 ) ;
  assign n7182 = ( n6897 & n7180 ) | ( n6897 & ~n7181 ) | ( n7180 & ~n7181 ) ;
  assign n7183 = ~x14 & x64 ;
  assign n7184 = ~x15 & n7177 ;
  assign n7185 = ( x15 & ~x64 ) | ( x15 & n7177 ) | ( ~x64 & n7177 ) ;
  assign n7186 = ( n6898 & ~n7184 ) | ( n6898 & n7185 ) | ( ~n7184 & n7185 ) ;
  assign n7187 = ( x65 & n7183 ) | ( x65 & ~n7186 ) | ( n7183 & ~n7186 ) ;
  assign n7188 = ( x65 & n6898 ) | ( x65 & n7177 ) | ( n6898 & n7177 ) ;
  assign n7189 = x65 | n6898 ;
  assign n7190 = ( ~n6901 & n7188 ) | ( ~n6901 & n7189 ) | ( n7188 & n7189 ) ;
  assign n7191 = ( n6901 & n7188 ) | ( n6901 & n7189 ) | ( n7188 & n7189 ) ;
  assign n7192 = ( n6901 & n7190 ) | ( n6901 & ~n7191 ) | ( n7190 & ~n7191 ) ;
  assign n7193 = ( x66 & n7187 ) | ( x66 & ~n7192 ) | ( n7187 & ~n7192 ) ;
  assign n7194 = ( x66 & n6902 ) | ( x66 & n7177 ) | ( n6902 & n7177 ) ;
  assign n7195 = x66 | n6902 ;
  assign n7196 = ( ~n6907 & n7194 ) | ( ~n6907 & n7195 ) | ( n7194 & n7195 ) ;
  assign n7197 = ( n6907 & n7194 ) | ( n6907 & n7195 ) | ( n7194 & n7195 ) ;
  assign n7198 = ( n6907 & n7196 ) | ( n6907 & ~n7197 ) | ( n7196 & ~n7197 ) ;
  assign n7199 = ( x67 & n7193 ) | ( x67 & ~n7198 ) | ( n7193 & ~n7198 ) ;
  assign n7200 = ( x67 & n6908 ) | ( x67 & ~n7177 ) | ( n6908 & ~n7177 ) ;
  assign n7201 = x67 & n6908 ;
  assign n7202 = ( ~n6913 & n7200 ) | ( ~n6913 & n7201 ) | ( n7200 & n7201 ) ;
  assign n7203 = ( n6913 & n7200 ) | ( n6913 & n7201 ) | ( n7200 & n7201 ) ;
  assign n7204 = ( n6913 & n7202 ) | ( n6913 & ~n7203 ) | ( n7202 & ~n7203 ) ;
  assign n7205 = ( x68 & n7199 ) | ( x68 & ~n7204 ) | ( n7199 & ~n7204 ) ;
  assign n7206 = ( x68 & n6914 ) | ( x68 & ~n7177 ) | ( n6914 & ~n7177 ) ;
  assign n7207 = x68 & n6914 ;
  assign n7208 = ( ~n6919 & n7206 ) | ( ~n6919 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( n6919 & n7206 ) | ( n6919 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7210 = ( n6919 & n7208 ) | ( n6919 & ~n7209 ) | ( n7208 & ~n7209 ) ;
  assign n7211 = ( x69 & n7205 ) | ( x69 & ~n7210 ) | ( n7205 & ~n7210 ) ;
  assign n7212 = ( x69 & n6920 ) | ( x69 & ~n7177 ) | ( n6920 & ~n7177 ) ;
  assign n7213 = x69 & n6920 ;
  assign n7214 = ( ~n6925 & n7212 ) | ( ~n6925 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7215 = ( n6925 & n7212 ) | ( n6925 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7216 = ( n6925 & n7214 ) | ( n6925 & ~n7215 ) | ( n7214 & ~n7215 ) ;
  assign n7217 = ( x70 & n7211 ) | ( x70 & ~n7216 ) | ( n7211 & ~n7216 ) ;
  assign n7218 = ( x70 & n6926 ) | ( x70 & ~n7177 ) | ( n6926 & ~n7177 ) ;
  assign n7219 = x70 & n6926 ;
  assign n7220 = ( ~n6931 & n7218 ) | ( ~n6931 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7221 = ( n6931 & n7218 ) | ( n6931 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7222 = ( n6931 & n7220 ) | ( n6931 & ~n7221 ) | ( n7220 & ~n7221 ) ;
  assign n7223 = ( x71 & n7217 ) | ( x71 & ~n7222 ) | ( n7217 & ~n7222 ) ;
  assign n7224 = ( x71 & n6932 ) | ( x71 & ~n7177 ) | ( n6932 & ~n7177 ) ;
  assign n7225 = x71 & n6932 ;
  assign n7226 = ( ~n6937 & n7224 ) | ( ~n6937 & n7225 ) | ( n7224 & n7225 ) ;
  assign n7227 = ( n6937 & n7224 ) | ( n6937 & n7225 ) | ( n7224 & n7225 ) ;
  assign n7228 = ( n6937 & n7226 ) | ( n6937 & ~n7227 ) | ( n7226 & ~n7227 ) ;
  assign n7229 = ( x72 & n7223 ) | ( x72 & ~n7228 ) | ( n7223 & ~n7228 ) ;
  assign n7230 = ( x72 & n6938 ) | ( x72 & ~n7177 ) | ( n6938 & ~n7177 ) ;
  assign n7231 = x72 & n6938 ;
  assign n7232 = ( ~n6943 & n7230 ) | ( ~n6943 & n7231 ) | ( n7230 & n7231 ) ;
  assign n7233 = ( n6943 & n7230 ) | ( n6943 & n7231 ) | ( n7230 & n7231 ) ;
  assign n7234 = ( n6943 & n7232 ) | ( n6943 & ~n7233 ) | ( n7232 & ~n7233 ) ;
  assign n7235 = ( x73 & n7229 ) | ( x73 & ~n7234 ) | ( n7229 & ~n7234 ) ;
  assign n7236 = ( x73 & n6944 ) | ( x73 & ~n7177 ) | ( n6944 & ~n7177 ) ;
  assign n7237 = x73 & n6944 ;
  assign n7238 = ( ~n6949 & n7236 ) | ( ~n6949 & n7237 ) | ( n7236 & n7237 ) ;
  assign n7239 = ( n6949 & n7236 ) | ( n6949 & n7237 ) | ( n7236 & n7237 ) ;
  assign n7240 = ( n6949 & n7238 ) | ( n6949 & ~n7239 ) | ( n7238 & ~n7239 ) ;
  assign n7241 = ( x74 & n7235 ) | ( x74 & ~n7240 ) | ( n7235 & ~n7240 ) ;
  assign n7242 = ( x74 & n6950 ) | ( x74 & ~n7177 ) | ( n6950 & ~n7177 ) ;
  assign n7243 = x74 & n6950 ;
  assign n7244 = ( ~n6955 & n7242 ) | ( ~n6955 & n7243 ) | ( n7242 & n7243 ) ;
  assign n7245 = ( n6955 & n7242 ) | ( n6955 & n7243 ) | ( n7242 & n7243 ) ;
  assign n7246 = ( n6955 & n7244 ) | ( n6955 & ~n7245 ) | ( n7244 & ~n7245 ) ;
  assign n7247 = ( x75 & n7241 ) | ( x75 & ~n7246 ) | ( n7241 & ~n7246 ) ;
  assign n7248 = ( x75 & n6956 ) | ( x75 & ~n7177 ) | ( n6956 & ~n7177 ) ;
  assign n7249 = x75 & n6956 ;
  assign n7250 = ( ~n6961 & n7248 ) | ( ~n6961 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7251 = ( n6961 & n7248 ) | ( n6961 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7252 = ( n6961 & n7250 ) | ( n6961 & ~n7251 ) | ( n7250 & ~n7251 ) ;
  assign n7253 = ( x76 & n7247 ) | ( x76 & ~n7252 ) | ( n7247 & ~n7252 ) ;
  assign n7254 = ( x76 & n6962 ) | ( x76 & ~n7177 ) | ( n6962 & ~n7177 ) ;
  assign n7255 = x76 & n6962 ;
  assign n7256 = ( ~n6967 & n7254 ) | ( ~n6967 & n7255 ) | ( n7254 & n7255 ) ;
  assign n7257 = ( n6967 & n7254 ) | ( n6967 & n7255 ) | ( n7254 & n7255 ) ;
  assign n7258 = ( n6967 & n7256 ) | ( n6967 & ~n7257 ) | ( n7256 & ~n7257 ) ;
  assign n7259 = ( x77 & n7253 ) | ( x77 & ~n7258 ) | ( n7253 & ~n7258 ) ;
  assign n7260 = ( x77 & n6968 ) | ( x77 & ~n7177 ) | ( n6968 & ~n7177 ) ;
  assign n7261 = x77 & n6968 ;
  assign n7262 = ( ~n6973 & n7260 ) | ( ~n6973 & n7261 ) | ( n7260 & n7261 ) ;
  assign n7263 = ( n6973 & n7260 ) | ( n6973 & n7261 ) | ( n7260 & n7261 ) ;
  assign n7264 = ( n6973 & n7262 ) | ( n6973 & ~n7263 ) | ( n7262 & ~n7263 ) ;
  assign n7265 = ( x78 & n7259 ) | ( x78 & ~n7264 ) | ( n7259 & ~n7264 ) ;
  assign n7266 = ( x78 & n6974 ) | ( x78 & ~n7177 ) | ( n6974 & ~n7177 ) ;
  assign n7267 = x78 & n6974 ;
  assign n7268 = ( ~n6979 & n7266 ) | ( ~n6979 & n7267 ) | ( n7266 & n7267 ) ;
  assign n7269 = ( n6979 & n7266 ) | ( n6979 & n7267 ) | ( n7266 & n7267 ) ;
  assign n7270 = ( n6979 & n7268 ) | ( n6979 & ~n7269 ) | ( n7268 & ~n7269 ) ;
  assign n7271 = ( x79 & n7265 ) | ( x79 & ~n7270 ) | ( n7265 & ~n7270 ) ;
  assign n7272 = ( x79 & n6980 ) | ( x79 & ~n7177 ) | ( n6980 & ~n7177 ) ;
  assign n7273 = x79 & n6980 ;
  assign n7274 = ( ~n6985 & n7272 ) | ( ~n6985 & n7273 ) | ( n7272 & n7273 ) ;
  assign n7275 = ( n6985 & n7272 ) | ( n6985 & n7273 ) | ( n7272 & n7273 ) ;
  assign n7276 = ( n6985 & n7274 ) | ( n6985 & ~n7275 ) | ( n7274 & ~n7275 ) ;
  assign n7277 = ( x80 & n7271 ) | ( x80 & ~n7276 ) | ( n7271 & ~n7276 ) ;
  assign n7278 = ( x80 & n6986 ) | ( x80 & ~n7177 ) | ( n6986 & ~n7177 ) ;
  assign n7279 = x80 & n6986 ;
  assign n7280 = ( ~n6991 & n7278 ) | ( ~n6991 & n7279 ) | ( n7278 & n7279 ) ;
  assign n7281 = ( n6991 & n7278 ) | ( n6991 & n7279 ) | ( n7278 & n7279 ) ;
  assign n7282 = ( n6991 & n7280 ) | ( n6991 & ~n7281 ) | ( n7280 & ~n7281 ) ;
  assign n7283 = ( x81 & n7277 ) | ( x81 & ~n7282 ) | ( n7277 & ~n7282 ) ;
  assign n7284 = ( x81 & n6992 ) | ( x81 & ~n7177 ) | ( n6992 & ~n7177 ) ;
  assign n7285 = x81 & n6992 ;
  assign n7286 = ( ~n6997 & n7284 ) | ( ~n6997 & n7285 ) | ( n7284 & n7285 ) ;
  assign n7287 = ( n6997 & n7284 ) | ( n6997 & n7285 ) | ( n7284 & n7285 ) ;
  assign n7288 = ( n6997 & n7286 ) | ( n6997 & ~n7287 ) | ( n7286 & ~n7287 ) ;
  assign n7289 = ( x82 & n7283 ) | ( x82 & ~n7288 ) | ( n7283 & ~n7288 ) ;
  assign n7290 = ( x82 & n6998 ) | ( x82 & ~n7177 ) | ( n6998 & ~n7177 ) ;
  assign n7291 = x82 & n6998 ;
  assign n7292 = ( ~n7003 & n7290 ) | ( ~n7003 & n7291 ) | ( n7290 & n7291 ) ;
  assign n7293 = ( n7003 & n7290 ) | ( n7003 & n7291 ) | ( n7290 & n7291 ) ;
  assign n7294 = ( n7003 & n7292 ) | ( n7003 & ~n7293 ) | ( n7292 & ~n7293 ) ;
  assign n7295 = ( x83 & n7289 ) | ( x83 & ~n7294 ) | ( n7289 & ~n7294 ) ;
  assign n7296 = ( x83 & n7004 ) | ( x83 & ~n7177 ) | ( n7004 & ~n7177 ) ;
  assign n7297 = x83 & n7004 ;
  assign n7298 = ( ~n7009 & n7296 ) | ( ~n7009 & n7297 ) | ( n7296 & n7297 ) ;
  assign n7299 = ( n7009 & n7296 ) | ( n7009 & n7297 ) | ( n7296 & n7297 ) ;
  assign n7300 = ( n7009 & n7298 ) | ( n7009 & ~n7299 ) | ( n7298 & ~n7299 ) ;
  assign n7301 = ( x84 & n7295 ) | ( x84 & ~n7300 ) | ( n7295 & ~n7300 ) ;
  assign n7302 = ( x84 & n7010 ) | ( x84 & ~n7177 ) | ( n7010 & ~n7177 ) ;
  assign n7303 = x84 & n7010 ;
  assign n7304 = ( ~n7015 & n7302 ) | ( ~n7015 & n7303 ) | ( n7302 & n7303 ) ;
  assign n7305 = ( n7015 & n7302 ) | ( n7015 & n7303 ) | ( n7302 & n7303 ) ;
  assign n7306 = ( n7015 & n7304 ) | ( n7015 & ~n7305 ) | ( n7304 & ~n7305 ) ;
  assign n7307 = ( x85 & n7301 ) | ( x85 & ~n7306 ) | ( n7301 & ~n7306 ) ;
  assign n7308 = ( x85 & n7016 ) | ( x85 & ~n7177 ) | ( n7016 & ~n7177 ) ;
  assign n7309 = x85 & n7016 ;
  assign n7310 = ( ~n7021 & n7308 ) | ( ~n7021 & n7309 ) | ( n7308 & n7309 ) ;
  assign n7311 = ( n7021 & n7308 ) | ( n7021 & n7309 ) | ( n7308 & n7309 ) ;
  assign n7312 = ( n7021 & n7310 ) | ( n7021 & ~n7311 ) | ( n7310 & ~n7311 ) ;
  assign n7313 = ( x86 & n7307 ) | ( x86 & ~n7312 ) | ( n7307 & ~n7312 ) ;
  assign n7314 = ( x86 & n7022 ) | ( x86 & ~n7177 ) | ( n7022 & ~n7177 ) ;
  assign n7315 = x86 & n7022 ;
  assign n7316 = ( ~n7027 & n7314 ) | ( ~n7027 & n7315 ) | ( n7314 & n7315 ) ;
  assign n7317 = ( n7027 & n7314 ) | ( n7027 & n7315 ) | ( n7314 & n7315 ) ;
  assign n7318 = ( n7027 & n7316 ) | ( n7027 & ~n7317 ) | ( n7316 & ~n7317 ) ;
  assign n7319 = ( x87 & n7313 ) | ( x87 & ~n7318 ) | ( n7313 & ~n7318 ) ;
  assign n7320 = ( x87 & n7028 ) | ( x87 & ~n7177 ) | ( n7028 & ~n7177 ) ;
  assign n7321 = x87 & n7028 ;
  assign n7322 = ( ~n7033 & n7320 ) | ( ~n7033 & n7321 ) | ( n7320 & n7321 ) ;
  assign n7323 = ( n7033 & n7320 ) | ( n7033 & n7321 ) | ( n7320 & n7321 ) ;
  assign n7324 = ( n7033 & n7322 ) | ( n7033 & ~n7323 ) | ( n7322 & ~n7323 ) ;
  assign n7325 = ( x88 & n7319 ) | ( x88 & ~n7324 ) | ( n7319 & ~n7324 ) ;
  assign n7326 = ( x88 & n7034 ) | ( x88 & ~n7177 ) | ( n7034 & ~n7177 ) ;
  assign n7327 = x88 & n7034 ;
  assign n7328 = ( ~n7039 & n7326 ) | ( ~n7039 & n7327 ) | ( n7326 & n7327 ) ;
  assign n7329 = ( n7039 & n7326 ) | ( n7039 & n7327 ) | ( n7326 & n7327 ) ;
  assign n7330 = ( n7039 & n7328 ) | ( n7039 & ~n7329 ) | ( n7328 & ~n7329 ) ;
  assign n7331 = ( x89 & n7325 ) | ( x89 & ~n7330 ) | ( n7325 & ~n7330 ) ;
  assign n7332 = ( x89 & n7040 ) | ( x89 & ~n7177 ) | ( n7040 & ~n7177 ) ;
  assign n7333 = x89 & n7040 ;
  assign n7334 = ( ~n7045 & n7332 ) | ( ~n7045 & n7333 ) | ( n7332 & n7333 ) ;
  assign n7335 = ( n7045 & n7332 ) | ( n7045 & n7333 ) | ( n7332 & n7333 ) ;
  assign n7336 = ( n7045 & n7334 ) | ( n7045 & ~n7335 ) | ( n7334 & ~n7335 ) ;
  assign n7337 = ( x90 & n7331 ) | ( x90 & ~n7336 ) | ( n7331 & ~n7336 ) ;
  assign n7338 = ( x90 & n7046 ) | ( x90 & ~n7177 ) | ( n7046 & ~n7177 ) ;
  assign n7339 = x90 & n7046 ;
  assign n7340 = ( ~n7051 & n7338 ) | ( ~n7051 & n7339 ) | ( n7338 & n7339 ) ;
  assign n7341 = ( n7051 & n7338 ) | ( n7051 & n7339 ) | ( n7338 & n7339 ) ;
  assign n7342 = ( n7051 & n7340 ) | ( n7051 & ~n7341 ) | ( n7340 & ~n7341 ) ;
  assign n7343 = ( x91 & n7337 ) | ( x91 & ~n7342 ) | ( n7337 & ~n7342 ) ;
  assign n7344 = ( x91 & n7052 ) | ( x91 & ~n7177 ) | ( n7052 & ~n7177 ) ;
  assign n7345 = x91 & n7052 ;
  assign n7346 = ( ~n7057 & n7344 ) | ( ~n7057 & n7345 ) | ( n7344 & n7345 ) ;
  assign n7347 = ( n7057 & n7344 ) | ( n7057 & n7345 ) | ( n7344 & n7345 ) ;
  assign n7348 = ( n7057 & n7346 ) | ( n7057 & ~n7347 ) | ( n7346 & ~n7347 ) ;
  assign n7349 = ( x92 & n7343 ) | ( x92 & ~n7348 ) | ( n7343 & ~n7348 ) ;
  assign n7350 = ( x92 & n7058 ) | ( x92 & ~n7177 ) | ( n7058 & ~n7177 ) ;
  assign n7351 = x92 & n7058 ;
  assign n7352 = ( ~n7063 & n7350 ) | ( ~n7063 & n7351 ) | ( n7350 & n7351 ) ;
  assign n7353 = ( n7063 & n7350 ) | ( n7063 & n7351 ) | ( n7350 & n7351 ) ;
  assign n7354 = ( n7063 & n7352 ) | ( n7063 & ~n7353 ) | ( n7352 & ~n7353 ) ;
  assign n7355 = ( x93 & n7349 ) | ( x93 & ~n7354 ) | ( n7349 & ~n7354 ) ;
  assign n7356 = ( x93 & n7064 ) | ( x93 & ~n7177 ) | ( n7064 & ~n7177 ) ;
  assign n7357 = x93 & n7064 ;
  assign n7358 = ( ~n7069 & n7356 ) | ( ~n7069 & n7357 ) | ( n7356 & n7357 ) ;
  assign n7359 = ( n7069 & n7356 ) | ( n7069 & n7357 ) | ( n7356 & n7357 ) ;
  assign n7360 = ( n7069 & n7358 ) | ( n7069 & ~n7359 ) | ( n7358 & ~n7359 ) ;
  assign n7361 = ( x94 & n7355 ) | ( x94 & ~n7360 ) | ( n7355 & ~n7360 ) ;
  assign n7362 = ( x94 & n7070 ) | ( x94 & ~n7177 ) | ( n7070 & ~n7177 ) ;
  assign n7363 = x94 & n7070 ;
  assign n7364 = ( ~n7075 & n7362 ) | ( ~n7075 & n7363 ) | ( n7362 & n7363 ) ;
  assign n7365 = ( n7075 & n7362 ) | ( n7075 & n7363 ) | ( n7362 & n7363 ) ;
  assign n7366 = ( n7075 & n7364 ) | ( n7075 & ~n7365 ) | ( n7364 & ~n7365 ) ;
  assign n7367 = ( x95 & n7361 ) | ( x95 & ~n7366 ) | ( n7361 & ~n7366 ) ;
  assign n7368 = ( x95 & n7076 ) | ( x95 & ~n7177 ) | ( n7076 & ~n7177 ) ;
  assign n7369 = x95 & n7076 ;
  assign n7370 = ( ~n7081 & n7368 ) | ( ~n7081 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7371 = ( n7081 & n7368 ) | ( n7081 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7372 = ( n7081 & n7370 ) | ( n7081 & ~n7371 ) | ( n7370 & ~n7371 ) ;
  assign n7373 = ( x96 & n7367 ) | ( x96 & ~n7372 ) | ( n7367 & ~n7372 ) ;
  assign n7374 = ( x96 & n7082 ) | ( x96 & ~n7177 ) | ( n7082 & ~n7177 ) ;
  assign n7375 = x96 & n7082 ;
  assign n7376 = ( ~n7087 & n7374 ) | ( ~n7087 & n7375 ) | ( n7374 & n7375 ) ;
  assign n7377 = ( n7087 & n7374 ) | ( n7087 & n7375 ) | ( n7374 & n7375 ) ;
  assign n7378 = ( n7087 & n7376 ) | ( n7087 & ~n7377 ) | ( n7376 & ~n7377 ) ;
  assign n7379 = ( x97 & n7373 ) | ( x97 & ~n7378 ) | ( n7373 & ~n7378 ) ;
  assign n7380 = ( x97 & n7088 ) | ( x97 & ~n7177 ) | ( n7088 & ~n7177 ) ;
  assign n7381 = x97 & n7088 ;
  assign n7382 = ( ~n7093 & n7380 ) | ( ~n7093 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7383 = ( n7093 & n7380 ) | ( n7093 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7384 = ( n7093 & n7382 ) | ( n7093 & ~n7383 ) | ( n7382 & ~n7383 ) ;
  assign n7385 = ( x98 & n7379 ) | ( x98 & ~n7384 ) | ( n7379 & ~n7384 ) ;
  assign n7386 = ( x98 & n7094 ) | ( x98 & ~n7177 ) | ( n7094 & ~n7177 ) ;
  assign n7387 = x98 & n7094 ;
  assign n7388 = ( ~n7099 & n7386 ) | ( ~n7099 & n7387 ) | ( n7386 & n7387 ) ;
  assign n7389 = ( n7099 & n7386 ) | ( n7099 & n7387 ) | ( n7386 & n7387 ) ;
  assign n7390 = ( n7099 & n7388 ) | ( n7099 & ~n7389 ) | ( n7388 & ~n7389 ) ;
  assign n7391 = ( x99 & n7385 ) | ( x99 & ~n7390 ) | ( n7385 & ~n7390 ) ;
  assign n7392 = ( x99 & n7100 ) | ( x99 & ~n7177 ) | ( n7100 & ~n7177 ) ;
  assign n7393 = x99 & n7100 ;
  assign n7394 = ( ~n7105 & n7392 ) | ( ~n7105 & n7393 ) | ( n7392 & n7393 ) ;
  assign n7395 = ( n7105 & n7392 ) | ( n7105 & n7393 ) | ( n7392 & n7393 ) ;
  assign n7396 = ( n7105 & n7394 ) | ( n7105 & ~n7395 ) | ( n7394 & ~n7395 ) ;
  assign n7397 = ( x100 & n7391 ) | ( x100 & ~n7396 ) | ( n7391 & ~n7396 ) ;
  assign n7398 = ( x100 & n7106 ) | ( x100 & ~n7177 ) | ( n7106 & ~n7177 ) ;
  assign n7399 = x100 & n7106 ;
  assign n7400 = ( ~n7111 & n7398 ) | ( ~n7111 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7401 = ( n7111 & n7398 ) | ( n7111 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7402 = ( n7111 & n7400 ) | ( n7111 & ~n7401 ) | ( n7400 & ~n7401 ) ;
  assign n7403 = ( x101 & n7397 ) | ( x101 & ~n7402 ) | ( n7397 & ~n7402 ) ;
  assign n7404 = ( x101 & n7112 ) | ( x101 & ~n7177 ) | ( n7112 & ~n7177 ) ;
  assign n7405 = x101 & n7112 ;
  assign n7406 = ( ~n7117 & n7404 ) | ( ~n7117 & n7405 ) | ( n7404 & n7405 ) ;
  assign n7407 = ( n7117 & n7404 ) | ( n7117 & n7405 ) | ( n7404 & n7405 ) ;
  assign n7408 = ( n7117 & n7406 ) | ( n7117 & ~n7407 ) | ( n7406 & ~n7407 ) ;
  assign n7409 = ( x102 & n7403 ) | ( x102 & ~n7408 ) | ( n7403 & ~n7408 ) ;
  assign n7410 = ( x102 & n7118 ) | ( x102 & ~n7177 ) | ( n7118 & ~n7177 ) ;
  assign n7411 = x102 & n7118 ;
  assign n7412 = ( ~n7123 & n7410 ) | ( ~n7123 & n7411 ) | ( n7410 & n7411 ) ;
  assign n7413 = ( n7123 & n7410 ) | ( n7123 & n7411 ) | ( n7410 & n7411 ) ;
  assign n7414 = ( n7123 & n7412 ) | ( n7123 & ~n7413 ) | ( n7412 & ~n7413 ) ;
  assign n7415 = ( x103 & n7409 ) | ( x103 & ~n7414 ) | ( n7409 & ~n7414 ) ;
  assign n7416 = ( x103 & n7124 ) | ( x103 & ~n7177 ) | ( n7124 & ~n7177 ) ;
  assign n7417 = x103 & n7124 ;
  assign n7418 = ( ~n7129 & n7416 ) | ( ~n7129 & n7417 ) | ( n7416 & n7417 ) ;
  assign n7419 = ( n7129 & n7416 ) | ( n7129 & n7417 ) | ( n7416 & n7417 ) ;
  assign n7420 = ( n7129 & n7418 ) | ( n7129 & ~n7419 ) | ( n7418 & ~n7419 ) ;
  assign n7421 = ( x104 & n7415 ) | ( x104 & ~n7420 ) | ( n7415 & ~n7420 ) ;
  assign n7422 = ( x104 & n7130 ) | ( x104 & ~n7177 ) | ( n7130 & ~n7177 ) ;
  assign n7423 = x104 & n7130 ;
  assign n7424 = ( ~n7135 & n7422 ) | ( ~n7135 & n7423 ) | ( n7422 & n7423 ) ;
  assign n7425 = ( n7135 & n7422 ) | ( n7135 & n7423 ) | ( n7422 & n7423 ) ;
  assign n7426 = ( n7135 & n7424 ) | ( n7135 & ~n7425 ) | ( n7424 & ~n7425 ) ;
  assign n7427 = ( x105 & n7421 ) | ( x105 & ~n7426 ) | ( n7421 & ~n7426 ) ;
  assign n7428 = ( x105 & n7136 ) | ( x105 & ~n7177 ) | ( n7136 & ~n7177 ) ;
  assign n7429 = x105 & n7136 ;
  assign n7430 = ( ~n7141 & n7428 ) | ( ~n7141 & n7429 ) | ( n7428 & n7429 ) ;
  assign n7431 = ( n7141 & n7428 ) | ( n7141 & n7429 ) | ( n7428 & n7429 ) ;
  assign n7432 = ( n7141 & n7430 ) | ( n7141 & ~n7431 ) | ( n7430 & ~n7431 ) ;
  assign n7433 = ( x106 & n7427 ) | ( x106 & ~n7432 ) | ( n7427 & ~n7432 ) ;
  assign n7434 = ( x106 & n7142 ) | ( x106 & ~n7177 ) | ( n7142 & ~n7177 ) ;
  assign n7435 = x106 & n7142 ;
  assign n7436 = ( ~n7147 & n7434 ) | ( ~n7147 & n7435 ) | ( n7434 & n7435 ) ;
  assign n7437 = ( n7147 & n7434 ) | ( n7147 & n7435 ) | ( n7434 & n7435 ) ;
  assign n7438 = ( n7147 & n7436 ) | ( n7147 & ~n7437 ) | ( n7436 & ~n7437 ) ;
  assign n7439 = ( x107 & n7433 ) | ( x107 & ~n7438 ) | ( n7433 & ~n7438 ) ;
  assign n7440 = ( x107 & n7148 ) | ( x107 & ~n7177 ) | ( n7148 & ~n7177 ) ;
  assign n7441 = x107 & n7148 ;
  assign n7442 = ( ~n7153 & n7440 ) | ( ~n7153 & n7441 ) | ( n7440 & n7441 ) ;
  assign n7443 = ( n7153 & n7440 ) | ( n7153 & n7441 ) | ( n7440 & n7441 ) ;
  assign n7444 = ( n7153 & n7442 ) | ( n7153 & ~n7443 ) | ( n7442 & ~n7443 ) ;
  assign n7445 = ( x108 & n7439 ) | ( x108 & ~n7444 ) | ( n7439 & ~n7444 ) ;
  assign n7446 = ( x108 & n7154 ) | ( x108 & ~n7177 ) | ( n7154 & ~n7177 ) ;
  assign n7447 = x108 & n7154 ;
  assign n7448 = ( ~n7159 & n7446 ) | ( ~n7159 & n7447 ) | ( n7446 & n7447 ) ;
  assign n7449 = ( n7159 & n7446 ) | ( n7159 & n7447 ) | ( n7446 & n7447 ) ;
  assign n7450 = ( n7159 & n7448 ) | ( n7159 & ~n7449 ) | ( n7448 & ~n7449 ) ;
  assign n7451 = ( x109 & n7445 ) | ( x109 & ~n7450 ) | ( n7445 & ~n7450 ) ;
  assign n7452 = ( x109 & n7160 ) | ( x109 & ~n7177 ) | ( n7160 & ~n7177 ) ;
  assign n7453 = x109 & n7160 ;
  assign n7454 = ( ~n7165 & n7452 ) | ( ~n7165 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7455 = ( n7165 & n7452 ) | ( n7165 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7456 = ( n7165 & n7454 ) | ( n7165 & ~n7455 ) | ( n7454 & ~n7455 ) ;
  assign n7457 = ( x110 & n7451 ) | ( x110 & ~n7456 ) | ( n7451 & ~n7456 ) ;
  assign n7458 = ( x110 & n7166 ) | ( x110 & ~n7177 ) | ( n7166 & ~n7177 ) ;
  assign n7459 = x110 & n7166 ;
  assign n7460 = ( ~n7171 & n7458 ) | ( ~n7171 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7461 = ( n7171 & n7458 ) | ( n7171 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7462 = ( n7171 & n7460 ) | ( n7171 & ~n7461 ) | ( n7460 & ~n7461 ) ;
  assign n7463 = ( x111 & n7457 ) | ( x111 & ~n7462 ) | ( n7457 & ~n7462 ) ;
  assign n7464 = ( x112 & ~n7182 ) | ( x112 & n7463 ) | ( ~n7182 & n7463 ) ;
  assign n7465 = ( n143 & n144 ) | ( n143 & ~n6888 ) | ( n144 & ~n6888 ) ;
  assign n7466 = ( ~x112 & n7174 ) | ( ~x112 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7467 = ( ~x112 & n144 ) | ( ~x112 & n7175 ) | ( n144 & n7175 ) ;
  assign n7468 = ( n7465 & n7466 ) | ( n7465 & n7467 ) | ( n7466 & n7467 ) ;
  assign n7469 = n7466 & ~n7468 ;
  assign n7470 = ( n7464 & n7465 ) | ( n7464 & ~n7469 ) | ( n7465 & ~n7469 ) ;
  assign n7471 = ( x112 & n7463 ) | ( x112 & n7470 ) | ( n7463 & n7470 ) ;
  assign n7472 = x112 | n7463 ;
  assign n7473 = ( ~n7182 & n7471 ) | ( ~n7182 & n7472 ) | ( n7471 & n7472 ) ;
  assign n7474 = ( n7182 & n7471 ) | ( n7182 & n7472 ) | ( n7471 & n7472 ) ;
  assign n7475 = ( n7182 & n7473 ) | ( n7182 & ~n7474 ) | ( n7473 & ~n7474 ) ;
  assign n7476 = ~x13 & x64 ;
  assign n7477 = ~x14 & n7470 ;
  assign n7478 = ( x14 & ~x64 ) | ( x14 & n7470 ) | ( ~x64 & n7470 ) ;
  assign n7479 = ( n7183 & ~n7477 ) | ( n7183 & n7478 ) | ( ~n7477 & n7478 ) ;
  assign n7480 = ( x65 & n7476 ) | ( x65 & ~n7479 ) | ( n7476 & ~n7479 ) ;
  assign n7481 = ( x65 & n7183 ) | ( x65 & n7470 ) | ( n7183 & n7470 ) ;
  assign n7482 = x65 | n7183 ;
  assign n7483 = ( ~n7186 & n7481 ) | ( ~n7186 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7484 = ( n7186 & n7481 ) | ( n7186 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7485 = ( n7186 & n7483 ) | ( n7186 & ~n7484 ) | ( n7483 & ~n7484 ) ;
  assign n7486 = ( x66 & n7480 ) | ( x66 & ~n7485 ) | ( n7480 & ~n7485 ) ;
  assign n7487 = ( x66 & n7187 ) | ( x66 & n7470 ) | ( n7187 & n7470 ) ;
  assign n7488 = x66 | n7187 ;
  assign n7489 = ( ~n7192 & n7487 ) | ( ~n7192 & n7488 ) | ( n7487 & n7488 ) ;
  assign n7490 = ( n7192 & n7487 ) | ( n7192 & n7488 ) | ( n7487 & n7488 ) ;
  assign n7491 = ( n7192 & n7489 ) | ( n7192 & ~n7490 ) | ( n7489 & ~n7490 ) ;
  assign n7492 = ( x67 & n7486 ) | ( x67 & ~n7491 ) | ( n7486 & ~n7491 ) ;
  assign n7493 = ( x67 & n7193 ) | ( x67 & ~n7470 ) | ( n7193 & ~n7470 ) ;
  assign n7494 = x67 & n7193 ;
  assign n7495 = ( ~n7198 & n7493 ) | ( ~n7198 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7496 = ( n7198 & n7493 ) | ( n7198 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7497 = ( n7198 & n7495 ) | ( n7198 & ~n7496 ) | ( n7495 & ~n7496 ) ;
  assign n7498 = ( x68 & n7492 ) | ( x68 & ~n7497 ) | ( n7492 & ~n7497 ) ;
  assign n7499 = ( x68 & n7199 ) | ( x68 & ~n7470 ) | ( n7199 & ~n7470 ) ;
  assign n7500 = x68 & n7199 ;
  assign n7501 = ( ~n7204 & n7499 ) | ( ~n7204 & n7500 ) | ( n7499 & n7500 ) ;
  assign n7502 = ( n7204 & n7499 ) | ( n7204 & n7500 ) | ( n7499 & n7500 ) ;
  assign n7503 = ( n7204 & n7501 ) | ( n7204 & ~n7502 ) | ( n7501 & ~n7502 ) ;
  assign n7504 = ( x69 & n7498 ) | ( x69 & ~n7503 ) | ( n7498 & ~n7503 ) ;
  assign n7505 = ( x69 & n7205 ) | ( x69 & ~n7470 ) | ( n7205 & ~n7470 ) ;
  assign n7506 = x69 & n7205 ;
  assign n7507 = ( ~n7210 & n7505 ) | ( ~n7210 & n7506 ) | ( n7505 & n7506 ) ;
  assign n7508 = ( n7210 & n7505 ) | ( n7210 & n7506 ) | ( n7505 & n7506 ) ;
  assign n7509 = ( n7210 & n7507 ) | ( n7210 & ~n7508 ) | ( n7507 & ~n7508 ) ;
  assign n7510 = ( x70 & n7504 ) | ( x70 & ~n7509 ) | ( n7504 & ~n7509 ) ;
  assign n7511 = ( x70 & n7211 ) | ( x70 & ~n7470 ) | ( n7211 & ~n7470 ) ;
  assign n7512 = x70 & n7211 ;
  assign n7513 = ( ~n7216 & n7511 ) | ( ~n7216 & n7512 ) | ( n7511 & n7512 ) ;
  assign n7514 = ( n7216 & n7511 ) | ( n7216 & n7512 ) | ( n7511 & n7512 ) ;
  assign n7515 = ( n7216 & n7513 ) | ( n7216 & ~n7514 ) | ( n7513 & ~n7514 ) ;
  assign n7516 = ( x71 & n7510 ) | ( x71 & ~n7515 ) | ( n7510 & ~n7515 ) ;
  assign n7517 = ( x71 & n7217 ) | ( x71 & ~n7470 ) | ( n7217 & ~n7470 ) ;
  assign n7518 = x71 & n7217 ;
  assign n7519 = ( ~n7222 & n7517 ) | ( ~n7222 & n7518 ) | ( n7517 & n7518 ) ;
  assign n7520 = ( n7222 & n7517 ) | ( n7222 & n7518 ) | ( n7517 & n7518 ) ;
  assign n7521 = ( n7222 & n7519 ) | ( n7222 & ~n7520 ) | ( n7519 & ~n7520 ) ;
  assign n7522 = ( x72 & n7516 ) | ( x72 & ~n7521 ) | ( n7516 & ~n7521 ) ;
  assign n7523 = ( x72 & n7223 ) | ( x72 & ~n7470 ) | ( n7223 & ~n7470 ) ;
  assign n7524 = x72 & n7223 ;
  assign n7525 = ( ~n7228 & n7523 ) | ( ~n7228 & n7524 ) | ( n7523 & n7524 ) ;
  assign n7526 = ( n7228 & n7523 ) | ( n7228 & n7524 ) | ( n7523 & n7524 ) ;
  assign n7527 = ( n7228 & n7525 ) | ( n7228 & ~n7526 ) | ( n7525 & ~n7526 ) ;
  assign n7528 = ( x73 & n7522 ) | ( x73 & ~n7527 ) | ( n7522 & ~n7527 ) ;
  assign n7529 = ( x73 & n7229 ) | ( x73 & ~n7470 ) | ( n7229 & ~n7470 ) ;
  assign n7530 = x73 & n7229 ;
  assign n7531 = ( ~n7234 & n7529 ) | ( ~n7234 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7532 = ( n7234 & n7529 ) | ( n7234 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7533 = ( n7234 & n7531 ) | ( n7234 & ~n7532 ) | ( n7531 & ~n7532 ) ;
  assign n7534 = ( x74 & n7528 ) | ( x74 & ~n7533 ) | ( n7528 & ~n7533 ) ;
  assign n7535 = ( x74 & n7235 ) | ( x74 & ~n7470 ) | ( n7235 & ~n7470 ) ;
  assign n7536 = x74 & n7235 ;
  assign n7537 = ( ~n7240 & n7535 ) | ( ~n7240 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7538 = ( n7240 & n7535 ) | ( n7240 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7539 = ( n7240 & n7537 ) | ( n7240 & ~n7538 ) | ( n7537 & ~n7538 ) ;
  assign n7540 = ( x75 & n7534 ) | ( x75 & ~n7539 ) | ( n7534 & ~n7539 ) ;
  assign n7541 = ( x75 & n7241 ) | ( x75 & ~n7470 ) | ( n7241 & ~n7470 ) ;
  assign n7542 = x75 & n7241 ;
  assign n7543 = ( ~n7246 & n7541 ) | ( ~n7246 & n7542 ) | ( n7541 & n7542 ) ;
  assign n7544 = ( n7246 & n7541 ) | ( n7246 & n7542 ) | ( n7541 & n7542 ) ;
  assign n7545 = ( n7246 & n7543 ) | ( n7246 & ~n7544 ) | ( n7543 & ~n7544 ) ;
  assign n7546 = ( x76 & n7540 ) | ( x76 & ~n7545 ) | ( n7540 & ~n7545 ) ;
  assign n7547 = ( x76 & n7247 ) | ( x76 & ~n7470 ) | ( n7247 & ~n7470 ) ;
  assign n7548 = x76 & n7247 ;
  assign n7549 = ( ~n7252 & n7547 ) | ( ~n7252 & n7548 ) | ( n7547 & n7548 ) ;
  assign n7550 = ( n7252 & n7547 ) | ( n7252 & n7548 ) | ( n7547 & n7548 ) ;
  assign n7551 = ( n7252 & n7549 ) | ( n7252 & ~n7550 ) | ( n7549 & ~n7550 ) ;
  assign n7552 = ( x77 & n7546 ) | ( x77 & ~n7551 ) | ( n7546 & ~n7551 ) ;
  assign n7553 = ( x77 & n7253 ) | ( x77 & ~n7470 ) | ( n7253 & ~n7470 ) ;
  assign n7554 = x77 & n7253 ;
  assign n7555 = ( ~n7258 & n7553 ) | ( ~n7258 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7556 = ( n7258 & n7553 ) | ( n7258 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7557 = ( n7258 & n7555 ) | ( n7258 & ~n7556 ) | ( n7555 & ~n7556 ) ;
  assign n7558 = ( x78 & n7552 ) | ( x78 & ~n7557 ) | ( n7552 & ~n7557 ) ;
  assign n7559 = ( x78 & n7259 ) | ( x78 & ~n7470 ) | ( n7259 & ~n7470 ) ;
  assign n7560 = x78 & n7259 ;
  assign n7561 = ( ~n7264 & n7559 ) | ( ~n7264 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7562 = ( n7264 & n7559 ) | ( n7264 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7563 = ( n7264 & n7561 ) | ( n7264 & ~n7562 ) | ( n7561 & ~n7562 ) ;
  assign n7564 = ( x79 & n7558 ) | ( x79 & ~n7563 ) | ( n7558 & ~n7563 ) ;
  assign n7565 = ( x79 & n7265 ) | ( x79 & ~n7470 ) | ( n7265 & ~n7470 ) ;
  assign n7566 = x79 & n7265 ;
  assign n7567 = ( ~n7270 & n7565 ) | ( ~n7270 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7568 = ( n7270 & n7565 ) | ( n7270 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7569 = ( n7270 & n7567 ) | ( n7270 & ~n7568 ) | ( n7567 & ~n7568 ) ;
  assign n7570 = ( x80 & n7564 ) | ( x80 & ~n7569 ) | ( n7564 & ~n7569 ) ;
  assign n7571 = ( x80 & n7271 ) | ( x80 & ~n7470 ) | ( n7271 & ~n7470 ) ;
  assign n7572 = x80 & n7271 ;
  assign n7573 = ( ~n7276 & n7571 ) | ( ~n7276 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = ( n7276 & n7571 ) | ( n7276 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7575 = ( n7276 & n7573 ) | ( n7276 & ~n7574 ) | ( n7573 & ~n7574 ) ;
  assign n7576 = ( x81 & n7570 ) | ( x81 & ~n7575 ) | ( n7570 & ~n7575 ) ;
  assign n7577 = ( x81 & n7277 ) | ( x81 & ~n7470 ) | ( n7277 & ~n7470 ) ;
  assign n7578 = x81 & n7277 ;
  assign n7579 = ( ~n7282 & n7577 ) | ( ~n7282 & n7578 ) | ( n7577 & n7578 ) ;
  assign n7580 = ( n7282 & n7577 ) | ( n7282 & n7578 ) | ( n7577 & n7578 ) ;
  assign n7581 = ( n7282 & n7579 ) | ( n7282 & ~n7580 ) | ( n7579 & ~n7580 ) ;
  assign n7582 = ( x82 & n7576 ) | ( x82 & ~n7581 ) | ( n7576 & ~n7581 ) ;
  assign n7583 = ( x82 & n7283 ) | ( x82 & ~n7470 ) | ( n7283 & ~n7470 ) ;
  assign n7584 = x82 & n7283 ;
  assign n7585 = ( ~n7288 & n7583 ) | ( ~n7288 & n7584 ) | ( n7583 & n7584 ) ;
  assign n7586 = ( n7288 & n7583 ) | ( n7288 & n7584 ) | ( n7583 & n7584 ) ;
  assign n7587 = ( n7288 & n7585 ) | ( n7288 & ~n7586 ) | ( n7585 & ~n7586 ) ;
  assign n7588 = ( x83 & n7582 ) | ( x83 & ~n7587 ) | ( n7582 & ~n7587 ) ;
  assign n7589 = ( x83 & n7289 ) | ( x83 & ~n7470 ) | ( n7289 & ~n7470 ) ;
  assign n7590 = x83 & n7289 ;
  assign n7591 = ( ~n7294 & n7589 ) | ( ~n7294 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7592 = ( n7294 & n7589 ) | ( n7294 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7593 = ( n7294 & n7591 ) | ( n7294 & ~n7592 ) | ( n7591 & ~n7592 ) ;
  assign n7594 = ( x84 & n7588 ) | ( x84 & ~n7593 ) | ( n7588 & ~n7593 ) ;
  assign n7595 = ( x84 & n7295 ) | ( x84 & ~n7470 ) | ( n7295 & ~n7470 ) ;
  assign n7596 = x84 & n7295 ;
  assign n7597 = ( ~n7300 & n7595 ) | ( ~n7300 & n7596 ) | ( n7595 & n7596 ) ;
  assign n7598 = ( n7300 & n7595 ) | ( n7300 & n7596 ) | ( n7595 & n7596 ) ;
  assign n7599 = ( n7300 & n7597 ) | ( n7300 & ~n7598 ) | ( n7597 & ~n7598 ) ;
  assign n7600 = ( x85 & n7594 ) | ( x85 & ~n7599 ) | ( n7594 & ~n7599 ) ;
  assign n7601 = ( x85 & n7301 ) | ( x85 & ~n7470 ) | ( n7301 & ~n7470 ) ;
  assign n7602 = x85 & n7301 ;
  assign n7603 = ( ~n7306 & n7601 ) | ( ~n7306 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7604 = ( n7306 & n7601 ) | ( n7306 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7605 = ( n7306 & n7603 ) | ( n7306 & ~n7604 ) | ( n7603 & ~n7604 ) ;
  assign n7606 = ( x86 & n7600 ) | ( x86 & ~n7605 ) | ( n7600 & ~n7605 ) ;
  assign n7607 = ( x86 & n7307 ) | ( x86 & ~n7470 ) | ( n7307 & ~n7470 ) ;
  assign n7608 = x86 & n7307 ;
  assign n7609 = ( ~n7312 & n7607 ) | ( ~n7312 & n7608 ) | ( n7607 & n7608 ) ;
  assign n7610 = ( n7312 & n7607 ) | ( n7312 & n7608 ) | ( n7607 & n7608 ) ;
  assign n7611 = ( n7312 & n7609 ) | ( n7312 & ~n7610 ) | ( n7609 & ~n7610 ) ;
  assign n7612 = ( x87 & n7606 ) | ( x87 & ~n7611 ) | ( n7606 & ~n7611 ) ;
  assign n7613 = ( x87 & n7313 ) | ( x87 & ~n7470 ) | ( n7313 & ~n7470 ) ;
  assign n7614 = x87 & n7313 ;
  assign n7615 = ( ~n7318 & n7613 ) | ( ~n7318 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7616 = ( n7318 & n7613 ) | ( n7318 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7617 = ( n7318 & n7615 ) | ( n7318 & ~n7616 ) | ( n7615 & ~n7616 ) ;
  assign n7618 = ( x88 & n7612 ) | ( x88 & ~n7617 ) | ( n7612 & ~n7617 ) ;
  assign n7619 = ( x88 & n7319 ) | ( x88 & ~n7470 ) | ( n7319 & ~n7470 ) ;
  assign n7620 = x88 & n7319 ;
  assign n7621 = ( ~n7324 & n7619 ) | ( ~n7324 & n7620 ) | ( n7619 & n7620 ) ;
  assign n7622 = ( n7324 & n7619 ) | ( n7324 & n7620 ) | ( n7619 & n7620 ) ;
  assign n7623 = ( n7324 & n7621 ) | ( n7324 & ~n7622 ) | ( n7621 & ~n7622 ) ;
  assign n7624 = ( x89 & n7618 ) | ( x89 & ~n7623 ) | ( n7618 & ~n7623 ) ;
  assign n7625 = ( x89 & n7325 ) | ( x89 & ~n7470 ) | ( n7325 & ~n7470 ) ;
  assign n7626 = x89 & n7325 ;
  assign n7627 = ( ~n7330 & n7625 ) | ( ~n7330 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7628 = ( n7330 & n7625 ) | ( n7330 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7629 = ( n7330 & n7627 ) | ( n7330 & ~n7628 ) | ( n7627 & ~n7628 ) ;
  assign n7630 = ( x90 & n7624 ) | ( x90 & ~n7629 ) | ( n7624 & ~n7629 ) ;
  assign n7631 = ( x90 & n7331 ) | ( x90 & ~n7470 ) | ( n7331 & ~n7470 ) ;
  assign n7632 = x90 & n7331 ;
  assign n7633 = ( ~n7336 & n7631 ) | ( ~n7336 & n7632 ) | ( n7631 & n7632 ) ;
  assign n7634 = ( n7336 & n7631 ) | ( n7336 & n7632 ) | ( n7631 & n7632 ) ;
  assign n7635 = ( n7336 & n7633 ) | ( n7336 & ~n7634 ) | ( n7633 & ~n7634 ) ;
  assign n7636 = ( x91 & n7630 ) | ( x91 & ~n7635 ) | ( n7630 & ~n7635 ) ;
  assign n7637 = ( x91 & n7337 ) | ( x91 & ~n7470 ) | ( n7337 & ~n7470 ) ;
  assign n7638 = x91 & n7337 ;
  assign n7639 = ( ~n7342 & n7637 ) | ( ~n7342 & n7638 ) | ( n7637 & n7638 ) ;
  assign n7640 = ( n7342 & n7637 ) | ( n7342 & n7638 ) | ( n7637 & n7638 ) ;
  assign n7641 = ( n7342 & n7639 ) | ( n7342 & ~n7640 ) | ( n7639 & ~n7640 ) ;
  assign n7642 = ( x92 & n7636 ) | ( x92 & ~n7641 ) | ( n7636 & ~n7641 ) ;
  assign n7643 = ( x92 & n7343 ) | ( x92 & ~n7470 ) | ( n7343 & ~n7470 ) ;
  assign n7644 = x92 & n7343 ;
  assign n7645 = ( ~n7348 & n7643 ) | ( ~n7348 & n7644 ) | ( n7643 & n7644 ) ;
  assign n7646 = ( n7348 & n7643 ) | ( n7348 & n7644 ) | ( n7643 & n7644 ) ;
  assign n7647 = ( n7348 & n7645 ) | ( n7348 & ~n7646 ) | ( n7645 & ~n7646 ) ;
  assign n7648 = ( x93 & n7642 ) | ( x93 & ~n7647 ) | ( n7642 & ~n7647 ) ;
  assign n7649 = ( x93 & n7349 ) | ( x93 & ~n7470 ) | ( n7349 & ~n7470 ) ;
  assign n7650 = x93 & n7349 ;
  assign n7651 = ( ~n7354 & n7649 ) | ( ~n7354 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7652 = ( n7354 & n7649 ) | ( n7354 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7653 = ( n7354 & n7651 ) | ( n7354 & ~n7652 ) | ( n7651 & ~n7652 ) ;
  assign n7654 = ( x94 & n7648 ) | ( x94 & ~n7653 ) | ( n7648 & ~n7653 ) ;
  assign n7655 = ( x94 & n7355 ) | ( x94 & ~n7470 ) | ( n7355 & ~n7470 ) ;
  assign n7656 = x94 & n7355 ;
  assign n7657 = ( ~n7360 & n7655 ) | ( ~n7360 & n7656 ) | ( n7655 & n7656 ) ;
  assign n7658 = ( n7360 & n7655 ) | ( n7360 & n7656 ) | ( n7655 & n7656 ) ;
  assign n7659 = ( n7360 & n7657 ) | ( n7360 & ~n7658 ) | ( n7657 & ~n7658 ) ;
  assign n7660 = ( x95 & n7654 ) | ( x95 & ~n7659 ) | ( n7654 & ~n7659 ) ;
  assign n7661 = ( x95 & n7361 ) | ( x95 & ~n7470 ) | ( n7361 & ~n7470 ) ;
  assign n7662 = x95 & n7361 ;
  assign n7663 = ( ~n7366 & n7661 ) | ( ~n7366 & n7662 ) | ( n7661 & n7662 ) ;
  assign n7664 = ( n7366 & n7661 ) | ( n7366 & n7662 ) | ( n7661 & n7662 ) ;
  assign n7665 = ( n7366 & n7663 ) | ( n7366 & ~n7664 ) | ( n7663 & ~n7664 ) ;
  assign n7666 = ( x96 & n7660 ) | ( x96 & ~n7665 ) | ( n7660 & ~n7665 ) ;
  assign n7667 = ( x96 & n7367 ) | ( x96 & ~n7470 ) | ( n7367 & ~n7470 ) ;
  assign n7668 = x96 & n7367 ;
  assign n7669 = ( ~n7372 & n7667 ) | ( ~n7372 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7670 = ( n7372 & n7667 ) | ( n7372 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7671 = ( n7372 & n7669 ) | ( n7372 & ~n7670 ) | ( n7669 & ~n7670 ) ;
  assign n7672 = ( x97 & n7666 ) | ( x97 & ~n7671 ) | ( n7666 & ~n7671 ) ;
  assign n7673 = ( x97 & n7373 ) | ( x97 & ~n7470 ) | ( n7373 & ~n7470 ) ;
  assign n7674 = x97 & n7373 ;
  assign n7675 = ( ~n7378 & n7673 ) | ( ~n7378 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7676 = ( n7378 & n7673 ) | ( n7378 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7677 = ( n7378 & n7675 ) | ( n7378 & ~n7676 ) | ( n7675 & ~n7676 ) ;
  assign n7678 = ( x98 & n7672 ) | ( x98 & ~n7677 ) | ( n7672 & ~n7677 ) ;
  assign n7679 = ( x98 & n7379 ) | ( x98 & ~n7470 ) | ( n7379 & ~n7470 ) ;
  assign n7680 = x98 & n7379 ;
  assign n7681 = ( ~n7384 & n7679 ) | ( ~n7384 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7682 = ( n7384 & n7679 ) | ( n7384 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7683 = ( n7384 & n7681 ) | ( n7384 & ~n7682 ) | ( n7681 & ~n7682 ) ;
  assign n7684 = ( x99 & n7678 ) | ( x99 & ~n7683 ) | ( n7678 & ~n7683 ) ;
  assign n7685 = ( x99 & n7385 ) | ( x99 & ~n7470 ) | ( n7385 & ~n7470 ) ;
  assign n7686 = x99 & n7385 ;
  assign n7687 = ( ~n7390 & n7685 ) | ( ~n7390 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7688 = ( n7390 & n7685 ) | ( n7390 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7689 = ( n7390 & n7687 ) | ( n7390 & ~n7688 ) | ( n7687 & ~n7688 ) ;
  assign n7690 = ( x100 & n7684 ) | ( x100 & ~n7689 ) | ( n7684 & ~n7689 ) ;
  assign n7691 = ( x100 & n7391 ) | ( x100 & ~n7470 ) | ( n7391 & ~n7470 ) ;
  assign n7692 = x100 & n7391 ;
  assign n7693 = ( ~n7396 & n7691 ) | ( ~n7396 & n7692 ) | ( n7691 & n7692 ) ;
  assign n7694 = ( n7396 & n7691 ) | ( n7396 & n7692 ) | ( n7691 & n7692 ) ;
  assign n7695 = ( n7396 & n7693 ) | ( n7396 & ~n7694 ) | ( n7693 & ~n7694 ) ;
  assign n7696 = ( x101 & n7690 ) | ( x101 & ~n7695 ) | ( n7690 & ~n7695 ) ;
  assign n7697 = ( x101 & n7397 ) | ( x101 & ~n7470 ) | ( n7397 & ~n7470 ) ;
  assign n7698 = x101 & n7397 ;
  assign n7699 = ( ~n7402 & n7697 ) | ( ~n7402 & n7698 ) | ( n7697 & n7698 ) ;
  assign n7700 = ( n7402 & n7697 ) | ( n7402 & n7698 ) | ( n7697 & n7698 ) ;
  assign n7701 = ( n7402 & n7699 ) | ( n7402 & ~n7700 ) | ( n7699 & ~n7700 ) ;
  assign n7702 = ( x102 & n7696 ) | ( x102 & ~n7701 ) | ( n7696 & ~n7701 ) ;
  assign n7703 = ( x102 & n7403 ) | ( x102 & ~n7470 ) | ( n7403 & ~n7470 ) ;
  assign n7704 = x102 & n7403 ;
  assign n7705 = ( ~n7408 & n7703 ) | ( ~n7408 & n7704 ) | ( n7703 & n7704 ) ;
  assign n7706 = ( n7408 & n7703 ) | ( n7408 & n7704 ) | ( n7703 & n7704 ) ;
  assign n7707 = ( n7408 & n7705 ) | ( n7408 & ~n7706 ) | ( n7705 & ~n7706 ) ;
  assign n7708 = ( x103 & n7702 ) | ( x103 & ~n7707 ) | ( n7702 & ~n7707 ) ;
  assign n7709 = ( x103 & n7409 ) | ( x103 & ~n7470 ) | ( n7409 & ~n7470 ) ;
  assign n7710 = x103 & n7409 ;
  assign n7711 = ( ~n7414 & n7709 ) | ( ~n7414 & n7710 ) | ( n7709 & n7710 ) ;
  assign n7712 = ( n7414 & n7709 ) | ( n7414 & n7710 ) | ( n7709 & n7710 ) ;
  assign n7713 = ( n7414 & n7711 ) | ( n7414 & ~n7712 ) | ( n7711 & ~n7712 ) ;
  assign n7714 = ( x104 & n7708 ) | ( x104 & ~n7713 ) | ( n7708 & ~n7713 ) ;
  assign n7715 = ( x104 & n7415 ) | ( x104 & ~n7470 ) | ( n7415 & ~n7470 ) ;
  assign n7716 = x104 & n7415 ;
  assign n7717 = ( ~n7420 & n7715 ) | ( ~n7420 & n7716 ) | ( n7715 & n7716 ) ;
  assign n7718 = ( n7420 & n7715 ) | ( n7420 & n7716 ) | ( n7715 & n7716 ) ;
  assign n7719 = ( n7420 & n7717 ) | ( n7420 & ~n7718 ) | ( n7717 & ~n7718 ) ;
  assign n7720 = ( x105 & n7714 ) | ( x105 & ~n7719 ) | ( n7714 & ~n7719 ) ;
  assign n7721 = ( x105 & n7421 ) | ( x105 & ~n7470 ) | ( n7421 & ~n7470 ) ;
  assign n7722 = x105 & n7421 ;
  assign n7723 = ( ~n7426 & n7721 ) | ( ~n7426 & n7722 ) | ( n7721 & n7722 ) ;
  assign n7724 = ( n7426 & n7721 ) | ( n7426 & n7722 ) | ( n7721 & n7722 ) ;
  assign n7725 = ( n7426 & n7723 ) | ( n7426 & ~n7724 ) | ( n7723 & ~n7724 ) ;
  assign n7726 = ( x106 & n7720 ) | ( x106 & ~n7725 ) | ( n7720 & ~n7725 ) ;
  assign n7727 = ( x106 & n7427 ) | ( x106 & ~n7470 ) | ( n7427 & ~n7470 ) ;
  assign n7728 = x106 & n7427 ;
  assign n7729 = ( ~n7432 & n7727 ) | ( ~n7432 & n7728 ) | ( n7727 & n7728 ) ;
  assign n7730 = ( n7432 & n7727 ) | ( n7432 & n7728 ) | ( n7727 & n7728 ) ;
  assign n7731 = ( n7432 & n7729 ) | ( n7432 & ~n7730 ) | ( n7729 & ~n7730 ) ;
  assign n7732 = ( x107 & n7726 ) | ( x107 & ~n7731 ) | ( n7726 & ~n7731 ) ;
  assign n7733 = ( x107 & n7433 ) | ( x107 & ~n7470 ) | ( n7433 & ~n7470 ) ;
  assign n7734 = x107 & n7433 ;
  assign n7735 = ( ~n7438 & n7733 ) | ( ~n7438 & n7734 ) | ( n7733 & n7734 ) ;
  assign n7736 = ( n7438 & n7733 ) | ( n7438 & n7734 ) | ( n7733 & n7734 ) ;
  assign n7737 = ( n7438 & n7735 ) | ( n7438 & ~n7736 ) | ( n7735 & ~n7736 ) ;
  assign n7738 = ( x108 & n7732 ) | ( x108 & ~n7737 ) | ( n7732 & ~n7737 ) ;
  assign n7739 = ( x108 & n7439 ) | ( x108 & ~n7470 ) | ( n7439 & ~n7470 ) ;
  assign n7740 = x108 & n7439 ;
  assign n7741 = ( ~n7444 & n7739 ) | ( ~n7444 & n7740 ) | ( n7739 & n7740 ) ;
  assign n7742 = ( n7444 & n7739 ) | ( n7444 & n7740 ) | ( n7739 & n7740 ) ;
  assign n7743 = ( n7444 & n7741 ) | ( n7444 & ~n7742 ) | ( n7741 & ~n7742 ) ;
  assign n7744 = ( x109 & n7738 ) | ( x109 & ~n7743 ) | ( n7738 & ~n7743 ) ;
  assign n7745 = ( x109 & n7445 ) | ( x109 & ~n7470 ) | ( n7445 & ~n7470 ) ;
  assign n7746 = x109 & n7445 ;
  assign n7747 = ( ~n7450 & n7745 ) | ( ~n7450 & n7746 ) | ( n7745 & n7746 ) ;
  assign n7748 = ( n7450 & n7745 ) | ( n7450 & n7746 ) | ( n7745 & n7746 ) ;
  assign n7749 = ( n7450 & n7747 ) | ( n7450 & ~n7748 ) | ( n7747 & ~n7748 ) ;
  assign n7750 = ( x110 & n7744 ) | ( x110 & ~n7749 ) | ( n7744 & ~n7749 ) ;
  assign n7751 = ( x110 & n7451 ) | ( x110 & ~n7470 ) | ( n7451 & ~n7470 ) ;
  assign n7752 = x110 & n7451 ;
  assign n7753 = ( ~n7456 & n7751 ) | ( ~n7456 & n7752 ) | ( n7751 & n7752 ) ;
  assign n7754 = ( n7456 & n7751 ) | ( n7456 & n7752 ) | ( n7751 & n7752 ) ;
  assign n7755 = ( n7456 & n7753 ) | ( n7456 & ~n7754 ) | ( n7753 & ~n7754 ) ;
  assign n7756 = ( x111 & n7750 ) | ( x111 & ~n7755 ) | ( n7750 & ~n7755 ) ;
  assign n7757 = ( x111 & n7457 ) | ( x111 & ~n7470 ) | ( n7457 & ~n7470 ) ;
  assign n7758 = x111 & n7457 ;
  assign n7759 = ( ~n7462 & n7757 ) | ( ~n7462 & n7758 ) | ( n7757 & n7758 ) ;
  assign n7760 = ( n7462 & n7757 ) | ( n7462 & n7758 ) | ( n7757 & n7758 ) ;
  assign n7761 = ( n7462 & n7759 ) | ( n7462 & ~n7760 ) | ( n7759 & ~n7760 ) ;
  assign n7762 = ( x112 & n7756 ) | ( x112 & ~n7761 ) | ( n7756 & ~n7761 ) ;
  assign n7763 = ( x113 & ~n7475 ) | ( x113 & n7762 ) | ( ~n7475 & n7762 ) ;
  assign n7764 = ( n143 & n144 ) | ( n143 & n7464 ) | ( n144 & n7464 ) ;
  assign n7765 = ( n389 & n6888 ) | ( n389 & n7764 ) | ( n6888 & n7764 ) ;
  assign n7766 = ( x114 & n7763 ) | ( x114 & ~n7765 ) | ( n7763 & ~n7765 ) ;
  assign n7767 = n142 | n7766 ;
  assign n7768 = ( x113 & n7762 ) | ( x113 & n7767 ) | ( n7762 & n7767 ) ;
  assign n7769 = x113 | n7762 ;
  assign n7770 = ( ~n7475 & n7768 ) | ( ~n7475 & n7769 ) | ( n7768 & n7769 ) ;
  assign n7771 = ( n7475 & n7768 ) | ( n7475 & n7769 ) | ( n7768 & n7769 ) ;
  assign n7772 = ( n7475 & n7770 ) | ( n7475 & ~n7771 ) | ( n7770 & ~n7771 ) ;
  assign n7773 = ~x12 & x64 ;
  assign n7774 = ~x13 & n7767 ;
  assign n7775 = ( x13 & ~x64 ) | ( x13 & n7767 ) | ( ~x64 & n7767 ) ;
  assign n7776 = ( n7476 & ~n7774 ) | ( n7476 & n7775 ) | ( ~n7774 & n7775 ) ;
  assign n7777 = ( x65 & n7773 ) | ( x65 & ~n7776 ) | ( n7773 & ~n7776 ) ;
  assign n7778 = ( x65 & n7476 ) | ( x65 & n7767 ) | ( n7476 & n7767 ) ;
  assign n7779 = x65 | n7476 ;
  assign n7780 = ( ~n7479 & n7778 ) | ( ~n7479 & n7779 ) | ( n7778 & n7779 ) ;
  assign n7781 = ( n7479 & n7778 ) | ( n7479 & n7779 ) | ( n7778 & n7779 ) ;
  assign n7782 = ( n7479 & n7780 ) | ( n7479 & ~n7781 ) | ( n7780 & ~n7781 ) ;
  assign n7783 = ( x66 & n7777 ) | ( x66 & ~n7782 ) | ( n7777 & ~n7782 ) ;
  assign n7784 = ( x66 & n7480 ) | ( x66 & n7767 ) | ( n7480 & n7767 ) ;
  assign n7785 = x66 | n7480 ;
  assign n7786 = ( ~n7485 & n7784 ) | ( ~n7485 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7787 = ( n7485 & n7784 ) | ( n7485 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7788 = ( n7485 & n7786 ) | ( n7485 & ~n7787 ) | ( n7786 & ~n7787 ) ;
  assign n7789 = ( x67 & n7783 ) | ( x67 & ~n7788 ) | ( n7783 & ~n7788 ) ;
  assign n7790 = ( x67 & n7486 ) | ( x67 & ~n7767 ) | ( n7486 & ~n7767 ) ;
  assign n7791 = x67 & n7486 ;
  assign n7792 = ( ~n7491 & n7790 ) | ( ~n7491 & n7791 ) | ( n7790 & n7791 ) ;
  assign n7793 = ( n7491 & n7790 ) | ( n7491 & n7791 ) | ( n7790 & n7791 ) ;
  assign n7794 = ( n7491 & n7792 ) | ( n7491 & ~n7793 ) | ( n7792 & ~n7793 ) ;
  assign n7795 = ( x68 & n7789 ) | ( x68 & ~n7794 ) | ( n7789 & ~n7794 ) ;
  assign n7796 = ( x68 & n7492 ) | ( x68 & ~n7767 ) | ( n7492 & ~n7767 ) ;
  assign n7797 = x68 & n7492 ;
  assign n7798 = ( ~n7497 & n7796 ) | ( ~n7497 & n7797 ) | ( n7796 & n7797 ) ;
  assign n7799 = ( n7497 & n7796 ) | ( n7497 & n7797 ) | ( n7796 & n7797 ) ;
  assign n7800 = ( n7497 & n7798 ) | ( n7497 & ~n7799 ) | ( n7798 & ~n7799 ) ;
  assign n7801 = ( x69 & n7795 ) | ( x69 & ~n7800 ) | ( n7795 & ~n7800 ) ;
  assign n7802 = ( x69 & n7498 ) | ( x69 & ~n7767 ) | ( n7498 & ~n7767 ) ;
  assign n7803 = x69 & n7498 ;
  assign n7804 = ( ~n7503 & n7802 ) | ( ~n7503 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7805 = ( n7503 & n7802 ) | ( n7503 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7806 = ( n7503 & n7804 ) | ( n7503 & ~n7805 ) | ( n7804 & ~n7805 ) ;
  assign n7807 = ( x70 & n7801 ) | ( x70 & ~n7806 ) | ( n7801 & ~n7806 ) ;
  assign n7808 = ( x70 & n7504 ) | ( x70 & ~n7767 ) | ( n7504 & ~n7767 ) ;
  assign n7809 = x70 & n7504 ;
  assign n7810 = ( ~n7509 & n7808 ) | ( ~n7509 & n7809 ) | ( n7808 & n7809 ) ;
  assign n7811 = ( n7509 & n7808 ) | ( n7509 & n7809 ) | ( n7808 & n7809 ) ;
  assign n7812 = ( n7509 & n7810 ) | ( n7509 & ~n7811 ) | ( n7810 & ~n7811 ) ;
  assign n7813 = ( x71 & n7807 ) | ( x71 & ~n7812 ) | ( n7807 & ~n7812 ) ;
  assign n7814 = ( x71 & n7510 ) | ( x71 & ~n7767 ) | ( n7510 & ~n7767 ) ;
  assign n7815 = x71 & n7510 ;
  assign n7816 = ( ~n7515 & n7814 ) | ( ~n7515 & n7815 ) | ( n7814 & n7815 ) ;
  assign n7817 = ( n7515 & n7814 ) | ( n7515 & n7815 ) | ( n7814 & n7815 ) ;
  assign n7818 = ( n7515 & n7816 ) | ( n7515 & ~n7817 ) | ( n7816 & ~n7817 ) ;
  assign n7819 = ( x72 & n7813 ) | ( x72 & ~n7818 ) | ( n7813 & ~n7818 ) ;
  assign n7820 = ( x72 & n7516 ) | ( x72 & ~n7767 ) | ( n7516 & ~n7767 ) ;
  assign n7821 = x72 & n7516 ;
  assign n7822 = ( ~n7521 & n7820 ) | ( ~n7521 & n7821 ) | ( n7820 & n7821 ) ;
  assign n7823 = ( n7521 & n7820 ) | ( n7521 & n7821 ) | ( n7820 & n7821 ) ;
  assign n7824 = ( n7521 & n7822 ) | ( n7521 & ~n7823 ) | ( n7822 & ~n7823 ) ;
  assign n7825 = ( x73 & n7819 ) | ( x73 & ~n7824 ) | ( n7819 & ~n7824 ) ;
  assign n7826 = ( x73 & n7522 ) | ( x73 & ~n7767 ) | ( n7522 & ~n7767 ) ;
  assign n7827 = x73 & n7522 ;
  assign n7828 = ( ~n7527 & n7826 ) | ( ~n7527 & n7827 ) | ( n7826 & n7827 ) ;
  assign n7829 = ( n7527 & n7826 ) | ( n7527 & n7827 ) | ( n7826 & n7827 ) ;
  assign n7830 = ( n7527 & n7828 ) | ( n7527 & ~n7829 ) | ( n7828 & ~n7829 ) ;
  assign n7831 = ( x74 & n7825 ) | ( x74 & ~n7830 ) | ( n7825 & ~n7830 ) ;
  assign n7832 = ( x74 & n7528 ) | ( x74 & ~n7767 ) | ( n7528 & ~n7767 ) ;
  assign n7833 = x74 & n7528 ;
  assign n7834 = ( ~n7533 & n7832 ) | ( ~n7533 & n7833 ) | ( n7832 & n7833 ) ;
  assign n7835 = ( n7533 & n7832 ) | ( n7533 & n7833 ) | ( n7832 & n7833 ) ;
  assign n7836 = ( n7533 & n7834 ) | ( n7533 & ~n7835 ) | ( n7834 & ~n7835 ) ;
  assign n7837 = ( x75 & n7831 ) | ( x75 & ~n7836 ) | ( n7831 & ~n7836 ) ;
  assign n7838 = ( x75 & n7534 ) | ( x75 & ~n7767 ) | ( n7534 & ~n7767 ) ;
  assign n7839 = x75 & n7534 ;
  assign n7840 = ( ~n7539 & n7838 ) | ( ~n7539 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7841 = ( n7539 & n7838 ) | ( n7539 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7842 = ( n7539 & n7840 ) | ( n7539 & ~n7841 ) | ( n7840 & ~n7841 ) ;
  assign n7843 = ( x76 & n7837 ) | ( x76 & ~n7842 ) | ( n7837 & ~n7842 ) ;
  assign n7844 = ( x76 & n7540 ) | ( x76 & ~n7767 ) | ( n7540 & ~n7767 ) ;
  assign n7845 = x76 & n7540 ;
  assign n7846 = ( ~n7545 & n7844 ) | ( ~n7545 & n7845 ) | ( n7844 & n7845 ) ;
  assign n7847 = ( n7545 & n7844 ) | ( n7545 & n7845 ) | ( n7844 & n7845 ) ;
  assign n7848 = ( n7545 & n7846 ) | ( n7545 & ~n7847 ) | ( n7846 & ~n7847 ) ;
  assign n7849 = ( x77 & n7843 ) | ( x77 & ~n7848 ) | ( n7843 & ~n7848 ) ;
  assign n7850 = ( x77 & n7546 ) | ( x77 & ~n7767 ) | ( n7546 & ~n7767 ) ;
  assign n7851 = x77 & n7546 ;
  assign n7852 = ( ~n7551 & n7850 ) | ( ~n7551 & n7851 ) | ( n7850 & n7851 ) ;
  assign n7853 = ( n7551 & n7850 ) | ( n7551 & n7851 ) | ( n7850 & n7851 ) ;
  assign n7854 = ( n7551 & n7852 ) | ( n7551 & ~n7853 ) | ( n7852 & ~n7853 ) ;
  assign n7855 = ( x78 & n7849 ) | ( x78 & ~n7854 ) | ( n7849 & ~n7854 ) ;
  assign n7856 = ( x78 & n7552 ) | ( x78 & ~n7767 ) | ( n7552 & ~n7767 ) ;
  assign n7857 = x78 & n7552 ;
  assign n7858 = ( ~n7557 & n7856 ) | ( ~n7557 & n7857 ) | ( n7856 & n7857 ) ;
  assign n7859 = ( n7557 & n7856 ) | ( n7557 & n7857 ) | ( n7856 & n7857 ) ;
  assign n7860 = ( n7557 & n7858 ) | ( n7557 & ~n7859 ) | ( n7858 & ~n7859 ) ;
  assign n7861 = ( x79 & n7855 ) | ( x79 & ~n7860 ) | ( n7855 & ~n7860 ) ;
  assign n7862 = ( x79 & n7558 ) | ( x79 & ~n7767 ) | ( n7558 & ~n7767 ) ;
  assign n7863 = x79 & n7558 ;
  assign n7864 = ( ~n7563 & n7862 ) | ( ~n7563 & n7863 ) | ( n7862 & n7863 ) ;
  assign n7865 = ( n7563 & n7862 ) | ( n7563 & n7863 ) | ( n7862 & n7863 ) ;
  assign n7866 = ( n7563 & n7864 ) | ( n7563 & ~n7865 ) | ( n7864 & ~n7865 ) ;
  assign n7867 = ( x80 & n7861 ) | ( x80 & ~n7866 ) | ( n7861 & ~n7866 ) ;
  assign n7868 = ( x80 & n7564 ) | ( x80 & ~n7767 ) | ( n7564 & ~n7767 ) ;
  assign n7869 = x80 & n7564 ;
  assign n7870 = ( ~n7569 & n7868 ) | ( ~n7569 & n7869 ) | ( n7868 & n7869 ) ;
  assign n7871 = ( n7569 & n7868 ) | ( n7569 & n7869 ) | ( n7868 & n7869 ) ;
  assign n7872 = ( n7569 & n7870 ) | ( n7569 & ~n7871 ) | ( n7870 & ~n7871 ) ;
  assign n7873 = ( x81 & n7867 ) | ( x81 & ~n7872 ) | ( n7867 & ~n7872 ) ;
  assign n7874 = ( x81 & n7570 ) | ( x81 & ~n7767 ) | ( n7570 & ~n7767 ) ;
  assign n7875 = x81 & n7570 ;
  assign n7876 = ( ~n7575 & n7874 ) | ( ~n7575 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7877 = ( n7575 & n7874 ) | ( n7575 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7878 = ( n7575 & n7876 ) | ( n7575 & ~n7877 ) | ( n7876 & ~n7877 ) ;
  assign n7879 = ( x82 & n7873 ) | ( x82 & ~n7878 ) | ( n7873 & ~n7878 ) ;
  assign n7880 = ( x82 & n7576 ) | ( x82 & ~n7767 ) | ( n7576 & ~n7767 ) ;
  assign n7881 = x82 & n7576 ;
  assign n7882 = ( ~n7581 & n7880 ) | ( ~n7581 & n7881 ) | ( n7880 & n7881 ) ;
  assign n7883 = ( n7581 & n7880 ) | ( n7581 & n7881 ) | ( n7880 & n7881 ) ;
  assign n7884 = ( n7581 & n7882 ) | ( n7581 & ~n7883 ) | ( n7882 & ~n7883 ) ;
  assign n7885 = ( x83 & n7879 ) | ( x83 & ~n7884 ) | ( n7879 & ~n7884 ) ;
  assign n7886 = ( x83 & n7582 ) | ( x83 & ~n7767 ) | ( n7582 & ~n7767 ) ;
  assign n7887 = x83 & n7582 ;
  assign n7888 = ( ~n7587 & n7886 ) | ( ~n7587 & n7887 ) | ( n7886 & n7887 ) ;
  assign n7889 = ( n7587 & n7886 ) | ( n7587 & n7887 ) | ( n7886 & n7887 ) ;
  assign n7890 = ( n7587 & n7888 ) | ( n7587 & ~n7889 ) | ( n7888 & ~n7889 ) ;
  assign n7891 = ( x84 & n7885 ) | ( x84 & ~n7890 ) | ( n7885 & ~n7890 ) ;
  assign n7892 = ( x84 & n7588 ) | ( x84 & ~n7767 ) | ( n7588 & ~n7767 ) ;
  assign n7893 = x84 & n7588 ;
  assign n7894 = ( ~n7593 & n7892 ) | ( ~n7593 & n7893 ) | ( n7892 & n7893 ) ;
  assign n7895 = ( n7593 & n7892 ) | ( n7593 & n7893 ) | ( n7892 & n7893 ) ;
  assign n7896 = ( n7593 & n7894 ) | ( n7593 & ~n7895 ) | ( n7894 & ~n7895 ) ;
  assign n7897 = ( x85 & n7891 ) | ( x85 & ~n7896 ) | ( n7891 & ~n7896 ) ;
  assign n7898 = ( x85 & n7594 ) | ( x85 & ~n7767 ) | ( n7594 & ~n7767 ) ;
  assign n7899 = x85 & n7594 ;
  assign n7900 = ( ~n7599 & n7898 ) | ( ~n7599 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7901 = ( n7599 & n7898 ) | ( n7599 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7902 = ( n7599 & n7900 ) | ( n7599 & ~n7901 ) | ( n7900 & ~n7901 ) ;
  assign n7903 = ( x86 & n7897 ) | ( x86 & ~n7902 ) | ( n7897 & ~n7902 ) ;
  assign n7904 = ( x86 & n7600 ) | ( x86 & ~n7767 ) | ( n7600 & ~n7767 ) ;
  assign n7905 = x86 & n7600 ;
  assign n7906 = ( ~n7605 & n7904 ) | ( ~n7605 & n7905 ) | ( n7904 & n7905 ) ;
  assign n7907 = ( n7605 & n7904 ) | ( n7605 & n7905 ) | ( n7904 & n7905 ) ;
  assign n7908 = ( n7605 & n7906 ) | ( n7605 & ~n7907 ) | ( n7906 & ~n7907 ) ;
  assign n7909 = ( x87 & n7903 ) | ( x87 & ~n7908 ) | ( n7903 & ~n7908 ) ;
  assign n7910 = ( x87 & n7606 ) | ( x87 & ~n7767 ) | ( n7606 & ~n7767 ) ;
  assign n7911 = x87 & n7606 ;
  assign n7912 = ( ~n7611 & n7910 ) | ( ~n7611 & n7911 ) | ( n7910 & n7911 ) ;
  assign n7913 = ( n7611 & n7910 ) | ( n7611 & n7911 ) | ( n7910 & n7911 ) ;
  assign n7914 = ( n7611 & n7912 ) | ( n7611 & ~n7913 ) | ( n7912 & ~n7913 ) ;
  assign n7915 = ( x88 & n7909 ) | ( x88 & ~n7914 ) | ( n7909 & ~n7914 ) ;
  assign n7916 = ( x88 & n7612 ) | ( x88 & ~n7767 ) | ( n7612 & ~n7767 ) ;
  assign n7917 = x88 & n7612 ;
  assign n7918 = ( ~n7617 & n7916 ) | ( ~n7617 & n7917 ) | ( n7916 & n7917 ) ;
  assign n7919 = ( n7617 & n7916 ) | ( n7617 & n7917 ) | ( n7916 & n7917 ) ;
  assign n7920 = ( n7617 & n7918 ) | ( n7617 & ~n7919 ) | ( n7918 & ~n7919 ) ;
  assign n7921 = ( x89 & n7915 ) | ( x89 & ~n7920 ) | ( n7915 & ~n7920 ) ;
  assign n7922 = ( x89 & n7618 ) | ( x89 & ~n7767 ) | ( n7618 & ~n7767 ) ;
  assign n7923 = x89 & n7618 ;
  assign n7924 = ( ~n7623 & n7922 ) | ( ~n7623 & n7923 ) | ( n7922 & n7923 ) ;
  assign n7925 = ( n7623 & n7922 ) | ( n7623 & n7923 ) | ( n7922 & n7923 ) ;
  assign n7926 = ( n7623 & n7924 ) | ( n7623 & ~n7925 ) | ( n7924 & ~n7925 ) ;
  assign n7927 = ( x90 & n7921 ) | ( x90 & ~n7926 ) | ( n7921 & ~n7926 ) ;
  assign n7928 = ( x90 & n7624 ) | ( x90 & ~n7767 ) | ( n7624 & ~n7767 ) ;
  assign n7929 = x90 & n7624 ;
  assign n7930 = ( ~n7629 & n7928 ) | ( ~n7629 & n7929 ) | ( n7928 & n7929 ) ;
  assign n7931 = ( n7629 & n7928 ) | ( n7629 & n7929 ) | ( n7928 & n7929 ) ;
  assign n7932 = ( n7629 & n7930 ) | ( n7629 & ~n7931 ) | ( n7930 & ~n7931 ) ;
  assign n7933 = ( x91 & n7927 ) | ( x91 & ~n7932 ) | ( n7927 & ~n7932 ) ;
  assign n7934 = ( x91 & n7630 ) | ( x91 & ~n7767 ) | ( n7630 & ~n7767 ) ;
  assign n7935 = x91 & n7630 ;
  assign n7936 = ( ~n7635 & n7934 ) | ( ~n7635 & n7935 ) | ( n7934 & n7935 ) ;
  assign n7937 = ( n7635 & n7934 ) | ( n7635 & n7935 ) | ( n7934 & n7935 ) ;
  assign n7938 = ( n7635 & n7936 ) | ( n7635 & ~n7937 ) | ( n7936 & ~n7937 ) ;
  assign n7939 = ( x92 & n7933 ) | ( x92 & ~n7938 ) | ( n7933 & ~n7938 ) ;
  assign n7940 = ( x92 & n7636 ) | ( x92 & ~n7767 ) | ( n7636 & ~n7767 ) ;
  assign n7941 = x92 & n7636 ;
  assign n7942 = ( ~n7641 & n7940 ) | ( ~n7641 & n7941 ) | ( n7940 & n7941 ) ;
  assign n7943 = ( n7641 & n7940 ) | ( n7641 & n7941 ) | ( n7940 & n7941 ) ;
  assign n7944 = ( n7641 & n7942 ) | ( n7641 & ~n7943 ) | ( n7942 & ~n7943 ) ;
  assign n7945 = ( x93 & n7939 ) | ( x93 & ~n7944 ) | ( n7939 & ~n7944 ) ;
  assign n7946 = ( x93 & n7642 ) | ( x93 & ~n7767 ) | ( n7642 & ~n7767 ) ;
  assign n7947 = x93 & n7642 ;
  assign n7948 = ( ~n7647 & n7946 ) | ( ~n7647 & n7947 ) | ( n7946 & n7947 ) ;
  assign n7949 = ( n7647 & n7946 ) | ( n7647 & n7947 ) | ( n7946 & n7947 ) ;
  assign n7950 = ( n7647 & n7948 ) | ( n7647 & ~n7949 ) | ( n7948 & ~n7949 ) ;
  assign n7951 = ( x94 & n7945 ) | ( x94 & ~n7950 ) | ( n7945 & ~n7950 ) ;
  assign n7952 = ( x94 & n7648 ) | ( x94 & ~n7767 ) | ( n7648 & ~n7767 ) ;
  assign n7953 = x94 & n7648 ;
  assign n7954 = ( ~n7653 & n7952 ) | ( ~n7653 & n7953 ) | ( n7952 & n7953 ) ;
  assign n7955 = ( n7653 & n7952 ) | ( n7653 & n7953 ) | ( n7952 & n7953 ) ;
  assign n7956 = ( n7653 & n7954 ) | ( n7653 & ~n7955 ) | ( n7954 & ~n7955 ) ;
  assign n7957 = ( x95 & n7951 ) | ( x95 & ~n7956 ) | ( n7951 & ~n7956 ) ;
  assign n7958 = ( x95 & n7654 ) | ( x95 & ~n7767 ) | ( n7654 & ~n7767 ) ;
  assign n7959 = x95 & n7654 ;
  assign n7960 = ( ~n7659 & n7958 ) | ( ~n7659 & n7959 ) | ( n7958 & n7959 ) ;
  assign n7961 = ( n7659 & n7958 ) | ( n7659 & n7959 ) | ( n7958 & n7959 ) ;
  assign n7962 = ( n7659 & n7960 ) | ( n7659 & ~n7961 ) | ( n7960 & ~n7961 ) ;
  assign n7963 = ( x96 & n7957 ) | ( x96 & ~n7962 ) | ( n7957 & ~n7962 ) ;
  assign n7964 = ( x96 & n7660 ) | ( x96 & ~n7767 ) | ( n7660 & ~n7767 ) ;
  assign n7965 = x96 & n7660 ;
  assign n7966 = ( ~n7665 & n7964 ) | ( ~n7665 & n7965 ) | ( n7964 & n7965 ) ;
  assign n7967 = ( n7665 & n7964 ) | ( n7665 & n7965 ) | ( n7964 & n7965 ) ;
  assign n7968 = ( n7665 & n7966 ) | ( n7665 & ~n7967 ) | ( n7966 & ~n7967 ) ;
  assign n7969 = ( x97 & n7963 ) | ( x97 & ~n7968 ) | ( n7963 & ~n7968 ) ;
  assign n7970 = ( x97 & n7666 ) | ( x97 & ~n7767 ) | ( n7666 & ~n7767 ) ;
  assign n7971 = x97 & n7666 ;
  assign n7972 = ( ~n7671 & n7970 ) | ( ~n7671 & n7971 ) | ( n7970 & n7971 ) ;
  assign n7973 = ( n7671 & n7970 ) | ( n7671 & n7971 ) | ( n7970 & n7971 ) ;
  assign n7974 = ( n7671 & n7972 ) | ( n7671 & ~n7973 ) | ( n7972 & ~n7973 ) ;
  assign n7975 = ( x98 & n7969 ) | ( x98 & ~n7974 ) | ( n7969 & ~n7974 ) ;
  assign n7976 = ( x98 & n7672 ) | ( x98 & ~n7767 ) | ( n7672 & ~n7767 ) ;
  assign n7977 = x98 & n7672 ;
  assign n7978 = ( ~n7677 & n7976 ) | ( ~n7677 & n7977 ) | ( n7976 & n7977 ) ;
  assign n7979 = ( n7677 & n7976 ) | ( n7677 & n7977 ) | ( n7976 & n7977 ) ;
  assign n7980 = ( n7677 & n7978 ) | ( n7677 & ~n7979 ) | ( n7978 & ~n7979 ) ;
  assign n7981 = ( x99 & n7975 ) | ( x99 & ~n7980 ) | ( n7975 & ~n7980 ) ;
  assign n7982 = ( x99 & n7678 ) | ( x99 & ~n7767 ) | ( n7678 & ~n7767 ) ;
  assign n7983 = x99 & n7678 ;
  assign n7984 = ( ~n7683 & n7982 ) | ( ~n7683 & n7983 ) | ( n7982 & n7983 ) ;
  assign n7985 = ( n7683 & n7982 ) | ( n7683 & n7983 ) | ( n7982 & n7983 ) ;
  assign n7986 = ( n7683 & n7984 ) | ( n7683 & ~n7985 ) | ( n7984 & ~n7985 ) ;
  assign n7987 = ( x100 & n7981 ) | ( x100 & ~n7986 ) | ( n7981 & ~n7986 ) ;
  assign n7988 = ( x100 & n7684 ) | ( x100 & ~n7767 ) | ( n7684 & ~n7767 ) ;
  assign n7989 = x100 & n7684 ;
  assign n7990 = ( ~n7689 & n7988 ) | ( ~n7689 & n7989 ) | ( n7988 & n7989 ) ;
  assign n7991 = ( n7689 & n7988 ) | ( n7689 & n7989 ) | ( n7988 & n7989 ) ;
  assign n7992 = ( n7689 & n7990 ) | ( n7689 & ~n7991 ) | ( n7990 & ~n7991 ) ;
  assign n7993 = ( x101 & n7987 ) | ( x101 & ~n7992 ) | ( n7987 & ~n7992 ) ;
  assign n7994 = ( x101 & n7690 ) | ( x101 & ~n7767 ) | ( n7690 & ~n7767 ) ;
  assign n7995 = x101 & n7690 ;
  assign n7996 = ( ~n7695 & n7994 ) | ( ~n7695 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7997 = ( n7695 & n7994 ) | ( n7695 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7998 = ( n7695 & n7996 ) | ( n7695 & ~n7997 ) | ( n7996 & ~n7997 ) ;
  assign n7999 = ( x102 & n7993 ) | ( x102 & ~n7998 ) | ( n7993 & ~n7998 ) ;
  assign n8000 = ( x102 & n7696 ) | ( x102 & ~n7767 ) | ( n7696 & ~n7767 ) ;
  assign n8001 = x102 & n7696 ;
  assign n8002 = ( ~n7701 & n8000 ) | ( ~n7701 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8003 = ( n7701 & n8000 ) | ( n7701 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8004 = ( n7701 & n8002 ) | ( n7701 & ~n8003 ) | ( n8002 & ~n8003 ) ;
  assign n8005 = ( x103 & n7999 ) | ( x103 & ~n8004 ) | ( n7999 & ~n8004 ) ;
  assign n8006 = ( x103 & n7702 ) | ( x103 & ~n7767 ) | ( n7702 & ~n7767 ) ;
  assign n8007 = x103 & n7702 ;
  assign n8008 = ( ~n7707 & n8006 ) | ( ~n7707 & n8007 ) | ( n8006 & n8007 ) ;
  assign n8009 = ( n7707 & n8006 ) | ( n7707 & n8007 ) | ( n8006 & n8007 ) ;
  assign n8010 = ( n7707 & n8008 ) | ( n7707 & ~n8009 ) | ( n8008 & ~n8009 ) ;
  assign n8011 = ( x104 & n8005 ) | ( x104 & ~n8010 ) | ( n8005 & ~n8010 ) ;
  assign n8012 = ( x104 & n7708 ) | ( x104 & ~n7767 ) | ( n7708 & ~n7767 ) ;
  assign n8013 = x104 & n7708 ;
  assign n8014 = ( ~n7713 & n8012 ) | ( ~n7713 & n8013 ) | ( n8012 & n8013 ) ;
  assign n8015 = ( n7713 & n8012 ) | ( n7713 & n8013 ) | ( n8012 & n8013 ) ;
  assign n8016 = ( n7713 & n8014 ) | ( n7713 & ~n8015 ) | ( n8014 & ~n8015 ) ;
  assign n8017 = ( x105 & n8011 ) | ( x105 & ~n8016 ) | ( n8011 & ~n8016 ) ;
  assign n8018 = ( x105 & n7714 ) | ( x105 & ~n7767 ) | ( n7714 & ~n7767 ) ;
  assign n8019 = x105 & n7714 ;
  assign n8020 = ( ~n7719 & n8018 ) | ( ~n7719 & n8019 ) | ( n8018 & n8019 ) ;
  assign n8021 = ( n7719 & n8018 ) | ( n7719 & n8019 ) | ( n8018 & n8019 ) ;
  assign n8022 = ( n7719 & n8020 ) | ( n7719 & ~n8021 ) | ( n8020 & ~n8021 ) ;
  assign n8023 = ( x106 & n8017 ) | ( x106 & ~n8022 ) | ( n8017 & ~n8022 ) ;
  assign n8024 = ( x106 & n7720 ) | ( x106 & ~n7767 ) | ( n7720 & ~n7767 ) ;
  assign n8025 = x106 & n7720 ;
  assign n8026 = ( ~n7725 & n8024 ) | ( ~n7725 & n8025 ) | ( n8024 & n8025 ) ;
  assign n8027 = ( n7725 & n8024 ) | ( n7725 & n8025 ) | ( n8024 & n8025 ) ;
  assign n8028 = ( n7725 & n8026 ) | ( n7725 & ~n8027 ) | ( n8026 & ~n8027 ) ;
  assign n8029 = ( x107 & n8023 ) | ( x107 & ~n8028 ) | ( n8023 & ~n8028 ) ;
  assign n8030 = ( x107 & n7726 ) | ( x107 & ~n7767 ) | ( n7726 & ~n7767 ) ;
  assign n8031 = x107 & n7726 ;
  assign n8032 = ( ~n7731 & n8030 ) | ( ~n7731 & n8031 ) | ( n8030 & n8031 ) ;
  assign n8033 = ( n7731 & n8030 ) | ( n7731 & n8031 ) | ( n8030 & n8031 ) ;
  assign n8034 = ( n7731 & n8032 ) | ( n7731 & ~n8033 ) | ( n8032 & ~n8033 ) ;
  assign n8035 = ( x108 & n8029 ) | ( x108 & ~n8034 ) | ( n8029 & ~n8034 ) ;
  assign n8036 = ( x108 & n7732 ) | ( x108 & ~n7767 ) | ( n7732 & ~n7767 ) ;
  assign n8037 = x108 & n7732 ;
  assign n8038 = ( ~n7737 & n8036 ) | ( ~n7737 & n8037 ) | ( n8036 & n8037 ) ;
  assign n8039 = ( n7737 & n8036 ) | ( n7737 & n8037 ) | ( n8036 & n8037 ) ;
  assign n8040 = ( n7737 & n8038 ) | ( n7737 & ~n8039 ) | ( n8038 & ~n8039 ) ;
  assign n8041 = ( x109 & n8035 ) | ( x109 & ~n8040 ) | ( n8035 & ~n8040 ) ;
  assign n8042 = ( x109 & n7738 ) | ( x109 & ~n7767 ) | ( n7738 & ~n7767 ) ;
  assign n8043 = x109 & n7738 ;
  assign n8044 = ( ~n7743 & n8042 ) | ( ~n7743 & n8043 ) | ( n8042 & n8043 ) ;
  assign n8045 = ( n7743 & n8042 ) | ( n7743 & n8043 ) | ( n8042 & n8043 ) ;
  assign n8046 = ( n7743 & n8044 ) | ( n7743 & ~n8045 ) | ( n8044 & ~n8045 ) ;
  assign n8047 = ( x110 & n8041 ) | ( x110 & ~n8046 ) | ( n8041 & ~n8046 ) ;
  assign n8048 = ( x110 & n7744 ) | ( x110 & ~n7767 ) | ( n7744 & ~n7767 ) ;
  assign n8049 = x110 & n7744 ;
  assign n8050 = ( ~n7749 & n8048 ) | ( ~n7749 & n8049 ) | ( n8048 & n8049 ) ;
  assign n8051 = ( n7749 & n8048 ) | ( n7749 & n8049 ) | ( n8048 & n8049 ) ;
  assign n8052 = ( n7749 & n8050 ) | ( n7749 & ~n8051 ) | ( n8050 & ~n8051 ) ;
  assign n8053 = ( x111 & n8047 ) | ( x111 & ~n8052 ) | ( n8047 & ~n8052 ) ;
  assign n8054 = ( x111 & n7750 ) | ( x111 & ~n7767 ) | ( n7750 & ~n7767 ) ;
  assign n8055 = x111 & n7750 ;
  assign n8056 = ( ~n7755 & n8054 ) | ( ~n7755 & n8055 ) | ( n8054 & n8055 ) ;
  assign n8057 = ( n7755 & n8054 ) | ( n7755 & n8055 ) | ( n8054 & n8055 ) ;
  assign n8058 = ( n7755 & n8056 ) | ( n7755 & ~n8057 ) | ( n8056 & ~n8057 ) ;
  assign n8059 = ( x112 & n8053 ) | ( x112 & ~n8058 ) | ( n8053 & ~n8058 ) ;
  assign n8060 = ( x112 & n7756 ) | ( x112 & ~n7767 ) | ( n7756 & ~n7767 ) ;
  assign n8061 = x112 & n7756 ;
  assign n8062 = ( ~n7761 & n8060 ) | ( ~n7761 & n8061 ) | ( n8060 & n8061 ) ;
  assign n8063 = ( n7761 & n8060 ) | ( n7761 & n8061 ) | ( n8060 & n8061 ) ;
  assign n8064 = ( n7761 & n8062 ) | ( n7761 & ~n8063 ) | ( n8062 & ~n8063 ) ;
  assign n8065 = ( x113 & n8059 ) | ( x113 & ~n8064 ) | ( n8059 & ~n8064 ) ;
  assign n8066 = ( x114 & n142 ) | ( x114 & n7763 ) | ( n142 & n7763 ) ;
  assign n8067 = x114 | n7763 ;
  assign n8068 = ( n7765 & n8066 ) | ( n7765 & ~n8067 ) | ( n8066 & ~n8067 ) ;
  assign n8069 = ( x114 & ~n7772 ) | ( x114 & n8065 ) | ( ~n7772 & n8065 ) ;
  assign n8070 = ( x115 & ~n8068 ) | ( x115 & n8069 ) | ( ~n8068 & n8069 ) ;
  assign n8071 = n141 | n8070 ;
  assign n8072 = ( x114 & n8065 ) | ( x114 & n8071 ) | ( n8065 & n8071 ) ;
  assign n8073 = x114 | n8065 ;
  assign n8074 = ( ~n7772 & n8072 ) | ( ~n7772 & n8073 ) | ( n8072 & n8073 ) ;
  assign n8075 = ( n7772 & n8072 ) | ( n7772 & n8073 ) | ( n8072 & n8073 ) ;
  assign n8076 = ( n7772 & n8074 ) | ( n7772 & ~n8075 ) | ( n8074 & ~n8075 ) ;
  assign n8077 = ~x11 & x64 ;
  assign n8078 = ~x12 & n8071 ;
  assign n8079 = ( x12 & ~x64 ) | ( x12 & n8071 ) | ( ~x64 & n8071 ) ;
  assign n8080 = ( n7773 & ~n8078 ) | ( n7773 & n8079 ) | ( ~n8078 & n8079 ) ;
  assign n8081 = ( x65 & n8077 ) | ( x65 & ~n8080 ) | ( n8077 & ~n8080 ) ;
  assign n8082 = ( x65 & n7773 ) | ( x65 & n8071 ) | ( n7773 & n8071 ) ;
  assign n8083 = x65 | n7773 ;
  assign n8084 = ( ~n7776 & n8082 ) | ( ~n7776 & n8083 ) | ( n8082 & n8083 ) ;
  assign n8085 = ( n7776 & n8082 ) | ( n7776 & n8083 ) | ( n8082 & n8083 ) ;
  assign n8086 = ( n7776 & n8084 ) | ( n7776 & ~n8085 ) | ( n8084 & ~n8085 ) ;
  assign n8087 = ( x66 & n8081 ) | ( x66 & ~n8086 ) | ( n8081 & ~n8086 ) ;
  assign n8088 = ( x66 & n7777 ) | ( x66 & n8071 ) | ( n7777 & n8071 ) ;
  assign n8089 = x66 | n7777 ;
  assign n8090 = ( ~n7782 & n8088 ) | ( ~n7782 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8091 = ( n7782 & n8088 ) | ( n7782 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8092 = ( n7782 & n8090 ) | ( n7782 & ~n8091 ) | ( n8090 & ~n8091 ) ;
  assign n8093 = ( x67 & n8087 ) | ( x67 & ~n8092 ) | ( n8087 & ~n8092 ) ;
  assign n8094 = ( x67 & n7783 ) | ( x67 & ~n8071 ) | ( n7783 & ~n8071 ) ;
  assign n8095 = x67 & n7783 ;
  assign n8096 = ( ~n7788 & n8094 ) | ( ~n7788 & n8095 ) | ( n8094 & n8095 ) ;
  assign n8097 = ( n7788 & n8094 ) | ( n7788 & n8095 ) | ( n8094 & n8095 ) ;
  assign n8098 = ( n7788 & n8096 ) | ( n7788 & ~n8097 ) | ( n8096 & ~n8097 ) ;
  assign n8099 = ( x68 & n8093 ) | ( x68 & ~n8098 ) | ( n8093 & ~n8098 ) ;
  assign n8100 = ( x68 & n7789 ) | ( x68 & ~n8071 ) | ( n7789 & ~n8071 ) ;
  assign n8101 = x68 & n7789 ;
  assign n8102 = ( ~n7794 & n8100 ) | ( ~n7794 & n8101 ) | ( n8100 & n8101 ) ;
  assign n8103 = ( n7794 & n8100 ) | ( n7794 & n8101 ) | ( n8100 & n8101 ) ;
  assign n8104 = ( n7794 & n8102 ) | ( n7794 & ~n8103 ) | ( n8102 & ~n8103 ) ;
  assign n8105 = ( x69 & n8099 ) | ( x69 & ~n8104 ) | ( n8099 & ~n8104 ) ;
  assign n8106 = ( x69 & n7795 ) | ( x69 & ~n8071 ) | ( n7795 & ~n8071 ) ;
  assign n8107 = x69 & n7795 ;
  assign n8108 = ( ~n7800 & n8106 ) | ( ~n7800 & n8107 ) | ( n8106 & n8107 ) ;
  assign n8109 = ( n7800 & n8106 ) | ( n7800 & n8107 ) | ( n8106 & n8107 ) ;
  assign n8110 = ( n7800 & n8108 ) | ( n7800 & ~n8109 ) | ( n8108 & ~n8109 ) ;
  assign n8111 = ( x70 & n8105 ) | ( x70 & ~n8110 ) | ( n8105 & ~n8110 ) ;
  assign n8112 = ( x70 & n7801 ) | ( x70 & ~n8071 ) | ( n7801 & ~n8071 ) ;
  assign n8113 = x70 & n7801 ;
  assign n8114 = ( ~n7806 & n8112 ) | ( ~n7806 & n8113 ) | ( n8112 & n8113 ) ;
  assign n8115 = ( n7806 & n8112 ) | ( n7806 & n8113 ) | ( n8112 & n8113 ) ;
  assign n8116 = ( n7806 & n8114 ) | ( n7806 & ~n8115 ) | ( n8114 & ~n8115 ) ;
  assign n8117 = ( x71 & n8111 ) | ( x71 & ~n8116 ) | ( n8111 & ~n8116 ) ;
  assign n8118 = ( x71 & n7807 ) | ( x71 & ~n8071 ) | ( n7807 & ~n8071 ) ;
  assign n8119 = x71 & n7807 ;
  assign n8120 = ( ~n7812 & n8118 ) | ( ~n7812 & n8119 ) | ( n8118 & n8119 ) ;
  assign n8121 = ( n7812 & n8118 ) | ( n7812 & n8119 ) | ( n8118 & n8119 ) ;
  assign n8122 = ( n7812 & n8120 ) | ( n7812 & ~n8121 ) | ( n8120 & ~n8121 ) ;
  assign n8123 = ( x72 & n8117 ) | ( x72 & ~n8122 ) | ( n8117 & ~n8122 ) ;
  assign n8124 = ( x72 & n7813 ) | ( x72 & ~n8071 ) | ( n7813 & ~n8071 ) ;
  assign n8125 = x72 & n7813 ;
  assign n8126 = ( ~n7818 & n8124 ) | ( ~n7818 & n8125 ) | ( n8124 & n8125 ) ;
  assign n8127 = ( n7818 & n8124 ) | ( n7818 & n8125 ) | ( n8124 & n8125 ) ;
  assign n8128 = ( n7818 & n8126 ) | ( n7818 & ~n8127 ) | ( n8126 & ~n8127 ) ;
  assign n8129 = ( x73 & n8123 ) | ( x73 & ~n8128 ) | ( n8123 & ~n8128 ) ;
  assign n8130 = ( x73 & n7819 ) | ( x73 & ~n8071 ) | ( n7819 & ~n8071 ) ;
  assign n8131 = x73 & n7819 ;
  assign n8132 = ( ~n7824 & n8130 ) | ( ~n7824 & n8131 ) | ( n8130 & n8131 ) ;
  assign n8133 = ( n7824 & n8130 ) | ( n7824 & n8131 ) | ( n8130 & n8131 ) ;
  assign n8134 = ( n7824 & n8132 ) | ( n7824 & ~n8133 ) | ( n8132 & ~n8133 ) ;
  assign n8135 = ( x74 & n8129 ) | ( x74 & ~n8134 ) | ( n8129 & ~n8134 ) ;
  assign n8136 = ( x74 & n7825 ) | ( x74 & ~n8071 ) | ( n7825 & ~n8071 ) ;
  assign n8137 = x74 & n7825 ;
  assign n8138 = ( ~n7830 & n8136 ) | ( ~n7830 & n8137 ) | ( n8136 & n8137 ) ;
  assign n8139 = ( n7830 & n8136 ) | ( n7830 & n8137 ) | ( n8136 & n8137 ) ;
  assign n8140 = ( n7830 & n8138 ) | ( n7830 & ~n8139 ) | ( n8138 & ~n8139 ) ;
  assign n8141 = ( x75 & n8135 ) | ( x75 & ~n8140 ) | ( n8135 & ~n8140 ) ;
  assign n8142 = ( x75 & n7831 ) | ( x75 & ~n8071 ) | ( n7831 & ~n8071 ) ;
  assign n8143 = x75 & n7831 ;
  assign n8144 = ( ~n7836 & n8142 ) | ( ~n7836 & n8143 ) | ( n8142 & n8143 ) ;
  assign n8145 = ( n7836 & n8142 ) | ( n7836 & n8143 ) | ( n8142 & n8143 ) ;
  assign n8146 = ( n7836 & n8144 ) | ( n7836 & ~n8145 ) | ( n8144 & ~n8145 ) ;
  assign n8147 = ( x76 & n8141 ) | ( x76 & ~n8146 ) | ( n8141 & ~n8146 ) ;
  assign n8148 = ( x76 & n7837 ) | ( x76 & ~n8071 ) | ( n7837 & ~n8071 ) ;
  assign n8149 = x76 & n7837 ;
  assign n8150 = ( ~n7842 & n8148 ) | ( ~n7842 & n8149 ) | ( n8148 & n8149 ) ;
  assign n8151 = ( n7842 & n8148 ) | ( n7842 & n8149 ) | ( n8148 & n8149 ) ;
  assign n8152 = ( n7842 & n8150 ) | ( n7842 & ~n8151 ) | ( n8150 & ~n8151 ) ;
  assign n8153 = ( x77 & n8147 ) | ( x77 & ~n8152 ) | ( n8147 & ~n8152 ) ;
  assign n8154 = ( x77 & n7843 ) | ( x77 & ~n8071 ) | ( n7843 & ~n8071 ) ;
  assign n8155 = x77 & n7843 ;
  assign n8156 = ( ~n7848 & n8154 ) | ( ~n7848 & n8155 ) | ( n8154 & n8155 ) ;
  assign n8157 = ( n7848 & n8154 ) | ( n7848 & n8155 ) | ( n8154 & n8155 ) ;
  assign n8158 = ( n7848 & n8156 ) | ( n7848 & ~n8157 ) | ( n8156 & ~n8157 ) ;
  assign n8159 = ( x78 & n8153 ) | ( x78 & ~n8158 ) | ( n8153 & ~n8158 ) ;
  assign n8160 = ( x78 & n7849 ) | ( x78 & ~n8071 ) | ( n7849 & ~n8071 ) ;
  assign n8161 = x78 & n7849 ;
  assign n8162 = ( ~n7854 & n8160 ) | ( ~n7854 & n8161 ) | ( n8160 & n8161 ) ;
  assign n8163 = ( n7854 & n8160 ) | ( n7854 & n8161 ) | ( n8160 & n8161 ) ;
  assign n8164 = ( n7854 & n8162 ) | ( n7854 & ~n8163 ) | ( n8162 & ~n8163 ) ;
  assign n8165 = ( x79 & n8159 ) | ( x79 & ~n8164 ) | ( n8159 & ~n8164 ) ;
  assign n8166 = ( x79 & n7855 ) | ( x79 & ~n8071 ) | ( n7855 & ~n8071 ) ;
  assign n8167 = x79 & n7855 ;
  assign n8168 = ( ~n7860 & n8166 ) | ( ~n7860 & n8167 ) | ( n8166 & n8167 ) ;
  assign n8169 = ( n7860 & n8166 ) | ( n7860 & n8167 ) | ( n8166 & n8167 ) ;
  assign n8170 = ( n7860 & n8168 ) | ( n7860 & ~n8169 ) | ( n8168 & ~n8169 ) ;
  assign n8171 = ( x80 & n8165 ) | ( x80 & ~n8170 ) | ( n8165 & ~n8170 ) ;
  assign n8172 = ( x80 & n7861 ) | ( x80 & ~n8071 ) | ( n7861 & ~n8071 ) ;
  assign n8173 = x80 & n7861 ;
  assign n8174 = ( ~n7866 & n8172 ) | ( ~n7866 & n8173 ) | ( n8172 & n8173 ) ;
  assign n8175 = ( n7866 & n8172 ) | ( n7866 & n8173 ) | ( n8172 & n8173 ) ;
  assign n8176 = ( n7866 & n8174 ) | ( n7866 & ~n8175 ) | ( n8174 & ~n8175 ) ;
  assign n8177 = ( x81 & n8171 ) | ( x81 & ~n8176 ) | ( n8171 & ~n8176 ) ;
  assign n8178 = ( x81 & n7867 ) | ( x81 & ~n8071 ) | ( n7867 & ~n8071 ) ;
  assign n8179 = x81 & n7867 ;
  assign n8180 = ( ~n7872 & n8178 ) | ( ~n7872 & n8179 ) | ( n8178 & n8179 ) ;
  assign n8181 = ( n7872 & n8178 ) | ( n7872 & n8179 ) | ( n8178 & n8179 ) ;
  assign n8182 = ( n7872 & n8180 ) | ( n7872 & ~n8181 ) | ( n8180 & ~n8181 ) ;
  assign n8183 = ( x82 & n8177 ) | ( x82 & ~n8182 ) | ( n8177 & ~n8182 ) ;
  assign n8184 = ( x82 & n7873 ) | ( x82 & ~n8071 ) | ( n7873 & ~n8071 ) ;
  assign n8185 = x82 & n7873 ;
  assign n8186 = ( ~n7878 & n8184 ) | ( ~n7878 & n8185 ) | ( n8184 & n8185 ) ;
  assign n8187 = ( n7878 & n8184 ) | ( n7878 & n8185 ) | ( n8184 & n8185 ) ;
  assign n8188 = ( n7878 & n8186 ) | ( n7878 & ~n8187 ) | ( n8186 & ~n8187 ) ;
  assign n8189 = ( x83 & n8183 ) | ( x83 & ~n8188 ) | ( n8183 & ~n8188 ) ;
  assign n8190 = ( x83 & n7879 ) | ( x83 & ~n8071 ) | ( n7879 & ~n8071 ) ;
  assign n8191 = x83 & n7879 ;
  assign n8192 = ( ~n7884 & n8190 ) | ( ~n7884 & n8191 ) | ( n8190 & n8191 ) ;
  assign n8193 = ( n7884 & n8190 ) | ( n7884 & n8191 ) | ( n8190 & n8191 ) ;
  assign n8194 = ( n7884 & n8192 ) | ( n7884 & ~n8193 ) | ( n8192 & ~n8193 ) ;
  assign n8195 = ( x84 & n8189 ) | ( x84 & ~n8194 ) | ( n8189 & ~n8194 ) ;
  assign n8196 = ( x84 & n7885 ) | ( x84 & ~n8071 ) | ( n7885 & ~n8071 ) ;
  assign n8197 = x84 & n7885 ;
  assign n8198 = ( ~n7890 & n8196 ) | ( ~n7890 & n8197 ) | ( n8196 & n8197 ) ;
  assign n8199 = ( n7890 & n8196 ) | ( n7890 & n8197 ) | ( n8196 & n8197 ) ;
  assign n8200 = ( n7890 & n8198 ) | ( n7890 & ~n8199 ) | ( n8198 & ~n8199 ) ;
  assign n8201 = ( x85 & n8195 ) | ( x85 & ~n8200 ) | ( n8195 & ~n8200 ) ;
  assign n8202 = ( x85 & n7891 ) | ( x85 & ~n8071 ) | ( n7891 & ~n8071 ) ;
  assign n8203 = x85 & n7891 ;
  assign n8204 = ( ~n7896 & n8202 ) | ( ~n7896 & n8203 ) | ( n8202 & n8203 ) ;
  assign n8205 = ( n7896 & n8202 ) | ( n7896 & n8203 ) | ( n8202 & n8203 ) ;
  assign n8206 = ( n7896 & n8204 ) | ( n7896 & ~n8205 ) | ( n8204 & ~n8205 ) ;
  assign n8207 = ( x86 & n8201 ) | ( x86 & ~n8206 ) | ( n8201 & ~n8206 ) ;
  assign n8208 = ( x86 & n7897 ) | ( x86 & ~n8071 ) | ( n7897 & ~n8071 ) ;
  assign n8209 = x86 & n7897 ;
  assign n8210 = ( ~n7902 & n8208 ) | ( ~n7902 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = ( n7902 & n8208 ) | ( n7902 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8212 = ( n7902 & n8210 ) | ( n7902 & ~n8211 ) | ( n8210 & ~n8211 ) ;
  assign n8213 = ( x87 & n8207 ) | ( x87 & ~n8212 ) | ( n8207 & ~n8212 ) ;
  assign n8214 = ( x87 & n7903 ) | ( x87 & ~n8071 ) | ( n7903 & ~n8071 ) ;
  assign n8215 = x87 & n7903 ;
  assign n8216 = ( ~n7908 & n8214 ) | ( ~n7908 & n8215 ) | ( n8214 & n8215 ) ;
  assign n8217 = ( n7908 & n8214 ) | ( n7908 & n8215 ) | ( n8214 & n8215 ) ;
  assign n8218 = ( n7908 & n8216 ) | ( n7908 & ~n8217 ) | ( n8216 & ~n8217 ) ;
  assign n8219 = ( x88 & n8213 ) | ( x88 & ~n8218 ) | ( n8213 & ~n8218 ) ;
  assign n8220 = ( x88 & n7909 ) | ( x88 & ~n8071 ) | ( n7909 & ~n8071 ) ;
  assign n8221 = x88 & n7909 ;
  assign n8222 = ( ~n7914 & n8220 ) | ( ~n7914 & n8221 ) | ( n8220 & n8221 ) ;
  assign n8223 = ( n7914 & n8220 ) | ( n7914 & n8221 ) | ( n8220 & n8221 ) ;
  assign n8224 = ( n7914 & n8222 ) | ( n7914 & ~n8223 ) | ( n8222 & ~n8223 ) ;
  assign n8225 = ( x89 & n8219 ) | ( x89 & ~n8224 ) | ( n8219 & ~n8224 ) ;
  assign n8226 = ( x89 & n7915 ) | ( x89 & ~n8071 ) | ( n7915 & ~n8071 ) ;
  assign n8227 = x89 & n7915 ;
  assign n8228 = ( ~n7920 & n8226 ) | ( ~n7920 & n8227 ) | ( n8226 & n8227 ) ;
  assign n8229 = ( n7920 & n8226 ) | ( n7920 & n8227 ) | ( n8226 & n8227 ) ;
  assign n8230 = ( n7920 & n8228 ) | ( n7920 & ~n8229 ) | ( n8228 & ~n8229 ) ;
  assign n8231 = ( x90 & n8225 ) | ( x90 & ~n8230 ) | ( n8225 & ~n8230 ) ;
  assign n8232 = ( x90 & n7921 ) | ( x90 & ~n8071 ) | ( n7921 & ~n8071 ) ;
  assign n8233 = x90 & n7921 ;
  assign n8234 = ( ~n7926 & n8232 ) | ( ~n7926 & n8233 ) | ( n8232 & n8233 ) ;
  assign n8235 = ( n7926 & n8232 ) | ( n7926 & n8233 ) | ( n8232 & n8233 ) ;
  assign n8236 = ( n7926 & n8234 ) | ( n7926 & ~n8235 ) | ( n8234 & ~n8235 ) ;
  assign n8237 = ( x91 & n8231 ) | ( x91 & ~n8236 ) | ( n8231 & ~n8236 ) ;
  assign n8238 = ( x91 & n7927 ) | ( x91 & ~n8071 ) | ( n7927 & ~n8071 ) ;
  assign n8239 = x91 & n7927 ;
  assign n8240 = ( ~n7932 & n8238 ) | ( ~n7932 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8241 = ( n7932 & n8238 ) | ( n7932 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8242 = ( n7932 & n8240 ) | ( n7932 & ~n8241 ) | ( n8240 & ~n8241 ) ;
  assign n8243 = ( x92 & n8237 ) | ( x92 & ~n8242 ) | ( n8237 & ~n8242 ) ;
  assign n8244 = ( x92 & n7933 ) | ( x92 & ~n8071 ) | ( n7933 & ~n8071 ) ;
  assign n8245 = x92 & n7933 ;
  assign n8246 = ( ~n7938 & n8244 ) | ( ~n7938 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8247 = ( n7938 & n8244 ) | ( n7938 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8248 = ( n7938 & n8246 ) | ( n7938 & ~n8247 ) | ( n8246 & ~n8247 ) ;
  assign n8249 = ( x93 & n8243 ) | ( x93 & ~n8248 ) | ( n8243 & ~n8248 ) ;
  assign n8250 = ( x93 & n7939 ) | ( x93 & ~n8071 ) | ( n7939 & ~n8071 ) ;
  assign n8251 = x93 & n7939 ;
  assign n8252 = ( ~n7944 & n8250 ) | ( ~n7944 & n8251 ) | ( n8250 & n8251 ) ;
  assign n8253 = ( n7944 & n8250 ) | ( n7944 & n8251 ) | ( n8250 & n8251 ) ;
  assign n8254 = ( n7944 & n8252 ) | ( n7944 & ~n8253 ) | ( n8252 & ~n8253 ) ;
  assign n8255 = ( x94 & n8249 ) | ( x94 & ~n8254 ) | ( n8249 & ~n8254 ) ;
  assign n8256 = ( x94 & n7945 ) | ( x94 & ~n8071 ) | ( n7945 & ~n8071 ) ;
  assign n8257 = x94 & n7945 ;
  assign n8258 = ( ~n7950 & n8256 ) | ( ~n7950 & n8257 ) | ( n8256 & n8257 ) ;
  assign n8259 = ( n7950 & n8256 ) | ( n7950 & n8257 ) | ( n8256 & n8257 ) ;
  assign n8260 = ( n7950 & n8258 ) | ( n7950 & ~n8259 ) | ( n8258 & ~n8259 ) ;
  assign n8261 = ( x95 & n8255 ) | ( x95 & ~n8260 ) | ( n8255 & ~n8260 ) ;
  assign n8262 = ( x95 & n7951 ) | ( x95 & ~n8071 ) | ( n7951 & ~n8071 ) ;
  assign n8263 = x95 & n7951 ;
  assign n8264 = ( ~n7956 & n8262 ) | ( ~n7956 & n8263 ) | ( n8262 & n8263 ) ;
  assign n8265 = ( n7956 & n8262 ) | ( n7956 & n8263 ) | ( n8262 & n8263 ) ;
  assign n8266 = ( n7956 & n8264 ) | ( n7956 & ~n8265 ) | ( n8264 & ~n8265 ) ;
  assign n8267 = ( x96 & n8261 ) | ( x96 & ~n8266 ) | ( n8261 & ~n8266 ) ;
  assign n8268 = ( x96 & n7957 ) | ( x96 & ~n8071 ) | ( n7957 & ~n8071 ) ;
  assign n8269 = x96 & n7957 ;
  assign n8270 = ( ~n7962 & n8268 ) | ( ~n7962 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8271 = ( n7962 & n8268 ) | ( n7962 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8272 = ( n7962 & n8270 ) | ( n7962 & ~n8271 ) | ( n8270 & ~n8271 ) ;
  assign n8273 = ( x97 & n8267 ) | ( x97 & ~n8272 ) | ( n8267 & ~n8272 ) ;
  assign n8274 = ( x97 & n7963 ) | ( x97 & ~n8071 ) | ( n7963 & ~n8071 ) ;
  assign n8275 = x97 & n7963 ;
  assign n8276 = ( ~n7968 & n8274 ) | ( ~n7968 & n8275 ) | ( n8274 & n8275 ) ;
  assign n8277 = ( n7968 & n8274 ) | ( n7968 & n8275 ) | ( n8274 & n8275 ) ;
  assign n8278 = ( n7968 & n8276 ) | ( n7968 & ~n8277 ) | ( n8276 & ~n8277 ) ;
  assign n8279 = ( x98 & n8273 ) | ( x98 & ~n8278 ) | ( n8273 & ~n8278 ) ;
  assign n8280 = ( x98 & n7969 ) | ( x98 & ~n8071 ) | ( n7969 & ~n8071 ) ;
  assign n8281 = x98 & n7969 ;
  assign n8282 = ( ~n7974 & n8280 ) | ( ~n7974 & n8281 ) | ( n8280 & n8281 ) ;
  assign n8283 = ( n7974 & n8280 ) | ( n7974 & n8281 ) | ( n8280 & n8281 ) ;
  assign n8284 = ( n7974 & n8282 ) | ( n7974 & ~n8283 ) | ( n8282 & ~n8283 ) ;
  assign n8285 = ( x99 & n8279 ) | ( x99 & ~n8284 ) | ( n8279 & ~n8284 ) ;
  assign n8286 = ( x99 & n7975 ) | ( x99 & ~n8071 ) | ( n7975 & ~n8071 ) ;
  assign n8287 = x99 & n7975 ;
  assign n8288 = ( ~n7980 & n8286 ) | ( ~n7980 & n8287 ) | ( n8286 & n8287 ) ;
  assign n8289 = ( n7980 & n8286 ) | ( n7980 & n8287 ) | ( n8286 & n8287 ) ;
  assign n8290 = ( n7980 & n8288 ) | ( n7980 & ~n8289 ) | ( n8288 & ~n8289 ) ;
  assign n8291 = ( x100 & n8285 ) | ( x100 & ~n8290 ) | ( n8285 & ~n8290 ) ;
  assign n8292 = ( x100 & n7981 ) | ( x100 & ~n8071 ) | ( n7981 & ~n8071 ) ;
  assign n8293 = x100 & n7981 ;
  assign n8294 = ( ~n7986 & n8292 ) | ( ~n7986 & n8293 ) | ( n8292 & n8293 ) ;
  assign n8295 = ( n7986 & n8292 ) | ( n7986 & n8293 ) | ( n8292 & n8293 ) ;
  assign n8296 = ( n7986 & n8294 ) | ( n7986 & ~n8295 ) | ( n8294 & ~n8295 ) ;
  assign n8297 = ( x101 & n8291 ) | ( x101 & ~n8296 ) | ( n8291 & ~n8296 ) ;
  assign n8298 = ( x101 & n7987 ) | ( x101 & ~n8071 ) | ( n7987 & ~n8071 ) ;
  assign n8299 = x101 & n7987 ;
  assign n8300 = ( ~n7992 & n8298 ) | ( ~n7992 & n8299 ) | ( n8298 & n8299 ) ;
  assign n8301 = ( n7992 & n8298 ) | ( n7992 & n8299 ) | ( n8298 & n8299 ) ;
  assign n8302 = ( n7992 & n8300 ) | ( n7992 & ~n8301 ) | ( n8300 & ~n8301 ) ;
  assign n8303 = ( x102 & n8297 ) | ( x102 & ~n8302 ) | ( n8297 & ~n8302 ) ;
  assign n8304 = ( x102 & n7993 ) | ( x102 & ~n8071 ) | ( n7993 & ~n8071 ) ;
  assign n8305 = x102 & n7993 ;
  assign n8306 = ( ~n7998 & n8304 ) | ( ~n7998 & n8305 ) | ( n8304 & n8305 ) ;
  assign n8307 = ( n7998 & n8304 ) | ( n7998 & n8305 ) | ( n8304 & n8305 ) ;
  assign n8308 = ( n7998 & n8306 ) | ( n7998 & ~n8307 ) | ( n8306 & ~n8307 ) ;
  assign n8309 = ( x103 & n8303 ) | ( x103 & ~n8308 ) | ( n8303 & ~n8308 ) ;
  assign n8310 = ( x103 & n7999 ) | ( x103 & ~n8071 ) | ( n7999 & ~n8071 ) ;
  assign n8311 = x103 & n7999 ;
  assign n8312 = ( ~n8004 & n8310 ) | ( ~n8004 & n8311 ) | ( n8310 & n8311 ) ;
  assign n8313 = ( n8004 & n8310 ) | ( n8004 & n8311 ) | ( n8310 & n8311 ) ;
  assign n8314 = ( n8004 & n8312 ) | ( n8004 & ~n8313 ) | ( n8312 & ~n8313 ) ;
  assign n8315 = ( x104 & n8309 ) | ( x104 & ~n8314 ) | ( n8309 & ~n8314 ) ;
  assign n8316 = ( x104 & n8005 ) | ( x104 & ~n8071 ) | ( n8005 & ~n8071 ) ;
  assign n8317 = x104 & n8005 ;
  assign n8318 = ( ~n8010 & n8316 ) | ( ~n8010 & n8317 ) | ( n8316 & n8317 ) ;
  assign n8319 = ( n8010 & n8316 ) | ( n8010 & n8317 ) | ( n8316 & n8317 ) ;
  assign n8320 = ( n8010 & n8318 ) | ( n8010 & ~n8319 ) | ( n8318 & ~n8319 ) ;
  assign n8321 = ( x105 & n8315 ) | ( x105 & ~n8320 ) | ( n8315 & ~n8320 ) ;
  assign n8322 = ( x105 & n8011 ) | ( x105 & ~n8071 ) | ( n8011 & ~n8071 ) ;
  assign n8323 = x105 & n8011 ;
  assign n8324 = ( ~n8016 & n8322 ) | ( ~n8016 & n8323 ) | ( n8322 & n8323 ) ;
  assign n8325 = ( n8016 & n8322 ) | ( n8016 & n8323 ) | ( n8322 & n8323 ) ;
  assign n8326 = ( n8016 & n8324 ) | ( n8016 & ~n8325 ) | ( n8324 & ~n8325 ) ;
  assign n8327 = ( x106 & n8321 ) | ( x106 & ~n8326 ) | ( n8321 & ~n8326 ) ;
  assign n8328 = ( x106 & n8017 ) | ( x106 & ~n8071 ) | ( n8017 & ~n8071 ) ;
  assign n8329 = x106 & n8017 ;
  assign n8330 = ( ~n8022 & n8328 ) | ( ~n8022 & n8329 ) | ( n8328 & n8329 ) ;
  assign n8331 = ( n8022 & n8328 ) | ( n8022 & n8329 ) | ( n8328 & n8329 ) ;
  assign n8332 = ( n8022 & n8330 ) | ( n8022 & ~n8331 ) | ( n8330 & ~n8331 ) ;
  assign n8333 = ( x107 & n8327 ) | ( x107 & ~n8332 ) | ( n8327 & ~n8332 ) ;
  assign n8334 = ( x107 & n8023 ) | ( x107 & ~n8071 ) | ( n8023 & ~n8071 ) ;
  assign n8335 = x107 & n8023 ;
  assign n8336 = ( ~n8028 & n8334 ) | ( ~n8028 & n8335 ) | ( n8334 & n8335 ) ;
  assign n8337 = ( n8028 & n8334 ) | ( n8028 & n8335 ) | ( n8334 & n8335 ) ;
  assign n8338 = ( n8028 & n8336 ) | ( n8028 & ~n8337 ) | ( n8336 & ~n8337 ) ;
  assign n8339 = ( x108 & n8333 ) | ( x108 & ~n8338 ) | ( n8333 & ~n8338 ) ;
  assign n8340 = ( x108 & n8029 ) | ( x108 & ~n8071 ) | ( n8029 & ~n8071 ) ;
  assign n8341 = x108 & n8029 ;
  assign n8342 = ( ~n8034 & n8340 ) | ( ~n8034 & n8341 ) | ( n8340 & n8341 ) ;
  assign n8343 = ( n8034 & n8340 ) | ( n8034 & n8341 ) | ( n8340 & n8341 ) ;
  assign n8344 = ( n8034 & n8342 ) | ( n8034 & ~n8343 ) | ( n8342 & ~n8343 ) ;
  assign n8345 = ( x109 & n8339 ) | ( x109 & ~n8344 ) | ( n8339 & ~n8344 ) ;
  assign n8346 = ( x109 & n8035 ) | ( x109 & ~n8071 ) | ( n8035 & ~n8071 ) ;
  assign n8347 = x109 & n8035 ;
  assign n8348 = ( ~n8040 & n8346 ) | ( ~n8040 & n8347 ) | ( n8346 & n8347 ) ;
  assign n8349 = ( n8040 & n8346 ) | ( n8040 & n8347 ) | ( n8346 & n8347 ) ;
  assign n8350 = ( n8040 & n8348 ) | ( n8040 & ~n8349 ) | ( n8348 & ~n8349 ) ;
  assign n8351 = ( x110 & n8345 ) | ( x110 & ~n8350 ) | ( n8345 & ~n8350 ) ;
  assign n8352 = ( x110 & n8041 ) | ( x110 & ~n8071 ) | ( n8041 & ~n8071 ) ;
  assign n8353 = x110 & n8041 ;
  assign n8354 = ( ~n8046 & n8352 ) | ( ~n8046 & n8353 ) | ( n8352 & n8353 ) ;
  assign n8355 = ( n8046 & n8352 ) | ( n8046 & n8353 ) | ( n8352 & n8353 ) ;
  assign n8356 = ( n8046 & n8354 ) | ( n8046 & ~n8355 ) | ( n8354 & ~n8355 ) ;
  assign n8357 = ( x111 & n8351 ) | ( x111 & ~n8356 ) | ( n8351 & ~n8356 ) ;
  assign n8358 = ( x111 & n8047 ) | ( x111 & ~n8071 ) | ( n8047 & ~n8071 ) ;
  assign n8359 = x111 & n8047 ;
  assign n8360 = ( ~n8052 & n8358 ) | ( ~n8052 & n8359 ) | ( n8358 & n8359 ) ;
  assign n8361 = ( n8052 & n8358 ) | ( n8052 & n8359 ) | ( n8358 & n8359 ) ;
  assign n8362 = ( n8052 & n8360 ) | ( n8052 & ~n8361 ) | ( n8360 & ~n8361 ) ;
  assign n8363 = ( x112 & n8357 ) | ( x112 & ~n8362 ) | ( n8357 & ~n8362 ) ;
  assign n8364 = ( x112 & n8053 ) | ( x112 & ~n8071 ) | ( n8053 & ~n8071 ) ;
  assign n8365 = x112 & n8053 ;
  assign n8366 = ( ~n8058 & n8364 ) | ( ~n8058 & n8365 ) | ( n8364 & n8365 ) ;
  assign n8367 = ( n8058 & n8364 ) | ( n8058 & n8365 ) | ( n8364 & n8365 ) ;
  assign n8368 = ( n8058 & n8366 ) | ( n8058 & ~n8367 ) | ( n8366 & ~n8367 ) ;
  assign n8369 = ( x113 & n8363 ) | ( x113 & ~n8368 ) | ( n8363 & ~n8368 ) ;
  assign n8370 = ( x113 & n8059 ) | ( x113 & ~n8071 ) | ( n8059 & ~n8071 ) ;
  assign n8371 = x113 & n8059 ;
  assign n8372 = ( ~n8064 & n8370 ) | ( ~n8064 & n8371 ) | ( n8370 & n8371 ) ;
  assign n8373 = ( n8064 & n8370 ) | ( n8064 & n8371 ) | ( n8370 & n8371 ) ;
  assign n8374 = ( n8064 & n8372 ) | ( n8064 & ~n8373 ) | ( n8372 & ~n8373 ) ;
  assign n8375 = ( x114 & n8369 ) | ( x114 & ~n8374 ) | ( n8369 & ~n8374 ) ;
  assign n8376 = ( x115 & ~n8076 ) | ( x115 & n8375 ) | ( ~n8076 & n8375 ) ;
  assign n8377 = ( x115 & n141 ) | ( x115 & n8069 ) | ( n141 & n8069 ) ;
  assign n8378 = x115 | n8069 ;
  assign n8379 = ( n8068 & n8377 ) | ( n8068 & ~n8378 ) | ( n8377 & ~n8378 ) ;
  assign n8380 = ( x116 & n8376 ) | ( x116 & ~n8379 ) | ( n8376 & ~n8379 ) ;
  assign n8381 = n140 | n8380 ;
  assign n8382 = ( x115 & n8375 ) | ( x115 & n8381 ) | ( n8375 & n8381 ) ;
  assign n8383 = x115 | n8375 ;
  assign n8384 = ( ~n8076 & n8382 ) | ( ~n8076 & n8383 ) | ( n8382 & n8383 ) ;
  assign n8385 = ( n8076 & n8382 ) | ( n8076 & n8383 ) | ( n8382 & n8383 ) ;
  assign n8386 = ( n8076 & n8384 ) | ( n8076 & ~n8385 ) | ( n8384 & ~n8385 ) ;
  assign n8387 = ~x10 & x64 ;
  assign n8388 = ~x11 & n8381 ;
  assign n8389 = ( x11 & ~x64 ) | ( x11 & n8381 ) | ( ~x64 & n8381 ) ;
  assign n8390 = ( n8077 & ~n8388 ) | ( n8077 & n8389 ) | ( ~n8388 & n8389 ) ;
  assign n8391 = ( x65 & n8387 ) | ( x65 & ~n8390 ) | ( n8387 & ~n8390 ) ;
  assign n8392 = ( x65 & n8077 ) | ( x65 & n8381 ) | ( n8077 & n8381 ) ;
  assign n8393 = x65 | n8077 ;
  assign n8394 = ( ~n8080 & n8392 ) | ( ~n8080 & n8393 ) | ( n8392 & n8393 ) ;
  assign n8395 = ( n8080 & n8392 ) | ( n8080 & n8393 ) | ( n8392 & n8393 ) ;
  assign n8396 = ( n8080 & n8394 ) | ( n8080 & ~n8395 ) | ( n8394 & ~n8395 ) ;
  assign n8397 = ( x66 & n8391 ) | ( x66 & ~n8396 ) | ( n8391 & ~n8396 ) ;
  assign n8398 = ( x66 & n8081 ) | ( x66 & n8381 ) | ( n8081 & n8381 ) ;
  assign n8399 = x66 | n8081 ;
  assign n8400 = ( ~n8086 & n8398 ) | ( ~n8086 & n8399 ) | ( n8398 & n8399 ) ;
  assign n8401 = ( n8086 & n8398 ) | ( n8086 & n8399 ) | ( n8398 & n8399 ) ;
  assign n8402 = ( n8086 & n8400 ) | ( n8086 & ~n8401 ) | ( n8400 & ~n8401 ) ;
  assign n8403 = ( x67 & n8397 ) | ( x67 & ~n8402 ) | ( n8397 & ~n8402 ) ;
  assign n8404 = ( x67 & n8087 ) | ( x67 & ~n8381 ) | ( n8087 & ~n8381 ) ;
  assign n8405 = x67 & n8087 ;
  assign n8406 = ( ~n8092 & n8404 ) | ( ~n8092 & n8405 ) | ( n8404 & n8405 ) ;
  assign n8407 = ( n8092 & n8404 ) | ( n8092 & n8405 ) | ( n8404 & n8405 ) ;
  assign n8408 = ( n8092 & n8406 ) | ( n8092 & ~n8407 ) | ( n8406 & ~n8407 ) ;
  assign n8409 = ( x68 & n8403 ) | ( x68 & ~n8408 ) | ( n8403 & ~n8408 ) ;
  assign n8410 = ( x68 & n8093 ) | ( x68 & ~n8381 ) | ( n8093 & ~n8381 ) ;
  assign n8411 = x68 & n8093 ;
  assign n8412 = ( ~n8098 & n8410 ) | ( ~n8098 & n8411 ) | ( n8410 & n8411 ) ;
  assign n8413 = ( n8098 & n8410 ) | ( n8098 & n8411 ) | ( n8410 & n8411 ) ;
  assign n8414 = ( n8098 & n8412 ) | ( n8098 & ~n8413 ) | ( n8412 & ~n8413 ) ;
  assign n8415 = ( x69 & n8409 ) | ( x69 & ~n8414 ) | ( n8409 & ~n8414 ) ;
  assign n8416 = ( x69 & n8099 ) | ( x69 & ~n8381 ) | ( n8099 & ~n8381 ) ;
  assign n8417 = x69 & n8099 ;
  assign n8418 = ( ~n8104 & n8416 ) | ( ~n8104 & n8417 ) | ( n8416 & n8417 ) ;
  assign n8419 = ( n8104 & n8416 ) | ( n8104 & n8417 ) | ( n8416 & n8417 ) ;
  assign n8420 = ( n8104 & n8418 ) | ( n8104 & ~n8419 ) | ( n8418 & ~n8419 ) ;
  assign n8421 = ( x70 & n8415 ) | ( x70 & ~n8420 ) | ( n8415 & ~n8420 ) ;
  assign n8422 = ( x70 & n8105 ) | ( x70 & ~n8381 ) | ( n8105 & ~n8381 ) ;
  assign n8423 = x70 & n8105 ;
  assign n8424 = ( ~n8110 & n8422 ) | ( ~n8110 & n8423 ) | ( n8422 & n8423 ) ;
  assign n8425 = ( n8110 & n8422 ) | ( n8110 & n8423 ) | ( n8422 & n8423 ) ;
  assign n8426 = ( n8110 & n8424 ) | ( n8110 & ~n8425 ) | ( n8424 & ~n8425 ) ;
  assign n8427 = ( x71 & n8421 ) | ( x71 & ~n8426 ) | ( n8421 & ~n8426 ) ;
  assign n8428 = ( x71 & n8111 ) | ( x71 & ~n8381 ) | ( n8111 & ~n8381 ) ;
  assign n8429 = x71 & n8111 ;
  assign n8430 = ( ~n8116 & n8428 ) | ( ~n8116 & n8429 ) | ( n8428 & n8429 ) ;
  assign n8431 = ( n8116 & n8428 ) | ( n8116 & n8429 ) | ( n8428 & n8429 ) ;
  assign n8432 = ( n8116 & n8430 ) | ( n8116 & ~n8431 ) | ( n8430 & ~n8431 ) ;
  assign n8433 = ( x72 & n8427 ) | ( x72 & ~n8432 ) | ( n8427 & ~n8432 ) ;
  assign n8434 = ( x72 & n8117 ) | ( x72 & ~n8381 ) | ( n8117 & ~n8381 ) ;
  assign n8435 = x72 & n8117 ;
  assign n8436 = ( ~n8122 & n8434 ) | ( ~n8122 & n8435 ) | ( n8434 & n8435 ) ;
  assign n8437 = ( n8122 & n8434 ) | ( n8122 & n8435 ) | ( n8434 & n8435 ) ;
  assign n8438 = ( n8122 & n8436 ) | ( n8122 & ~n8437 ) | ( n8436 & ~n8437 ) ;
  assign n8439 = ( x73 & n8433 ) | ( x73 & ~n8438 ) | ( n8433 & ~n8438 ) ;
  assign n8440 = ( x73 & n8123 ) | ( x73 & ~n8381 ) | ( n8123 & ~n8381 ) ;
  assign n8441 = x73 & n8123 ;
  assign n8442 = ( ~n8128 & n8440 ) | ( ~n8128 & n8441 ) | ( n8440 & n8441 ) ;
  assign n8443 = ( n8128 & n8440 ) | ( n8128 & n8441 ) | ( n8440 & n8441 ) ;
  assign n8444 = ( n8128 & n8442 ) | ( n8128 & ~n8443 ) | ( n8442 & ~n8443 ) ;
  assign n8445 = ( x74 & n8439 ) | ( x74 & ~n8444 ) | ( n8439 & ~n8444 ) ;
  assign n8446 = ( x74 & n8129 ) | ( x74 & ~n8381 ) | ( n8129 & ~n8381 ) ;
  assign n8447 = x74 & n8129 ;
  assign n8448 = ( ~n8134 & n8446 ) | ( ~n8134 & n8447 ) | ( n8446 & n8447 ) ;
  assign n8449 = ( n8134 & n8446 ) | ( n8134 & n8447 ) | ( n8446 & n8447 ) ;
  assign n8450 = ( n8134 & n8448 ) | ( n8134 & ~n8449 ) | ( n8448 & ~n8449 ) ;
  assign n8451 = ( x75 & n8445 ) | ( x75 & ~n8450 ) | ( n8445 & ~n8450 ) ;
  assign n8452 = ( x75 & n8135 ) | ( x75 & ~n8381 ) | ( n8135 & ~n8381 ) ;
  assign n8453 = x75 & n8135 ;
  assign n8454 = ( ~n8140 & n8452 ) | ( ~n8140 & n8453 ) | ( n8452 & n8453 ) ;
  assign n8455 = ( n8140 & n8452 ) | ( n8140 & n8453 ) | ( n8452 & n8453 ) ;
  assign n8456 = ( n8140 & n8454 ) | ( n8140 & ~n8455 ) | ( n8454 & ~n8455 ) ;
  assign n8457 = ( x76 & n8451 ) | ( x76 & ~n8456 ) | ( n8451 & ~n8456 ) ;
  assign n8458 = ( x76 & n8141 ) | ( x76 & ~n8381 ) | ( n8141 & ~n8381 ) ;
  assign n8459 = x76 & n8141 ;
  assign n8460 = ( ~n8146 & n8458 ) | ( ~n8146 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8461 = ( n8146 & n8458 ) | ( n8146 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8462 = ( n8146 & n8460 ) | ( n8146 & ~n8461 ) | ( n8460 & ~n8461 ) ;
  assign n8463 = ( x77 & n8457 ) | ( x77 & ~n8462 ) | ( n8457 & ~n8462 ) ;
  assign n8464 = ( x77 & n8147 ) | ( x77 & ~n8381 ) | ( n8147 & ~n8381 ) ;
  assign n8465 = x77 & n8147 ;
  assign n8466 = ( ~n8152 & n8464 ) | ( ~n8152 & n8465 ) | ( n8464 & n8465 ) ;
  assign n8467 = ( n8152 & n8464 ) | ( n8152 & n8465 ) | ( n8464 & n8465 ) ;
  assign n8468 = ( n8152 & n8466 ) | ( n8152 & ~n8467 ) | ( n8466 & ~n8467 ) ;
  assign n8469 = ( x78 & n8463 ) | ( x78 & ~n8468 ) | ( n8463 & ~n8468 ) ;
  assign n8470 = ( x78 & n8153 ) | ( x78 & ~n8381 ) | ( n8153 & ~n8381 ) ;
  assign n8471 = x78 & n8153 ;
  assign n8472 = ( ~n8158 & n8470 ) | ( ~n8158 & n8471 ) | ( n8470 & n8471 ) ;
  assign n8473 = ( n8158 & n8470 ) | ( n8158 & n8471 ) | ( n8470 & n8471 ) ;
  assign n8474 = ( n8158 & n8472 ) | ( n8158 & ~n8473 ) | ( n8472 & ~n8473 ) ;
  assign n8475 = ( x79 & n8469 ) | ( x79 & ~n8474 ) | ( n8469 & ~n8474 ) ;
  assign n8476 = ( x79 & n8159 ) | ( x79 & ~n8381 ) | ( n8159 & ~n8381 ) ;
  assign n8477 = x79 & n8159 ;
  assign n8478 = ( ~n8164 & n8476 ) | ( ~n8164 & n8477 ) | ( n8476 & n8477 ) ;
  assign n8479 = ( n8164 & n8476 ) | ( n8164 & n8477 ) | ( n8476 & n8477 ) ;
  assign n8480 = ( n8164 & n8478 ) | ( n8164 & ~n8479 ) | ( n8478 & ~n8479 ) ;
  assign n8481 = ( x80 & n8475 ) | ( x80 & ~n8480 ) | ( n8475 & ~n8480 ) ;
  assign n8482 = ( x80 & n8165 ) | ( x80 & ~n8381 ) | ( n8165 & ~n8381 ) ;
  assign n8483 = x80 & n8165 ;
  assign n8484 = ( ~n8170 & n8482 ) | ( ~n8170 & n8483 ) | ( n8482 & n8483 ) ;
  assign n8485 = ( n8170 & n8482 ) | ( n8170 & n8483 ) | ( n8482 & n8483 ) ;
  assign n8486 = ( n8170 & n8484 ) | ( n8170 & ~n8485 ) | ( n8484 & ~n8485 ) ;
  assign n8487 = ( x81 & n8481 ) | ( x81 & ~n8486 ) | ( n8481 & ~n8486 ) ;
  assign n8488 = ( x81 & n8171 ) | ( x81 & ~n8381 ) | ( n8171 & ~n8381 ) ;
  assign n8489 = x81 & n8171 ;
  assign n8490 = ( ~n8176 & n8488 ) | ( ~n8176 & n8489 ) | ( n8488 & n8489 ) ;
  assign n8491 = ( n8176 & n8488 ) | ( n8176 & n8489 ) | ( n8488 & n8489 ) ;
  assign n8492 = ( n8176 & n8490 ) | ( n8176 & ~n8491 ) | ( n8490 & ~n8491 ) ;
  assign n8493 = ( x82 & n8487 ) | ( x82 & ~n8492 ) | ( n8487 & ~n8492 ) ;
  assign n8494 = ( x82 & n8177 ) | ( x82 & ~n8381 ) | ( n8177 & ~n8381 ) ;
  assign n8495 = x82 & n8177 ;
  assign n8496 = ( ~n8182 & n8494 ) | ( ~n8182 & n8495 ) | ( n8494 & n8495 ) ;
  assign n8497 = ( n8182 & n8494 ) | ( n8182 & n8495 ) | ( n8494 & n8495 ) ;
  assign n8498 = ( n8182 & n8496 ) | ( n8182 & ~n8497 ) | ( n8496 & ~n8497 ) ;
  assign n8499 = ( x83 & n8493 ) | ( x83 & ~n8498 ) | ( n8493 & ~n8498 ) ;
  assign n8500 = ( x83 & n8183 ) | ( x83 & ~n8381 ) | ( n8183 & ~n8381 ) ;
  assign n8501 = x83 & n8183 ;
  assign n8502 = ( ~n8188 & n8500 ) | ( ~n8188 & n8501 ) | ( n8500 & n8501 ) ;
  assign n8503 = ( n8188 & n8500 ) | ( n8188 & n8501 ) | ( n8500 & n8501 ) ;
  assign n8504 = ( n8188 & n8502 ) | ( n8188 & ~n8503 ) | ( n8502 & ~n8503 ) ;
  assign n8505 = ( x84 & n8499 ) | ( x84 & ~n8504 ) | ( n8499 & ~n8504 ) ;
  assign n8506 = ( x84 & n8189 ) | ( x84 & ~n8381 ) | ( n8189 & ~n8381 ) ;
  assign n8507 = x84 & n8189 ;
  assign n8508 = ( ~n8194 & n8506 ) | ( ~n8194 & n8507 ) | ( n8506 & n8507 ) ;
  assign n8509 = ( n8194 & n8506 ) | ( n8194 & n8507 ) | ( n8506 & n8507 ) ;
  assign n8510 = ( n8194 & n8508 ) | ( n8194 & ~n8509 ) | ( n8508 & ~n8509 ) ;
  assign n8511 = ( x85 & n8505 ) | ( x85 & ~n8510 ) | ( n8505 & ~n8510 ) ;
  assign n8512 = ( x85 & n8195 ) | ( x85 & ~n8381 ) | ( n8195 & ~n8381 ) ;
  assign n8513 = x85 & n8195 ;
  assign n8514 = ( ~n8200 & n8512 ) | ( ~n8200 & n8513 ) | ( n8512 & n8513 ) ;
  assign n8515 = ( n8200 & n8512 ) | ( n8200 & n8513 ) | ( n8512 & n8513 ) ;
  assign n8516 = ( n8200 & n8514 ) | ( n8200 & ~n8515 ) | ( n8514 & ~n8515 ) ;
  assign n8517 = ( x86 & n8511 ) | ( x86 & ~n8516 ) | ( n8511 & ~n8516 ) ;
  assign n8518 = ( x86 & n8201 ) | ( x86 & ~n8381 ) | ( n8201 & ~n8381 ) ;
  assign n8519 = x86 & n8201 ;
  assign n8520 = ( ~n8206 & n8518 ) | ( ~n8206 & n8519 ) | ( n8518 & n8519 ) ;
  assign n8521 = ( n8206 & n8518 ) | ( n8206 & n8519 ) | ( n8518 & n8519 ) ;
  assign n8522 = ( n8206 & n8520 ) | ( n8206 & ~n8521 ) | ( n8520 & ~n8521 ) ;
  assign n8523 = ( x87 & n8517 ) | ( x87 & ~n8522 ) | ( n8517 & ~n8522 ) ;
  assign n8524 = ( x87 & n8207 ) | ( x87 & ~n8381 ) | ( n8207 & ~n8381 ) ;
  assign n8525 = x87 & n8207 ;
  assign n8526 = ( ~n8212 & n8524 ) | ( ~n8212 & n8525 ) | ( n8524 & n8525 ) ;
  assign n8527 = ( n8212 & n8524 ) | ( n8212 & n8525 ) | ( n8524 & n8525 ) ;
  assign n8528 = ( n8212 & n8526 ) | ( n8212 & ~n8527 ) | ( n8526 & ~n8527 ) ;
  assign n8529 = ( x88 & n8523 ) | ( x88 & ~n8528 ) | ( n8523 & ~n8528 ) ;
  assign n8530 = ( x88 & n8213 ) | ( x88 & ~n8381 ) | ( n8213 & ~n8381 ) ;
  assign n8531 = x88 & n8213 ;
  assign n8532 = ( ~n8218 & n8530 ) | ( ~n8218 & n8531 ) | ( n8530 & n8531 ) ;
  assign n8533 = ( n8218 & n8530 ) | ( n8218 & n8531 ) | ( n8530 & n8531 ) ;
  assign n8534 = ( n8218 & n8532 ) | ( n8218 & ~n8533 ) | ( n8532 & ~n8533 ) ;
  assign n8535 = ( x89 & n8529 ) | ( x89 & ~n8534 ) | ( n8529 & ~n8534 ) ;
  assign n8536 = ( x89 & n8219 ) | ( x89 & ~n8381 ) | ( n8219 & ~n8381 ) ;
  assign n8537 = x89 & n8219 ;
  assign n8538 = ( ~n8224 & n8536 ) | ( ~n8224 & n8537 ) | ( n8536 & n8537 ) ;
  assign n8539 = ( n8224 & n8536 ) | ( n8224 & n8537 ) | ( n8536 & n8537 ) ;
  assign n8540 = ( n8224 & n8538 ) | ( n8224 & ~n8539 ) | ( n8538 & ~n8539 ) ;
  assign n8541 = ( x90 & n8535 ) | ( x90 & ~n8540 ) | ( n8535 & ~n8540 ) ;
  assign n8542 = ( x90 & n8225 ) | ( x90 & ~n8381 ) | ( n8225 & ~n8381 ) ;
  assign n8543 = x90 & n8225 ;
  assign n8544 = ( ~n8230 & n8542 ) | ( ~n8230 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8545 = ( n8230 & n8542 ) | ( n8230 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8546 = ( n8230 & n8544 ) | ( n8230 & ~n8545 ) | ( n8544 & ~n8545 ) ;
  assign n8547 = ( x91 & n8541 ) | ( x91 & ~n8546 ) | ( n8541 & ~n8546 ) ;
  assign n8548 = ( x91 & n8231 ) | ( x91 & ~n8381 ) | ( n8231 & ~n8381 ) ;
  assign n8549 = x91 & n8231 ;
  assign n8550 = ( ~n8236 & n8548 ) | ( ~n8236 & n8549 ) | ( n8548 & n8549 ) ;
  assign n8551 = ( n8236 & n8548 ) | ( n8236 & n8549 ) | ( n8548 & n8549 ) ;
  assign n8552 = ( n8236 & n8550 ) | ( n8236 & ~n8551 ) | ( n8550 & ~n8551 ) ;
  assign n8553 = ( x92 & n8547 ) | ( x92 & ~n8552 ) | ( n8547 & ~n8552 ) ;
  assign n8554 = ( x92 & n8237 ) | ( x92 & ~n8381 ) | ( n8237 & ~n8381 ) ;
  assign n8555 = x92 & n8237 ;
  assign n8556 = ( ~n8242 & n8554 ) | ( ~n8242 & n8555 ) | ( n8554 & n8555 ) ;
  assign n8557 = ( n8242 & n8554 ) | ( n8242 & n8555 ) | ( n8554 & n8555 ) ;
  assign n8558 = ( n8242 & n8556 ) | ( n8242 & ~n8557 ) | ( n8556 & ~n8557 ) ;
  assign n8559 = ( x93 & n8553 ) | ( x93 & ~n8558 ) | ( n8553 & ~n8558 ) ;
  assign n8560 = ( x93 & n8243 ) | ( x93 & ~n8381 ) | ( n8243 & ~n8381 ) ;
  assign n8561 = x93 & n8243 ;
  assign n8562 = ( ~n8248 & n8560 ) | ( ~n8248 & n8561 ) | ( n8560 & n8561 ) ;
  assign n8563 = ( n8248 & n8560 ) | ( n8248 & n8561 ) | ( n8560 & n8561 ) ;
  assign n8564 = ( n8248 & n8562 ) | ( n8248 & ~n8563 ) | ( n8562 & ~n8563 ) ;
  assign n8565 = ( x94 & n8559 ) | ( x94 & ~n8564 ) | ( n8559 & ~n8564 ) ;
  assign n8566 = ( x94 & n8249 ) | ( x94 & ~n8381 ) | ( n8249 & ~n8381 ) ;
  assign n8567 = x94 & n8249 ;
  assign n8568 = ( ~n8254 & n8566 ) | ( ~n8254 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = ( n8254 & n8566 ) | ( n8254 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8570 = ( n8254 & n8568 ) | ( n8254 & ~n8569 ) | ( n8568 & ~n8569 ) ;
  assign n8571 = ( x95 & n8565 ) | ( x95 & ~n8570 ) | ( n8565 & ~n8570 ) ;
  assign n8572 = ( x95 & n8255 ) | ( x95 & ~n8381 ) | ( n8255 & ~n8381 ) ;
  assign n8573 = x95 & n8255 ;
  assign n8574 = ( ~n8260 & n8572 ) | ( ~n8260 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8575 = ( n8260 & n8572 ) | ( n8260 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8576 = ( n8260 & n8574 ) | ( n8260 & ~n8575 ) | ( n8574 & ~n8575 ) ;
  assign n8577 = ( x96 & n8571 ) | ( x96 & ~n8576 ) | ( n8571 & ~n8576 ) ;
  assign n8578 = ( x96 & n8261 ) | ( x96 & ~n8381 ) | ( n8261 & ~n8381 ) ;
  assign n8579 = x96 & n8261 ;
  assign n8580 = ( ~n8266 & n8578 ) | ( ~n8266 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = ( n8266 & n8578 ) | ( n8266 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8582 = ( n8266 & n8580 ) | ( n8266 & ~n8581 ) | ( n8580 & ~n8581 ) ;
  assign n8583 = ( x97 & n8577 ) | ( x97 & ~n8582 ) | ( n8577 & ~n8582 ) ;
  assign n8584 = ( x97 & n8267 ) | ( x97 & ~n8381 ) | ( n8267 & ~n8381 ) ;
  assign n8585 = x97 & n8267 ;
  assign n8586 = ( ~n8272 & n8584 ) | ( ~n8272 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8587 = ( n8272 & n8584 ) | ( n8272 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8588 = ( n8272 & n8586 ) | ( n8272 & ~n8587 ) | ( n8586 & ~n8587 ) ;
  assign n8589 = ( x98 & n8583 ) | ( x98 & ~n8588 ) | ( n8583 & ~n8588 ) ;
  assign n8590 = ( x98 & n8273 ) | ( x98 & ~n8381 ) | ( n8273 & ~n8381 ) ;
  assign n8591 = x98 & n8273 ;
  assign n8592 = ( ~n8278 & n8590 ) | ( ~n8278 & n8591 ) | ( n8590 & n8591 ) ;
  assign n8593 = ( n8278 & n8590 ) | ( n8278 & n8591 ) | ( n8590 & n8591 ) ;
  assign n8594 = ( n8278 & n8592 ) | ( n8278 & ~n8593 ) | ( n8592 & ~n8593 ) ;
  assign n8595 = ( x99 & n8589 ) | ( x99 & ~n8594 ) | ( n8589 & ~n8594 ) ;
  assign n8596 = ( x99 & n8279 ) | ( x99 & ~n8381 ) | ( n8279 & ~n8381 ) ;
  assign n8597 = x99 & n8279 ;
  assign n8598 = ( ~n8284 & n8596 ) | ( ~n8284 & n8597 ) | ( n8596 & n8597 ) ;
  assign n8599 = ( n8284 & n8596 ) | ( n8284 & n8597 ) | ( n8596 & n8597 ) ;
  assign n8600 = ( n8284 & n8598 ) | ( n8284 & ~n8599 ) | ( n8598 & ~n8599 ) ;
  assign n8601 = ( x100 & n8595 ) | ( x100 & ~n8600 ) | ( n8595 & ~n8600 ) ;
  assign n8602 = ( x100 & n8285 ) | ( x100 & ~n8381 ) | ( n8285 & ~n8381 ) ;
  assign n8603 = x100 & n8285 ;
  assign n8604 = ( ~n8290 & n8602 ) | ( ~n8290 & n8603 ) | ( n8602 & n8603 ) ;
  assign n8605 = ( n8290 & n8602 ) | ( n8290 & n8603 ) | ( n8602 & n8603 ) ;
  assign n8606 = ( n8290 & n8604 ) | ( n8290 & ~n8605 ) | ( n8604 & ~n8605 ) ;
  assign n8607 = ( x101 & n8601 ) | ( x101 & ~n8606 ) | ( n8601 & ~n8606 ) ;
  assign n8608 = ( x101 & n8291 ) | ( x101 & ~n8381 ) | ( n8291 & ~n8381 ) ;
  assign n8609 = x101 & n8291 ;
  assign n8610 = ( ~n8296 & n8608 ) | ( ~n8296 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = ( n8296 & n8608 ) | ( n8296 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8612 = ( n8296 & n8610 ) | ( n8296 & ~n8611 ) | ( n8610 & ~n8611 ) ;
  assign n8613 = ( x102 & n8607 ) | ( x102 & ~n8612 ) | ( n8607 & ~n8612 ) ;
  assign n8614 = ( x102 & n8297 ) | ( x102 & ~n8381 ) | ( n8297 & ~n8381 ) ;
  assign n8615 = x102 & n8297 ;
  assign n8616 = ( ~n8302 & n8614 ) | ( ~n8302 & n8615 ) | ( n8614 & n8615 ) ;
  assign n8617 = ( n8302 & n8614 ) | ( n8302 & n8615 ) | ( n8614 & n8615 ) ;
  assign n8618 = ( n8302 & n8616 ) | ( n8302 & ~n8617 ) | ( n8616 & ~n8617 ) ;
  assign n8619 = ( x103 & n8613 ) | ( x103 & ~n8618 ) | ( n8613 & ~n8618 ) ;
  assign n8620 = ( x103 & n8303 ) | ( x103 & ~n8381 ) | ( n8303 & ~n8381 ) ;
  assign n8621 = x103 & n8303 ;
  assign n8622 = ( ~n8308 & n8620 ) | ( ~n8308 & n8621 ) | ( n8620 & n8621 ) ;
  assign n8623 = ( n8308 & n8620 ) | ( n8308 & n8621 ) | ( n8620 & n8621 ) ;
  assign n8624 = ( n8308 & n8622 ) | ( n8308 & ~n8623 ) | ( n8622 & ~n8623 ) ;
  assign n8625 = ( x104 & n8619 ) | ( x104 & ~n8624 ) | ( n8619 & ~n8624 ) ;
  assign n8626 = ( x104 & n8309 ) | ( x104 & ~n8381 ) | ( n8309 & ~n8381 ) ;
  assign n8627 = x104 & n8309 ;
  assign n8628 = ( ~n8314 & n8626 ) | ( ~n8314 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8629 = ( n8314 & n8626 ) | ( n8314 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8630 = ( n8314 & n8628 ) | ( n8314 & ~n8629 ) | ( n8628 & ~n8629 ) ;
  assign n8631 = ( x105 & n8625 ) | ( x105 & ~n8630 ) | ( n8625 & ~n8630 ) ;
  assign n8632 = ( x105 & n8315 ) | ( x105 & ~n8381 ) | ( n8315 & ~n8381 ) ;
  assign n8633 = x105 & n8315 ;
  assign n8634 = ( ~n8320 & n8632 ) | ( ~n8320 & n8633 ) | ( n8632 & n8633 ) ;
  assign n8635 = ( n8320 & n8632 ) | ( n8320 & n8633 ) | ( n8632 & n8633 ) ;
  assign n8636 = ( n8320 & n8634 ) | ( n8320 & ~n8635 ) | ( n8634 & ~n8635 ) ;
  assign n8637 = ( x106 & n8631 ) | ( x106 & ~n8636 ) | ( n8631 & ~n8636 ) ;
  assign n8638 = ( x106 & n8321 ) | ( x106 & ~n8381 ) | ( n8321 & ~n8381 ) ;
  assign n8639 = x106 & n8321 ;
  assign n8640 = ( ~n8326 & n8638 ) | ( ~n8326 & n8639 ) | ( n8638 & n8639 ) ;
  assign n8641 = ( n8326 & n8638 ) | ( n8326 & n8639 ) | ( n8638 & n8639 ) ;
  assign n8642 = ( n8326 & n8640 ) | ( n8326 & ~n8641 ) | ( n8640 & ~n8641 ) ;
  assign n8643 = ( x107 & n8637 ) | ( x107 & ~n8642 ) | ( n8637 & ~n8642 ) ;
  assign n8644 = ( x107 & n8327 ) | ( x107 & ~n8381 ) | ( n8327 & ~n8381 ) ;
  assign n8645 = x107 & n8327 ;
  assign n8646 = ( ~n8332 & n8644 ) | ( ~n8332 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = ( n8332 & n8644 ) | ( n8332 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8648 = ( n8332 & n8646 ) | ( n8332 & ~n8647 ) | ( n8646 & ~n8647 ) ;
  assign n8649 = ( x108 & n8643 ) | ( x108 & ~n8648 ) | ( n8643 & ~n8648 ) ;
  assign n8650 = ( x108 & n8333 ) | ( x108 & ~n8381 ) | ( n8333 & ~n8381 ) ;
  assign n8651 = x108 & n8333 ;
  assign n8652 = ( ~n8338 & n8650 ) | ( ~n8338 & n8651 ) | ( n8650 & n8651 ) ;
  assign n8653 = ( n8338 & n8650 ) | ( n8338 & n8651 ) | ( n8650 & n8651 ) ;
  assign n8654 = ( n8338 & n8652 ) | ( n8338 & ~n8653 ) | ( n8652 & ~n8653 ) ;
  assign n8655 = ( x109 & n8649 ) | ( x109 & ~n8654 ) | ( n8649 & ~n8654 ) ;
  assign n8656 = ( x109 & n8339 ) | ( x109 & ~n8381 ) | ( n8339 & ~n8381 ) ;
  assign n8657 = x109 & n8339 ;
  assign n8658 = ( ~n8344 & n8656 ) | ( ~n8344 & n8657 ) | ( n8656 & n8657 ) ;
  assign n8659 = ( n8344 & n8656 ) | ( n8344 & n8657 ) | ( n8656 & n8657 ) ;
  assign n8660 = ( n8344 & n8658 ) | ( n8344 & ~n8659 ) | ( n8658 & ~n8659 ) ;
  assign n8661 = ( x110 & n8655 ) | ( x110 & ~n8660 ) | ( n8655 & ~n8660 ) ;
  assign n8662 = ( x110 & n8345 ) | ( x110 & ~n8381 ) | ( n8345 & ~n8381 ) ;
  assign n8663 = x110 & n8345 ;
  assign n8664 = ( ~n8350 & n8662 ) | ( ~n8350 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8665 = ( n8350 & n8662 ) | ( n8350 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8666 = ( n8350 & n8664 ) | ( n8350 & ~n8665 ) | ( n8664 & ~n8665 ) ;
  assign n8667 = ( x111 & n8661 ) | ( x111 & ~n8666 ) | ( n8661 & ~n8666 ) ;
  assign n8668 = ( x111 & n8351 ) | ( x111 & ~n8381 ) | ( n8351 & ~n8381 ) ;
  assign n8669 = x111 & n8351 ;
  assign n8670 = ( ~n8356 & n8668 ) | ( ~n8356 & n8669 ) | ( n8668 & n8669 ) ;
  assign n8671 = ( n8356 & n8668 ) | ( n8356 & n8669 ) | ( n8668 & n8669 ) ;
  assign n8672 = ( n8356 & n8670 ) | ( n8356 & ~n8671 ) | ( n8670 & ~n8671 ) ;
  assign n8673 = ( x112 & n8667 ) | ( x112 & ~n8672 ) | ( n8667 & ~n8672 ) ;
  assign n8674 = ( x112 & n8357 ) | ( x112 & ~n8381 ) | ( n8357 & ~n8381 ) ;
  assign n8675 = x112 & n8357 ;
  assign n8676 = ( ~n8362 & n8674 ) | ( ~n8362 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8677 = ( n8362 & n8674 ) | ( n8362 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8678 = ( n8362 & n8676 ) | ( n8362 & ~n8677 ) | ( n8676 & ~n8677 ) ;
  assign n8679 = ( x113 & n8673 ) | ( x113 & ~n8678 ) | ( n8673 & ~n8678 ) ;
  assign n8680 = ( x113 & n8363 ) | ( x113 & ~n8381 ) | ( n8363 & ~n8381 ) ;
  assign n8681 = x113 & n8363 ;
  assign n8682 = ( ~n8368 & n8680 ) | ( ~n8368 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8683 = ( n8368 & n8680 ) | ( n8368 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8684 = ( n8368 & n8682 ) | ( n8368 & ~n8683 ) | ( n8682 & ~n8683 ) ;
  assign n8685 = ( x114 & n8679 ) | ( x114 & ~n8684 ) | ( n8679 & ~n8684 ) ;
  assign n8686 = ( x114 & n8369 ) | ( x114 & ~n8381 ) | ( n8369 & ~n8381 ) ;
  assign n8687 = x114 & n8369 ;
  assign n8688 = ( ~n8374 & n8686 ) | ( ~n8374 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8689 = ( n8374 & n8686 ) | ( n8374 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8690 = ( n8374 & n8688 ) | ( n8374 & ~n8689 ) | ( n8688 & ~n8689 ) ;
  assign n8691 = ( x115 & n8685 ) | ( x115 & ~n8690 ) | ( n8685 & ~n8690 ) ;
  assign n8692 = ( x116 & ~n8386 ) | ( x116 & n8691 ) | ( ~n8386 & n8691 ) ;
  assign n8693 = ( n140 & n141 ) | ( n140 & n8376 ) | ( n141 & n8376 ) ;
  assign n8694 = n8068 & n8693 ;
  assign n8695 = n389 | n8694 ;
  assign n8696 = ( x117 & n8692 ) | ( x117 & ~n8695 ) | ( n8692 & ~n8695 ) ;
  assign n8697 = n139 | n8696 ;
  assign n8698 = ( x116 & n8691 ) | ( x116 & n8697 ) | ( n8691 & n8697 ) ;
  assign n8699 = x116 | n8691 ;
  assign n8700 = ( ~n8386 & n8698 ) | ( ~n8386 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8701 = ( n8386 & n8698 ) | ( n8386 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8702 = ( n8386 & n8700 ) | ( n8386 & ~n8701 ) | ( n8700 & ~n8701 ) ;
  assign n8703 = ~x9 & x64 ;
  assign n8704 = ~x10 & n8697 ;
  assign n8705 = ( x10 & ~x64 ) | ( x10 & n8697 ) | ( ~x64 & n8697 ) ;
  assign n8706 = ( n8387 & ~n8704 ) | ( n8387 & n8705 ) | ( ~n8704 & n8705 ) ;
  assign n8707 = ( x65 & n8703 ) | ( x65 & ~n8706 ) | ( n8703 & ~n8706 ) ;
  assign n8708 = ( x65 & n8387 ) | ( x65 & n8697 ) | ( n8387 & n8697 ) ;
  assign n8709 = x65 | n8387 ;
  assign n8710 = ( ~n8390 & n8708 ) | ( ~n8390 & n8709 ) | ( n8708 & n8709 ) ;
  assign n8711 = ( n8390 & n8708 ) | ( n8390 & n8709 ) | ( n8708 & n8709 ) ;
  assign n8712 = ( n8390 & n8710 ) | ( n8390 & ~n8711 ) | ( n8710 & ~n8711 ) ;
  assign n8713 = ( x66 & n8707 ) | ( x66 & ~n8712 ) | ( n8707 & ~n8712 ) ;
  assign n8714 = ( x66 & n8391 ) | ( x66 & n8697 ) | ( n8391 & n8697 ) ;
  assign n8715 = x66 | n8391 ;
  assign n8716 = ( ~n8396 & n8714 ) | ( ~n8396 & n8715 ) | ( n8714 & n8715 ) ;
  assign n8717 = ( n8396 & n8714 ) | ( n8396 & n8715 ) | ( n8714 & n8715 ) ;
  assign n8718 = ( n8396 & n8716 ) | ( n8396 & ~n8717 ) | ( n8716 & ~n8717 ) ;
  assign n8719 = ( x67 & n8713 ) | ( x67 & ~n8718 ) | ( n8713 & ~n8718 ) ;
  assign n8720 = ( x67 & n8397 ) | ( x67 & ~n8697 ) | ( n8397 & ~n8697 ) ;
  assign n8721 = x67 & n8397 ;
  assign n8722 = ( ~n8402 & n8720 ) | ( ~n8402 & n8721 ) | ( n8720 & n8721 ) ;
  assign n8723 = ( n8402 & n8720 ) | ( n8402 & n8721 ) | ( n8720 & n8721 ) ;
  assign n8724 = ( n8402 & n8722 ) | ( n8402 & ~n8723 ) | ( n8722 & ~n8723 ) ;
  assign n8725 = ( x68 & n8719 ) | ( x68 & ~n8724 ) | ( n8719 & ~n8724 ) ;
  assign n8726 = ( x68 & n8403 ) | ( x68 & ~n8697 ) | ( n8403 & ~n8697 ) ;
  assign n8727 = x68 & n8403 ;
  assign n8728 = ( ~n8408 & n8726 ) | ( ~n8408 & n8727 ) | ( n8726 & n8727 ) ;
  assign n8729 = ( n8408 & n8726 ) | ( n8408 & n8727 ) | ( n8726 & n8727 ) ;
  assign n8730 = ( n8408 & n8728 ) | ( n8408 & ~n8729 ) | ( n8728 & ~n8729 ) ;
  assign n8731 = ( x69 & n8725 ) | ( x69 & ~n8730 ) | ( n8725 & ~n8730 ) ;
  assign n8732 = ( x69 & n8409 ) | ( x69 & ~n8697 ) | ( n8409 & ~n8697 ) ;
  assign n8733 = x69 & n8409 ;
  assign n8734 = ( ~n8414 & n8732 ) | ( ~n8414 & n8733 ) | ( n8732 & n8733 ) ;
  assign n8735 = ( n8414 & n8732 ) | ( n8414 & n8733 ) | ( n8732 & n8733 ) ;
  assign n8736 = ( n8414 & n8734 ) | ( n8414 & ~n8735 ) | ( n8734 & ~n8735 ) ;
  assign n8737 = ( x70 & n8731 ) | ( x70 & ~n8736 ) | ( n8731 & ~n8736 ) ;
  assign n8738 = ( x70 & n8415 ) | ( x70 & ~n8697 ) | ( n8415 & ~n8697 ) ;
  assign n8739 = x70 & n8415 ;
  assign n8740 = ( ~n8420 & n8738 ) | ( ~n8420 & n8739 ) | ( n8738 & n8739 ) ;
  assign n8741 = ( n8420 & n8738 ) | ( n8420 & n8739 ) | ( n8738 & n8739 ) ;
  assign n8742 = ( n8420 & n8740 ) | ( n8420 & ~n8741 ) | ( n8740 & ~n8741 ) ;
  assign n8743 = ( x71 & n8737 ) | ( x71 & ~n8742 ) | ( n8737 & ~n8742 ) ;
  assign n8744 = ( x71 & n8421 ) | ( x71 & ~n8697 ) | ( n8421 & ~n8697 ) ;
  assign n8745 = x71 & n8421 ;
  assign n8746 = ( ~n8426 & n8744 ) | ( ~n8426 & n8745 ) | ( n8744 & n8745 ) ;
  assign n8747 = ( n8426 & n8744 ) | ( n8426 & n8745 ) | ( n8744 & n8745 ) ;
  assign n8748 = ( n8426 & n8746 ) | ( n8426 & ~n8747 ) | ( n8746 & ~n8747 ) ;
  assign n8749 = ( x72 & n8743 ) | ( x72 & ~n8748 ) | ( n8743 & ~n8748 ) ;
  assign n8750 = ( x72 & n8427 ) | ( x72 & ~n8697 ) | ( n8427 & ~n8697 ) ;
  assign n8751 = x72 & n8427 ;
  assign n8752 = ( ~n8432 & n8750 ) | ( ~n8432 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8753 = ( n8432 & n8750 ) | ( n8432 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8754 = ( n8432 & n8752 ) | ( n8432 & ~n8753 ) | ( n8752 & ~n8753 ) ;
  assign n8755 = ( x73 & n8749 ) | ( x73 & ~n8754 ) | ( n8749 & ~n8754 ) ;
  assign n8756 = ( x73 & n8433 ) | ( x73 & ~n8697 ) | ( n8433 & ~n8697 ) ;
  assign n8757 = x73 & n8433 ;
  assign n8758 = ( ~n8438 & n8756 ) | ( ~n8438 & n8757 ) | ( n8756 & n8757 ) ;
  assign n8759 = ( n8438 & n8756 ) | ( n8438 & n8757 ) | ( n8756 & n8757 ) ;
  assign n8760 = ( n8438 & n8758 ) | ( n8438 & ~n8759 ) | ( n8758 & ~n8759 ) ;
  assign n8761 = ( x74 & n8755 ) | ( x74 & ~n8760 ) | ( n8755 & ~n8760 ) ;
  assign n8762 = ( x74 & n8439 ) | ( x74 & ~n8697 ) | ( n8439 & ~n8697 ) ;
  assign n8763 = x74 & n8439 ;
  assign n8764 = ( ~n8444 & n8762 ) | ( ~n8444 & n8763 ) | ( n8762 & n8763 ) ;
  assign n8765 = ( n8444 & n8762 ) | ( n8444 & n8763 ) | ( n8762 & n8763 ) ;
  assign n8766 = ( n8444 & n8764 ) | ( n8444 & ~n8765 ) | ( n8764 & ~n8765 ) ;
  assign n8767 = ( x75 & n8761 ) | ( x75 & ~n8766 ) | ( n8761 & ~n8766 ) ;
  assign n8768 = ( x75 & n8445 ) | ( x75 & ~n8697 ) | ( n8445 & ~n8697 ) ;
  assign n8769 = x75 & n8445 ;
  assign n8770 = ( ~n8450 & n8768 ) | ( ~n8450 & n8769 ) | ( n8768 & n8769 ) ;
  assign n8771 = ( n8450 & n8768 ) | ( n8450 & n8769 ) | ( n8768 & n8769 ) ;
  assign n8772 = ( n8450 & n8770 ) | ( n8450 & ~n8771 ) | ( n8770 & ~n8771 ) ;
  assign n8773 = ( x76 & n8767 ) | ( x76 & ~n8772 ) | ( n8767 & ~n8772 ) ;
  assign n8774 = ( x76 & n8451 ) | ( x76 & ~n8697 ) | ( n8451 & ~n8697 ) ;
  assign n8775 = x76 & n8451 ;
  assign n8776 = ( ~n8456 & n8774 ) | ( ~n8456 & n8775 ) | ( n8774 & n8775 ) ;
  assign n8777 = ( n8456 & n8774 ) | ( n8456 & n8775 ) | ( n8774 & n8775 ) ;
  assign n8778 = ( n8456 & n8776 ) | ( n8456 & ~n8777 ) | ( n8776 & ~n8777 ) ;
  assign n8779 = ( x77 & n8773 ) | ( x77 & ~n8778 ) | ( n8773 & ~n8778 ) ;
  assign n8780 = ( x77 & n8457 ) | ( x77 & ~n8697 ) | ( n8457 & ~n8697 ) ;
  assign n8781 = x77 & n8457 ;
  assign n8782 = ( ~n8462 & n8780 ) | ( ~n8462 & n8781 ) | ( n8780 & n8781 ) ;
  assign n8783 = ( n8462 & n8780 ) | ( n8462 & n8781 ) | ( n8780 & n8781 ) ;
  assign n8784 = ( n8462 & n8782 ) | ( n8462 & ~n8783 ) | ( n8782 & ~n8783 ) ;
  assign n8785 = ( x78 & n8779 ) | ( x78 & ~n8784 ) | ( n8779 & ~n8784 ) ;
  assign n8786 = ( x78 & n8463 ) | ( x78 & ~n8697 ) | ( n8463 & ~n8697 ) ;
  assign n8787 = x78 & n8463 ;
  assign n8788 = ( ~n8468 & n8786 ) | ( ~n8468 & n8787 ) | ( n8786 & n8787 ) ;
  assign n8789 = ( n8468 & n8786 ) | ( n8468 & n8787 ) | ( n8786 & n8787 ) ;
  assign n8790 = ( n8468 & n8788 ) | ( n8468 & ~n8789 ) | ( n8788 & ~n8789 ) ;
  assign n8791 = ( x79 & n8785 ) | ( x79 & ~n8790 ) | ( n8785 & ~n8790 ) ;
  assign n8792 = ( x79 & n8469 ) | ( x79 & ~n8697 ) | ( n8469 & ~n8697 ) ;
  assign n8793 = x79 & n8469 ;
  assign n8794 = ( ~n8474 & n8792 ) | ( ~n8474 & n8793 ) | ( n8792 & n8793 ) ;
  assign n8795 = ( n8474 & n8792 ) | ( n8474 & n8793 ) | ( n8792 & n8793 ) ;
  assign n8796 = ( n8474 & n8794 ) | ( n8474 & ~n8795 ) | ( n8794 & ~n8795 ) ;
  assign n8797 = ( x80 & n8791 ) | ( x80 & ~n8796 ) | ( n8791 & ~n8796 ) ;
  assign n8798 = ( x80 & n8475 ) | ( x80 & ~n8697 ) | ( n8475 & ~n8697 ) ;
  assign n8799 = x80 & n8475 ;
  assign n8800 = ( ~n8480 & n8798 ) | ( ~n8480 & n8799 ) | ( n8798 & n8799 ) ;
  assign n8801 = ( n8480 & n8798 ) | ( n8480 & n8799 ) | ( n8798 & n8799 ) ;
  assign n8802 = ( n8480 & n8800 ) | ( n8480 & ~n8801 ) | ( n8800 & ~n8801 ) ;
  assign n8803 = ( x81 & n8797 ) | ( x81 & ~n8802 ) | ( n8797 & ~n8802 ) ;
  assign n8804 = ( x81 & n8481 ) | ( x81 & ~n8697 ) | ( n8481 & ~n8697 ) ;
  assign n8805 = x81 & n8481 ;
  assign n8806 = ( ~n8486 & n8804 ) | ( ~n8486 & n8805 ) | ( n8804 & n8805 ) ;
  assign n8807 = ( n8486 & n8804 ) | ( n8486 & n8805 ) | ( n8804 & n8805 ) ;
  assign n8808 = ( n8486 & n8806 ) | ( n8486 & ~n8807 ) | ( n8806 & ~n8807 ) ;
  assign n8809 = ( x82 & n8803 ) | ( x82 & ~n8808 ) | ( n8803 & ~n8808 ) ;
  assign n8810 = ( x82 & n8487 ) | ( x82 & ~n8697 ) | ( n8487 & ~n8697 ) ;
  assign n8811 = x82 & n8487 ;
  assign n8812 = ( ~n8492 & n8810 ) | ( ~n8492 & n8811 ) | ( n8810 & n8811 ) ;
  assign n8813 = ( n8492 & n8810 ) | ( n8492 & n8811 ) | ( n8810 & n8811 ) ;
  assign n8814 = ( n8492 & n8812 ) | ( n8492 & ~n8813 ) | ( n8812 & ~n8813 ) ;
  assign n8815 = ( x83 & n8809 ) | ( x83 & ~n8814 ) | ( n8809 & ~n8814 ) ;
  assign n8816 = ( x83 & n8493 ) | ( x83 & ~n8697 ) | ( n8493 & ~n8697 ) ;
  assign n8817 = x83 & n8493 ;
  assign n8818 = ( ~n8498 & n8816 ) | ( ~n8498 & n8817 ) | ( n8816 & n8817 ) ;
  assign n8819 = ( n8498 & n8816 ) | ( n8498 & n8817 ) | ( n8816 & n8817 ) ;
  assign n8820 = ( n8498 & n8818 ) | ( n8498 & ~n8819 ) | ( n8818 & ~n8819 ) ;
  assign n8821 = ( x84 & n8815 ) | ( x84 & ~n8820 ) | ( n8815 & ~n8820 ) ;
  assign n8822 = ( x84 & n8499 ) | ( x84 & ~n8697 ) | ( n8499 & ~n8697 ) ;
  assign n8823 = x84 & n8499 ;
  assign n8824 = ( ~n8504 & n8822 ) | ( ~n8504 & n8823 ) | ( n8822 & n8823 ) ;
  assign n8825 = ( n8504 & n8822 ) | ( n8504 & n8823 ) | ( n8822 & n8823 ) ;
  assign n8826 = ( n8504 & n8824 ) | ( n8504 & ~n8825 ) | ( n8824 & ~n8825 ) ;
  assign n8827 = ( x85 & n8821 ) | ( x85 & ~n8826 ) | ( n8821 & ~n8826 ) ;
  assign n8828 = ( x85 & n8505 ) | ( x85 & ~n8697 ) | ( n8505 & ~n8697 ) ;
  assign n8829 = x85 & n8505 ;
  assign n8830 = ( ~n8510 & n8828 ) | ( ~n8510 & n8829 ) | ( n8828 & n8829 ) ;
  assign n8831 = ( n8510 & n8828 ) | ( n8510 & n8829 ) | ( n8828 & n8829 ) ;
  assign n8832 = ( n8510 & n8830 ) | ( n8510 & ~n8831 ) | ( n8830 & ~n8831 ) ;
  assign n8833 = ( x86 & n8827 ) | ( x86 & ~n8832 ) | ( n8827 & ~n8832 ) ;
  assign n8834 = ( x86 & n8511 ) | ( x86 & ~n8697 ) | ( n8511 & ~n8697 ) ;
  assign n8835 = x86 & n8511 ;
  assign n8836 = ( ~n8516 & n8834 ) | ( ~n8516 & n8835 ) | ( n8834 & n8835 ) ;
  assign n8837 = ( n8516 & n8834 ) | ( n8516 & n8835 ) | ( n8834 & n8835 ) ;
  assign n8838 = ( n8516 & n8836 ) | ( n8516 & ~n8837 ) | ( n8836 & ~n8837 ) ;
  assign n8839 = ( x87 & n8833 ) | ( x87 & ~n8838 ) | ( n8833 & ~n8838 ) ;
  assign n8840 = ( x87 & n8517 ) | ( x87 & ~n8697 ) | ( n8517 & ~n8697 ) ;
  assign n8841 = x87 & n8517 ;
  assign n8842 = ( ~n8522 & n8840 ) | ( ~n8522 & n8841 ) | ( n8840 & n8841 ) ;
  assign n8843 = ( n8522 & n8840 ) | ( n8522 & n8841 ) | ( n8840 & n8841 ) ;
  assign n8844 = ( n8522 & n8842 ) | ( n8522 & ~n8843 ) | ( n8842 & ~n8843 ) ;
  assign n8845 = ( x88 & n8839 ) | ( x88 & ~n8844 ) | ( n8839 & ~n8844 ) ;
  assign n8846 = ( x88 & n8523 ) | ( x88 & ~n8697 ) | ( n8523 & ~n8697 ) ;
  assign n8847 = x88 & n8523 ;
  assign n8848 = ( ~n8528 & n8846 ) | ( ~n8528 & n8847 ) | ( n8846 & n8847 ) ;
  assign n8849 = ( n8528 & n8846 ) | ( n8528 & n8847 ) | ( n8846 & n8847 ) ;
  assign n8850 = ( n8528 & n8848 ) | ( n8528 & ~n8849 ) | ( n8848 & ~n8849 ) ;
  assign n8851 = ( x89 & n8845 ) | ( x89 & ~n8850 ) | ( n8845 & ~n8850 ) ;
  assign n8852 = ( x89 & n8529 ) | ( x89 & ~n8697 ) | ( n8529 & ~n8697 ) ;
  assign n8853 = x89 & n8529 ;
  assign n8854 = ( ~n8534 & n8852 ) | ( ~n8534 & n8853 ) | ( n8852 & n8853 ) ;
  assign n8855 = ( n8534 & n8852 ) | ( n8534 & n8853 ) | ( n8852 & n8853 ) ;
  assign n8856 = ( n8534 & n8854 ) | ( n8534 & ~n8855 ) | ( n8854 & ~n8855 ) ;
  assign n8857 = ( x90 & n8851 ) | ( x90 & ~n8856 ) | ( n8851 & ~n8856 ) ;
  assign n8858 = ( x90 & n8535 ) | ( x90 & ~n8697 ) | ( n8535 & ~n8697 ) ;
  assign n8859 = x90 & n8535 ;
  assign n8860 = ( ~n8540 & n8858 ) | ( ~n8540 & n8859 ) | ( n8858 & n8859 ) ;
  assign n8861 = ( n8540 & n8858 ) | ( n8540 & n8859 ) | ( n8858 & n8859 ) ;
  assign n8862 = ( n8540 & n8860 ) | ( n8540 & ~n8861 ) | ( n8860 & ~n8861 ) ;
  assign n8863 = ( x91 & n8857 ) | ( x91 & ~n8862 ) | ( n8857 & ~n8862 ) ;
  assign n8864 = ( x91 & n8541 ) | ( x91 & ~n8697 ) | ( n8541 & ~n8697 ) ;
  assign n8865 = x91 & n8541 ;
  assign n8866 = ( ~n8546 & n8864 ) | ( ~n8546 & n8865 ) | ( n8864 & n8865 ) ;
  assign n8867 = ( n8546 & n8864 ) | ( n8546 & n8865 ) | ( n8864 & n8865 ) ;
  assign n8868 = ( n8546 & n8866 ) | ( n8546 & ~n8867 ) | ( n8866 & ~n8867 ) ;
  assign n8869 = ( x92 & n8863 ) | ( x92 & ~n8868 ) | ( n8863 & ~n8868 ) ;
  assign n8870 = ( x92 & n8547 ) | ( x92 & ~n8697 ) | ( n8547 & ~n8697 ) ;
  assign n8871 = x92 & n8547 ;
  assign n8872 = ( ~n8552 & n8870 ) | ( ~n8552 & n8871 ) | ( n8870 & n8871 ) ;
  assign n8873 = ( n8552 & n8870 ) | ( n8552 & n8871 ) | ( n8870 & n8871 ) ;
  assign n8874 = ( n8552 & n8872 ) | ( n8552 & ~n8873 ) | ( n8872 & ~n8873 ) ;
  assign n8875 = ( x93 & n8869 ) | ( x93 & ~n8874 ) | ( n8869 & ~n8874 ) ;
  assign n8876 = ( x93 & n8553 ) | ( x93 & ~n8697 ) | ( n8553 & ~n8697 ) ;
  assign n8877 = x93 & n8553 ;
  assign n8878 = ( ~n8558 & n8876 ) | ( ~n8558 & n8877 ) | ( n8876 & n8877 ) ;
  assign n8879 = ( n8558 & n8876 ) | ( n8558 & n8877 ) | ( n8876 & n8877 ) ;
  assign n8880 = ( n8558 & n8878 ) | ( n8558 & ~n8879 ) | ( n8878 & ~n8879 ) ;
  assign n8881 = ( x94 & n8875 ) | ( x94 & ~n8880 ) | ( n8875 & ~n8880 ) ;
  assign n8882 = ( x94 & n8559 ) | ( x94 & ~n8697 ) | ( n8559 & ~n8697 ) ;
  assign n8883 = x94 & n8559 ;
  assign n8884 = ( ~n8564 & n8882 ) | ( ~n8564 & n8883 ) | ( n8882 & n8883 ) ;
  assign n8885 = ( n8564 & n8882 ) | ( n8564 & n8883 ) | ( n8882 & n8883 ) ;
  assign n8886 = ( n8564 & n8884 ) | ( n8564 & ~n8885 ) | ( n8884 & ~n8885 ) ;
  assign n8887 = ( x95 & n8881 ) | ( x95 & ~n8886 ) | ( n8881 & ~n8886 ) ;
  assign n8888 = ( x95 & n8565 ) | ( x95 & ~n8697 ) | ( n8565 & ~n8697 ) ;
  assign n8889 = x95 & n8565 ;
  assign n8890 = ( ~n8570 & n8888 ) | ( ~n8570 & n8889 ) | ( n8888 & n8889 ) ;
  assign n8891 = ( n8570 & n8888 ) | ( n8570 & n8889 ) | ( n8888 & n8889 ) ;
  assign n8892 = ( n8570 & n8890 ) | ( n8570 & ~n8891 ) | ( n8890 & ~n8891 ) ;
  assign n8893 = ( x96 & n8887 ) | ( x96 & ~n8892 ) | ( n8887 & ~n8892 ) ;
  assign n8894 = ( x96 & n8571 ) | ( x96 & ~n8697 ) | ( n8571 & ~n8697 ) ;
  assign n8895 = x96 & n8571 ;
  assign n8896 = ( ~n8576 & n8894 ) | ( ~n8576 & n8895 ) | ( n8894 & n8895 ) ;
  assign n8897 = ( n8576 & n8894 ) | ( n8576 & n8895 ) | ( n8894 & n8895 ) ;
  assign n8898 = ( n8576 & n8896 ) | ( n8576 & ~n8897 ) | ( n8896 & ~n8897 ) ;
  assign n8899 = ( x97 & n8893 ) | ( x97 & ~n8898 ) | ( n8893 & ~n8898 ) ;
  assign n8900 = ( x97 & n8577 ) | ( x97 & ~n8697 ) | ( n8577 & ~n8697 ) ;
  assign n8901 = x97 & n8577 ;
  assign n8902 = ( ~n8582 & n8900 ) | ( ~n8582 & n8901 ) | ( n8900 & n8901 ) ;
  assign n8903 = ( n8582 & n8900 ) | ( n8582 & n8901 ) | ( n8900 & n8901 ) ;
  assign n8904 = ( n8582 & n8902 ) | ( n8582 & ~n8903 ) | ( n8902 & ~n8903 ) ;
  assign n8905 = ( x98 & n8899 ) | ( x98 & ~n8904 ) | ( n8899 & ~n8904 ) ;
  assign n8906 = ( x98 & n8583 ) | ( x98 & ~n8697 ) | ( n8583 & ~n8697 ) ;
  assign n8907 = x98 & n8583 ;
  assign n8908 = ( ~n8588 & n8906 ) | ( ~n8588 & n8907 ) | ( n8906 & n8907 ) ;
  assign n8909 = ( n8588 & n8906 ) | ( n8588 & n8907 ) | ( n8906 & n8907 ) ;
  assign n8910 = ( n8588 & n8908 ) | ( n8588 & ~n8909 ) | ( n8908 & ~n8909 ) ;
  assign n8911 = ( x99 & n8905 ) | ( x99 & ~n8910 ) | ( n8905 & ~n8910 ) ;
  assign n8912 = ( x99 & n8589 ) | ( x99 & ~n8697 ) | ( n8589 & ~n8697 ) ;
  assign n8913 = x99 & n8589 ;
  assign n8914 = ( ~n8594 & n8912 ) | ( ~n8594 & n8913 ) | ( n8912 & n8913 ) ;
  assign n8915 = ( n8594 & n8912 ) | ( n8594 & n8913 ) | ( n8912 & n8913 ) ;
  assign n8916 = ( n8594 & n8914 ) | ( n8594 & ~n8915 ) | ( n8914 & ~n8915 ) ;
  assign n8917 = ( x100 & n8911 ) | ( x100 & ~n8916 ) | ( n8911 & ~n8916 ) ;
  assign n8918 = ( x100 & n8595 ) | ( x100 & ~n8697 ) | ( n8595 & ~n8697 ) ;
  assign n8919 = x100 & n8595 ;
  assign n8920 = ( ~n8600 & n8918 ) | ( ~n8600 & n8919 ) | ( n8918 & n8919 ) ;
  assign n8921 = ( n8600 & n8918 ) | ( n8600 & n8919 ) | ( n8918 & n8919 ) ;
  assign n8922 = ( n8600 & n8920 ) | ( n8600 & ~n8921 ) | ( n8920 & ~n8921 ) ;
  assign n8923 = ( x101 & n8917 ) | ( x101 & ~n8922 ) | ( n8917 & ~n8922 ) ;
  assign n8924 = ( x101 & n8601 ) | ( x101 & ~n8697 ) | ( n8601 & ~n8697 ) ;
  assign n8925 = x101 & n8601 ;
  assign n8926 = ( ~n8606 & n8924 ) | ( ~n8606 & n8925 ) | ( n8924 & n8925 ) ;
  assign n8927 = ( n8606 & n8924 ) | ( n8606 & n8925 ) | ( n8924 & n8925 ) ;
  assign n8928 = ( n8606 & n8926 ) | ( n8606 & ~n8927 ) | ( n8926 & ~n8927 ) ;
  assign n8929 = ( x102 & n8923 ) | ( x102 & ~n8928 ) | ( n8923 & ~n8928 ) ;
  assign n8930 = ( x102 & n8607 ) | ( x102 & ~n8697 ) | ( n8607 & ~n8697 ) ;
  assign n8931 = x102 & n8607 ;
  assign n8932 = ( ~n8612 & n8930 ) | ( ~n8612 & n8931 ) | ( n8930 & n8931 ) ;
  assign n8933 = ( n8612 & n8930 ) | ( n8612 & n8931 ) | ( n8930 & n8931 ) ;
  assign n8934 = ( n8612 & n8932 ) | ( n8612 & ~n8933 ) | ( n8932 & ~n8933 ) ;
  assign n8935 = ( x103 & n8929 ) | ( x103 & ~n8934 ) | ( n8929 & ~n8934 ) ;
  assign n8936 = ( x103 & n8613 ) | ( x103 & ~n8697 ) | ( n8613 & ~n8697 ) ;
  assign n8937 = x103 & n8613 ;
  assign n8938 = ( ~n8618 & n8936 ) | ( ~n8618 & n8937 ) | ( n8936 & n8937 ) ;
  assign n8939 = ( n8618 & n8936 ) | ( n8618 & n8937 ) | ( n8936 & n8937 ) ;
  assign n8940 = ( n8618 & n8938 ) | ( n8618 & ~n8939 ) | ( n8938 & ~n8939 ) ;
  assign n8941 = ( x104 & n8935 ) | ( x104 & ~n8940 ) | ( n8935 & ~n8940 ) ;
  assign n8942 = ( x104 & n8619 ) | ( x104 & ~n8697 ) | ( n8619 & ~n8697 ) ;
  assign n8943 = x104 & n8619 ;
  assign n8944 = ( ~n8624 & n8942 ) | ( ~n8624 & n8943 ) | ( n8942 & n8943 ) ;
  assign n8945 = ( n8624 & n8942 ) | ( n8624 & n8943 ) | ( n8942 & n8943 ) ;
  assign n8946 = ( n8624 & n8944 ) | ( n8624 & ~n8945 ) | ( n8944 & ~n8945 ) ;
  assign n8947 = ( x105 & n8941 ) | ( x105 & ~n8946 ) | ( n8941 & ~n8946 ) ;
  assign n8948 = ( x105 & n8625 ) | ( x105 & ~n8697 ) | ( n8625 & ~n8697 ) ;
  assign n8949 = x105 & n8625 ;
  assign n8950 = ( ~n8630 & n8948 ) | ( ~n8630 & n8949 ) | ( n8948 & n8949 ) ;
  assign n8951 = ( n8630 & n8948 ) | ( n8630 & n8949 ) | ( n8948 & n8949 ) ;
  assign n8952 = ( n8630 & n8950 ) | ( n8630 & ~n8951 ) | ( n8950 & ~n8951 ) ;
  assign n8953 = ( x106 & n8947 ) | ( x106 & ~n8952 ) | ( n8947 & ~n8952 ) ;
  assign n8954 = ( x106 & n8631 ) | ( x106 & ~n8697 ) | ( n8631 & ~n8697 ) ;
  assign n8955 = x106 & n8631 ;
  assign n8956 = ( ~n8636 & n8954 ) | ( ~n8636 & n8955 ) | ( n8954 & n8955 ) ;
  assign n8957 = ( n8636 & n8954 ) | ( n8636 & n8955 ) | ( n8954 & n8955 ) ;
  assign n8958 = ( n8636 & n8956 ) | ( n8636 & ~n8957 ) | ( n8956 & ~n8957 ) ;
  assign n8959 = ( x107 & n8953 ) | ( x107 & ~n8958 ) | ( n8953 & ~n8958 ) ;
  assign n8960 = ( x107 & n8637 ) | ( x107 & ~n8697 ) | ( n8637 & ~n8697 ) ;
  assign n8961 = x107 & n8637 ;
  assign n8962 = ( ~n8642 & n8960 ) | ( ~n8642 & n8961 ) | ( n8960 & n8961 ) ;
  assign n8963 = ( n8642 & n8960 ) | ( n8642 & n8961 ) | ( n8960 & n8961 ) ;
  assign n8964 = ( n8642 & n8962 ) | ( n8642 & ~n8963 ) | ( n8962 & ~n8963 ) ;
  assign n8965 = ( x108 & n8959 ) | ( x108 & ~n8964 ) | ( n8959 & ~n8964 ) ;
  assign n8966 = ( x108 & n8643 ) | ( x108 & ~n8697 ) | ( n8643 & ~n8697 ) ;
  assign n8967 = x108 & n8643 ;
  assign n8968 = ( ~n8648 & n8966 ) | ( ~n8648 & n8967 ) | ( n8966 & n8967 ) ;
  assign n8969 = ( n8648 & n8966 ) | ( n8648 & n8967 ) | ( n8966 & n8967 ) ;
  assign n8970 = ( n8648 & n8968 ) | ( n8648 & ~n8969 ) | ( n8968 & ~n8969 ) ;
  assign n8971 = ( x109 & n8965 ) | ( x109 & ~n8970 ) | ( n8965 & ~n8970 ) ;
  assign n8972 = ( x109 & n8649 ) | ( x109 & ~n8697 ) | ( n8649 & ~n8697 ) ;
  assign n8973 = x109 & n8649 ;
  assign n8974 = ( ~n8654 & n8972 ) | ( ~n8654 & n8973 ) | ( n8972 & n8973 ) ;
  assign n8975 = ( n8654 & n8972 ) | ( n8654 & n8973 ) | ( n8972 & n8973 ) ;
  assign n8976 = ( n8654 & n8974 ) | ( n8654 & ~n8975 ) | ( n8974 & ~n8975 ) ;
  assign n8977 = ( x110 & n8971 ) | ( x110 & ~n8976 ) | ( n8971 & ~n8976 ) ;
  assign n8978 = ( x110 & n8655 ) | ( x110 & ~n8697 ) | ( n8655 & ~n8697 ) ;
  assign n8979 = x110 & n8655 ;
  assign n8980 = ( ~n8660 & n8978 ) | ( ~n8660 & n8979 ) | ( n8978 & n8979 ) ;
  assign n8981 = ( n8660 & n8978 ) | ( n8660 & n8979 ) | ( n8978 & n8979 ) ;
  assign n8982 = ( n8660 & n8980 ) | ( n8660 & ~n8981 ) | ( n8980 & ~n8981 ) ;
  assign n8983 = ( x111 & n8977 ) | ( x111 & ~n8982 ) | ( n8977 & ~n8982 ) ;
  assign n8984 = ( x111 & n8661 ) | ( x111 & ~n8697 ) | ( n8661 & ~n8697 ) ;
  assign n8985 = x111 & n8661 ;
  assign n8986 = ( ~n8666 & n8984 ) | ( ~n8666 & n8985 ) | ( n8984 & n8985 ) ;
  assign n8987 = ( n8666 & n8984 ) | ( n8666 & n8985 ) | ( n8984 & n8985 ) ;
  assign n8988 = ( n8666 & n8986 ) | ( n8666 & ~n8987 ) | ( n8986 & ~n8987 ) ;
  assign n8989 = ( x112 & n8983 ) | ( x112 & ~n8988 ) | ( n8983 & ~n8988 ) ;
  assign n8990 = ( x112 & n8667 ) | ( x112 & ~n8697 ) | ( n8667 & ~n8697 ) ;
  assign n8991 = x112 & n8667 ;
  assign n8992 = ( ~n8672 & n8990 ) | ( ~n8672 & n8991 ) | ( n8990 & n8991 ) ;
  assign n8993 = ( n8672 & n8990 ) | ( n8672 & n8991 ) | ( n8990 & n8991 ) ;
  assign n8994 = ( n8672 & n8992 ) | ( n8672 & ~n8993 ) | ( n8992 & ~n8993 ) ;
  assign n8995 = ( x113 & n8989 ) | ( x113 & ~n8994 ) | ( n8989 & ~n8994 ) ;
  assign n8996 = ( x113 & n8673 ) | ( x113 & ~n8697 ) | ( n8673 & ~n8697 ) ;
  assign n8997 = x113 & n8673 ;
  assign n8998 = ( ~n8678 & n8996 ) | ( ~n8678 & n8997 ) | ( n8996 & n8997 ) ;
  assign n8999 = ( n8678 & n8996 ) | ( n8678 & n8997 ) | ( n8996 & n8997 ) ;
  assign n9000 = ( n8678 & n8998 ) | ( n8678 & ~n8999 ) | ( n8998 & ~n8999 ) ;
  assign n9001 = ( x114 & n8995 ) | ( x114 & ~n9000 ) | ( n8995 & ~n9000 ) ;
  assign n9002 = ( x114 & n8679 ) | ( x114 & ~n8697 ) | ( n8679 & ~n8697 ) ;
  assign n9003 = x114 & n8679 ;
  assign n9004 = ( ~n8684 & n9002 ) | ( ~n8684 & n9003 ) | ( n9002 & n9003 ) ;
  assign n9005 = ( n8684 & n9002 ) | ( n8684 & n9003 ) | ( n9002 & n9003 ) ;
  assign n9006 = ( n8684 & n9004 ) | ( n8684 & ~n9005 ) | ( n9004 & ~n9005 ) ;
  assign n9007 = ( x115 & n9001 ) | ( x115 & ~n9006 ) | ( n9001 & ~n9006 ) ;
  assign n9008 = ( x115 & n8685 ) | ( x115 & ~n8697 ) | ( n8685 & ~n8697 ) ;
  assign n9009 = x115 & n8685 ;
  assign n9010 = ( ~n8690 & n9008 ) | ( ~n8690 & n9009 ) | ( n9008 & n9009 ) ;
  assign n9011 = ( n8690 & n9008 ) | ( n8690 & n9009 ) | ( n9008 & n9009 ) ;
  assign n9012 = ( n8690 & n9010 ) | ( n8690 & ~n9011 ) | ( n9010 & ~n9011 ) ;
  assign n9013 = ( x116 & n9007 ) | ( x116 & ~n9012 ) | ( n9007 & ~n9012 ) ;
  assign n9014 = ( x117 & n139 ) | ( x117 & n8692 ) | ( n139 & n8692 ) ;
  assign n9015 = x117 | n8692 ;
  assign n9016 = ( n8695 & n9014 ) | ( n8695 & ~n9015 ) | ( n9014 & ~n9015 ) ;
  assign n9017 = ( x117 & ~n8702 ) | ( x117 & n9013 ) | ( ~n8702 & n9013 ) ;
  assign n9018 = ( x118 & ~n9016 ) | ( x118 & n9017 ) | ( ~n9016 & n9017 ) ;
  assign n9019 = n138 | n9018 ;
  assign n9020 = ( x117 & n9013 ) | ( x117 & n9019 ) | ( n9013 & n9019 ) ;
  assign n9021 = x117 | n9013 ;
  assign n9022 = ( ~n8702 & n9020 ) | ( ~n8702 & n9021 ) | ( n9020 & n9021 ) ;
  assign n9023 = ( n8702 & n9020 ) | ( n8702 & n9021 ) | ( n9020 & n9021 ) ;
  assign n9024 = ( n8702 & n9022 ) | ( n8702 & ~n9023 ) | ( n9022 & ~n9023 ) ;
  assign n9025 = ~x8 & x64 ;
  assign n9026 = ~x9 & n9019 ;
  assign n9027 = ( x9 & ~x64 ) | ( x9 & n9019 ) | ( ~x64 & n9019 ) ;
  assign n9028 = ( n8703 & ~n9026 ) | ( n8703 & n9027 ) | ( ~n9026 & n9027 ) ;
  assign n9029 = ( x65 & n9025 ) | ( x65 & ~n9028 ) | ( n9025 & ~n9028 ) ;
  assign n9030 = ( x65 & n8703 ) | ( x65 & n9019 ) | ( n8703 & n9019 ) ;
  assign n9031 = x65 | n8703 ;
  assign n9032 = ( ~n8706 & n9030 ) | ( ~n8706 & n9031 ) | ( n9030 & n9031 ) ;
  assign n9033 = ( n8706 & n9030 ) | ( n8706 & n9031 ) | ( n9030 & n9031 ) ;
  assign n9034 = ( n8706 & n9032 ) | ( n8706 & ~n9033 ) | ( n9032 & ~n9033 ) ;
  assign n9035 = ( x66 & n9029 ) | ( x66 & ~n9034 ) | ( n9029 & ~n9034 ) ;
  assign n9036 = ( x66 & n8707 ) | ( x66 & n9019 ) | ( n8707 & n9019 ) ;
  assign n9037 = x66 | n8707 ;
  assign n9038 = ( ~n8712 & n9036 ) | ( ~n8712 & n9037 ) | ( n9036 & n9037 ) ;
  assign n9039 = ( n8712 & n9036 ) | ( n8712 & n9037 ) | ( n9036 & n9037 ) ;
  assign n9040 = ( n8712 & n9038 ) | ( n8712 & ~n9039 ) | ( n9038 & ~n9039 ) ;
  assign n9041 = ( x67 & n9035 ) | ( x67 & ~n9040 ) | ( n9035 & ~n9040 ) ;
  assign n9042 = ( x67 & n8713 ) | ( x67 & ~n9019 ) | ( n8713 & ~n9019 ) ;
  assign n9043 = x67 & n8713 ;
  assign n9044 = ( ~n8718 & n9042 ) | ( ~n8718 & n9043 ) | ( n9042 & n9043 ) ;
  assign n9045 = ( n8718 & n9042 ) | ( n8718 & n9043 ) | ( n9042 & n9043 ) ;
  assign n9046 = ( n8718 & n9044 ) | ( n8718 & ~n9045 ) | ( n9044 & ~n9045 ) ;
  assign n9047 = ( x68 & n9041 ) | ( x68 & ~n9046 ) | ( n9041 & ~n9046 ) ;
  assign n9048 = ( x68 & n8719 ) | ( x68 & ~n9019 ) | ( n8719 & ~n9019 ) ;
  assign n9049 = x68 & n8719 ;
  assign n9050 = ( ~n8724 & n9048 ) | ( ~n8724 & n9049 ) | ( n9048 & n9049 ) ;
  assign n9051 = ( n8724 & n9048 ) | ( n8724 & n9049 ) | ( n9048 & n9049 ) ;
  assign n9052 = ( n8724 & n9050 ) | ( n8724 & ~n9051 ) | ( n9050 & ~n9051 ) ;
  assign n9053 = ( x69 & n9047 ) | ( x69 & ~n9052 ) | ( n9047 & ~n9052 ) ;
  assign n9054 = ( x69 & n8725 ) | ( x69 & ~n9019 ) | ( n8725 & ~n9019 ) ;
  assign n9055 = x69 & n8725 ;
  assign n9056 = ( ~n8730 & n9054 ) | ( ~n8730 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9057 = ( n8730 & n9054 ) | ( n8730 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9058 = ( n8730 & n9056 ) | ( n8730 & ~n9057 ) | ( n9056 & ~n9057 ) ;
  assign n9059 = ( x70 & n9053 ) | ( x70 & ~n9058 ) | ( n9053 & ~n9058 ) ;
  assign n9060 = ( x70 & n8731 ) | ( x70 & ~n9019 ) | ( n8731 & ~n9019 ) ;
  assign n9061 = x70 & n8731 ;
  assign n9062 = ( ~n8736 & n9060 ) | ( ~n8736 & n9061 ) | ( n9060 & n9061 ) ;
  assign n9063 = ( n8736 & n9060 ) | ( n8736 & n9061 ) | ( n9060 & n9061 ) ;
  assign n9064 = ( n8736 & n9062 ) | ( n8736 & ~n9063 ) | ( n9062 & ~n9063 ) ;
  assign n9065 = ( x71 & n9059 ) | ( x71 & ~n9064 ) | ( n9059 & ~n9064 ) ;
  assign n9066 = ( x71 & n8737 ) | ( x71 & ~n9019 ) | ( n8737 & ~n9019 ) ;
  assign n9067 = x71 & n8737 ;
  assign n9068 = ( ~n8742 & n9066 ) | ( ~n8742 & n9067 ) | ( n9066 & n9067 ) ;
  assign n9069 = ( n8742 & n9066 ) | ( n8742 & n9067 ) | ( n9066 & n9067 ) ;
  assign n9070 = ( n8742 & n9068 ) | ( n8742 & ~n9069 ) | ( n9068 & ~n9069 ) ;
  assign n9071 = ( x72 & n9065 ) | ( x72 & ~n9070 ) | ( n9065 & ~n9070 ) ;
  assign n9072 = ( x72 & n8743 ) | ( x72 & ~n9019 ) | ( n8743 & ~n9019 ) ;
  assign n9073 = x72 & n8743 ;
  assign n9074 = ( ~n8748 & n9072 ) | ( ~n8748 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9075 = ( n8748 & n9072 ) | ( n8748 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9076 = ( n8748 & n9074 ) | ( n8748 & ~n9075 ) | ( n9074 & ~n9075 ) ;
  assign n9077 = ( x73 & n9071 ) | ( x73 & ~n9076 ) | ( n9071 & ~n9076 ) ;
  assign n9078 = ( x73 & n8749 ) | ( x73 & ~n9019 ) | ( n8749 & ~n9019 ) ;
  assign n9079 = x73 & n8749 ;
  assign n9080 = ( ~n8754 & n9078 ) | ( ~n8754 & n9079 ) | ( n9078 & n9079 ) ;
  assign n9081 = ( n8754 & n9078 ) | ( n8754 & n9079 ) | ( n9078 & n9079 ) ;
  assign n9082 = ( n8754 & n9080 ) | ( n8754 & ~n9081 ) | ( n9080 & ~n9081 ) ;
  assign n9083 = ( x74 & n9077 ) | ( x74 & ~n9082 ) | ( n9077 & ~n9082 ) ;
  assign n9084 = ( x74 & n8755 ) | ( x74 & ~n9019 ) | ( n8755 & ~n9019 ) ;
  assign n9085 = x74 & n8755 ;
  assign n9086 = ( ~n8760 & n9084 ) | ( ~n8760 & n9085 ) | ( n9084 & n9085 ) ;
  assign n9087 = ( n8760 & n9084 ) | ( n8760 & n9085 ) | ( n9084 & n9085 ) ;
  assign n9088 = ( n8760 & n9086 ) | ( n8760 & ~n9087 ) | ( n9086 & ~n9087 ) ;
  assign n9089 = ( x75 & n9083 ) | ( x75 & ~n9088 ) | ( n9083 & ~n9088 ) ;
  assign n9090 = ( x75 & n8761 ) | ( x75 & ~n9019 ) | ( n8761 & ~n9019 ) ;
  assign n9091 = x75 & n8761 ;
  assign n9092 = ( ~n8766 & n9090 ) | ( ~n8766 & n9091 ) | ( n9090 & n9091 ) ;
  assign n9093 = ( n8766 & n9090 ) | ( n8766 & n9091 ) | ( n9090 & n9091 ) ;
  assign n9094 = ( n8766 & n9092 ) | ( n8766 & ~n9093 ) | ( n9092 & ~n9093 ) ;
  assign n9095 = ( x76 & n9089 ) | ( x76 & ~n9094 ) | ( n9089 & ~n9094 ) ;
  assign n9096 = ( x76 & n8767 ) | ( x76 & ~n9019 ) | ( n8767 & ~n9019 ) ;
  assign n9097 = x76 & n8767 ;
  assign n9098 = ( ~n8772 & n9096 ) | ( ~n8772 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9099 = ( n8772 & n9096 ) | ( n8772 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9100 = ( n8772 & n9098 ) | ( n8772 & ~n9099 ) | ( n9098 & ~n9099 ) ;
  assign n9101 = ( x77 & n9095 ) | ( x77 & ~n9100 ) | ( n9095 & ~n9100 ) ;
  assign n9102 = ( x77 & n8773 ) | ( x77 & ~n9019 ) | ( n8773 & ~n9019 ) ;
  assign n9103 = x77 & n8773 ;
  assign n9104 = ( ~n8778 & n9102 ) | ( ~n8778 & n9103 ) | ( n9102 & n9103 ) ;
  assign n9105 = ( n8778 & n9102 ) | ( n8778 & n9103 ) | ( n9102 & n9103 ) ;
  assign n9106 = ( n8778 & n9104 ) | ( n8778 & ~n9105 ) | ( n9104 & ~n9105 ) ;
  assign n9107 = ( x78 & n9101 ) | ( x78 & ~n9106 ) | ( n9101 & ~n9106 ) ;
  assign n9108 = ( x78 & n8779 ) | ( x78 & ~n9019 ) | ( n8779 & ~n9019 ) ;
  assign n9109 = x78 & n8779 ;
  assign n9110 = ( ~n8784 & n9108 ) | ( ~n8784 & n9109 ) | ( n9108 & n9109 ) ;
  assign n9111 = ( n8784 & n9108 ) | ( n8784 & n9109 ) | ( n9108 & n9109 ) ;
  assign n9112 = ( n8784 & n9110 ) | ( n8784 & ~n9111 ) | ( n9110 & ~n9111 ) ;
  assign n9113 = ( x79 & n9107 ) | ( x79 & ~n9112 ) | ( n9107 & ~n9112 ) ;
  assign n9114 = ( x79 & n8785 ) | ( x79 & ~n9019 ) | ( n8785 & ~n9019 ) ;
  assign n9115 = x79 & n8785 ;
  assign n9116 = ( ~n8790 & n9114 ) | ( ~n8790 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9117 = ( n8790 & n9114 ) | ( n8790 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9118 = ( n8790 & n9116 ) | ( n8790 & ~n9117 ) | ( n9116 & ~n9117 ) ;
  assign n9119 = ( x80 & n9113 ) | ( x80 & ~n9118 ) | ( n9113 & ~n9118 ) ;
  assign n9120 = ( x80 & n8791 ) | ( x80 & ~n9019 ) | ( n8791 & ~n9019 ) ;
  assign n9121 = x80 & n8791 ;
  assign n9122 = ( ~n8796 & n9120 ) | ( ~n8796 & n9121 ) | ( n9120 & n9121 ) ;
  assign n9123 = ( n8796 & n9120 ) | ( n8796 & n9121 ) | ( n9120 & n9121 ) ;
  assign n9124 = ( n8796 & n9122 ) | ( n8796 & ~n9123 ) | ( n9122 & ~n9123 ) ;
  assign n9125 = ( x81 & n9119 ) | ( x81 & ~n9124 ) | ( n9119 & ~n9124 ) ;
  assign n9126 = ( x81 & n8797 ) | ( x81 & ~n9019 ) | ( n8797 & ~n9019 ) ;
  assign n9127 = x81 & n8797 ;
  assign n9128 = ( ~n8802 & n9126 ) | ( ~n8802 & n9127 ) | ( n9126 & n9127 ) ;
  assign n9129 = ( n8802 & n9126 ) | ( n8802 & n9127 ) | ( n9126 & n9127 ) ;
  assign n9130 = ( n8802 & n9128 ) | ( n8802 & ~n9129 ) | ( n9128 & ~n9129 ) ;
  assign n9131 = ( x82 & n9125 ) | ( x82 & ~n9130 ) | ( n9125 & ~n9130 ) ;
  assign n9132 = ( x82 & n8803 ) | ( x82 & ~n9019 ) | ( n8803 & ~n9019 ) ;
  assign n9133 = x82 & n8803 ;
  assign n9134 = ( ~n8808 & n9132 ) | ( ~n8808 & n9133 ) | ( n9132 & n9133 ) ;
  assign n9135 = ( n8808 & n9132 ) | ( n8808 & n9133 ) | ( n9132 & n9133 ) ;
  assign n9136 = ( n8808 & n9134 ) | ( n8808 & ~n9135 ) | ( n9134 & ~n9135 ) ;
  assign n9137 = ( x83 & n9131 ) | ( x83 & ~n9136 ) | ( n9131 & ~n9136 ) ;
  assign n9138 = ( x83 & n8809 ) | ( x83 & ~n9019 ) | ( n8809 & ~n9019 ) ;
  assign n9139 = x83 & n8809 ;
  assign n9140 = ( ~n8814 & n9138 ) | ( ~n8814 & n9139 ) | ( n9138 & n9139 ) ;
  assign n9141 = ( n8814 & n9138 ) | ( n8814 & n9139 ) | ( n9138 & n9139 ) ;
  assign n9142 = ( n8814 & n9140 ) | ( n8814 & ~n9141 ) | ( n9140 & ~n9141 ) ;
  assign n9143 = ( x84 & n9137 ) | ( x84 & ~n9142 ) | ( n9137 & ~n9142 ) ;
  assign n9144 = ( x84 & n8815 ) | ( x84 & ~n9019 ) | ( n8815 & ~n9019 ) ;
  assign n9145 = x84 & n8815 ;
  assign n9146 = ( ~n8820 & n9144 ) | ( ~n8820 & n9145 ) | ( n9144 & n9145 ) ;
  assign n9147 = ( n8820 & n9144 ) | ( n8820 & n9145 ) | ( n9144 & n9145 ) ;
  assign n9148 = ( n8820 & n9146 ) | ( n8820 & ~n9147 ) | ( n9146 & ~n9147 ) ;
  assign n9149 = ( x85 & n9143 ) | ( x85 & ~n9148 ) | ( n9143 & ~n9148 ) ;
  assign n9150 = ( x85 & n8821 ) | ( x85 & ~n9019 ) | ( n8821 & ~n9019 ) ;
  assign n9151 = x85 & n8821 ;
  assign n9152 = ( ~n8826 & n9150 ) | ( ~n8826 & n9151 ) | ( n9150 & n9151 ) ;
  assign n9153 = ( n8826 & n9150 ) | ( n8826 & n9151 ) | ( n9150 & n9151 ) ;
  assign n9154 = ( n8826 & n9152 ) | ( n8826 & ~n9153 ) | ( n9152 & ~n9153 ) ;
  assign n9155 = ( x86 & n9149 ) | ( x86 & ~n9154 ) | ( n9149 & ~n9154 ) ;
  assign n9156 = ( x86 & n8827 ) | ( x86 & ~n9019 ) | ( n8827 & ~n9019 ) ;
  assign n9157 = x86 & n8827 ;
  assign n9158 = ( ~n8832 & n9156 ) | ( ~n8832 & n9157 ) | ( n9156 & n9157 ) ;
  assign n9159 = ( n8832 & n9156 ) | ( n8832 & n9157 ) | ( n9156 & n9157 ) ;
  assign n9160 = ( n8832 & n9158 ) | ( n8832 & ~n9159 ) | ( n9158 & ~n9159 ) ;
  assign n9161 = ( x87 & n9155 ) | ( x87 & ~n9160 ) | ( n9155 & ~n9160 ) ;
  assign n9162 = ( x87 & n8833 ) | ( x87 & ~n9019 ) | ( n8833 & ~n9019 ) ;
  assign n9163 = x87 & n8833 ;
  assign n9164 = ( ~n8838 & n9162 ) | ( ~n8838 & n9163 ) | ( n9162 & n9163 ) ;
  assign n9165 = ( n8838 & n9162 ) | ( n8838 & n9163 ) | ( n9162 & n9163 ) ;
  assign n9166 = ( n8838 & n9164 ) | ( n8838 & ~n9165 ) | ( n9164 & ~n9165 ) ;
  assign n9167 = ( x88 & n9161 ) | ( x88 & ~n9166 ) | ( n9161 & ~n9166 ) ;
  assign n9168 = ( x88 & n8839 ) | ( x88 & ~n9019 ) | ( n8839 & ~n9019 ) ;
  assign n9169 = x88 & n8839 ;
  assign n9170 = ( ~n8844 & n9168 ) | ( ~n8844 & n9169 ) | ( n9168 & n9169 ) ;
  assign n9171 = ( n8844 & n9168 ) | ( n8844 & n9169 ) | ( n9168 & n9169 ) ;
  assign n9172 = ( n8844 & n9170 ) | ( n8844 & ~n9171 ) | ( n9170 & ~n9171 ) ;
  assign n9173 = ( x89 & n9167 ) | ( x89 & ~n9172 ) | ( n9167 & ~n9172 ) ;
  assign n9174 = ( x89 & n8845 ) | ( x89 & ~n9019 ) | ( n8845 & ~n9019 ) ;
  assign n9175 = x89 & n8845 ;
  assign n9176 = ( ~n8850 & n9174 ) | ( ~n8850 & n9175 ) | ( n9174 & n9175 ) ;
  assign n9177 = ( n8850 & n9174 ) | ( n8850 & n9175 ) | ( n9174 & n9175 ) ;
  assign n9178 = ( n8850 & n9176 ) | ( n8850 & ~n9177 ) | ( n9176 & ~n9177 ) ;
  assign n9179 = ( x90 & n9173 ) | ( x90 & ~n9178 ) | ( n9173 & ~n9178 ) ;
  assign n9180 = ( x90 & n8851 ) | ( x90 & ~n9019 ) | ( n8851 & ~n9019 ) ;
  assign n9181 = x90 & n8851 ;
  assign n9182 = ( ~n8856 & n9180 ) | ( ~n8856 & n9181 ) | ( n9180 & n9181 ) ;
  assign n9183 = ( n8856 & n9180 ) | ( n8856 & n9181 ) | ( n9180 & n9181 ) ;
  assign n9184 = ( n8856 & n9182 ) | ( n8856 & ~n9183 ) | ( n9182 & ~n9183 ) ;
  assign n9185 = ( x91 & n9179 ) | ( x91 & ~n9184 ) | ( n9179 & ~n9184 ) ;
  assign n9186 = ( x91 & n8857 ) | ( x91 & ~n9019 ) | ( n8857 & ~n9019 ) ;
  assign n9187 = x91 & n8857 ;
  assign n9188 = ( ~n8862 & n9186 ) | ( ~n8862 & n9187 ) | ( n9186 & n9187 ) ;
  assign n9189 = ( n8862 & n9186 ) | ( n8862 & n9187 ) | ( n9186 & n9187 ) ;
  assign n9190 = ( n8862 & n9188 ) | ( n8862 & ~n9189 ) | ( n9188 & ~n9189 ) ;
  assign n9191 = ( x92 & n9185 ) | ( x92 & ~n9190 ) | ( n9185 & ~n9190 ) ;
  assign n9192 = ( x92 & n8863 ) | ( x92 & ~n9019 ) | ( n8863 & ~n9019 ) ;
  assign n9193 = x92 & n8863 ;
  assign n9194 = ( ~n8868 & n9192 ) | ( ~n8868 & n9193 ) | ( n9192 & n9193 ) ;
  assign n9195 = ( n8868 & n9192 ) | ( n8868 & n9193 ) | ( n9192 & n9193 ) ;
  assign n9196 = ( n8868 & n9194 ) | ( n8868 & ~n9195 ) | ( n9194 & ~n9195 ) ;
  assign n9197 = ( x93 & n9191 ) | ( x93 & ~n9196 ) | ( n9191 & ~n9196 ) ;
  assign n9198 = ( x93 & n8869 ) | ( x93 & ~n9019 ) | ( n8869 & ~n9019 ) ;
  assign n9199 = x93 & n8869 ;
  assign n9200 = ( ~n8874 & n9198 ) | ( ~n8874 & n9199 ) | ( n9198 & n9199 ) ;
  assign n9201 = ( n8874 & n9198 ) | ( n8874 & n9199 ) | ( n9198 & n9199 ) ;
  assign n9202 = ( n8874 & n9200 ) | ( n8874 & ~n9201 ) | ( n9200 & ~n9201 ) ;
  assign n9203 = ( x94 & n9197 ) | ( x94 & ~n9202 ) | ( n9197 & ~n9202 ) ;
  assign n9204 = ( x94 & n8875 ) | ( x94 & ~n9019 ) | ( n8875 & ~n9019 ) ;
  assign n9205 = x94 & n8875 ;
  assign n9206 = ( ~n8880 & n9204 ) | ( ~n8880 & n9205 ) | ( n9204 & n9205 ) ;
  assign n9207 = ( n8880 & n9204 ) | ( n8880 & n9205 ) | ( n9204 & n9205 ) ;
  assign n9208 = ( n8880 & n9206 ) | ( n8880 & ~n9207 ) | ( n9206 & ~n9207 ) ;
  assign n9209 = ( x95 & n9203 ) | ( x95 & ~n9208 ) | ( n9203 & ~n9208 ) ;
  assign n9210 = ( x95 & n8881 ) | ( x95 & ~n9019 ) | ( n8881 & ~n9019 ) ;
  assign n9211 = x95 & n8881 ;
  assign n9212 = ( ~n8886 & n9210 ) | ( ~n8886 & n9211 ) | ( n9210 & n9211 ) ;
  assign n9213 = ( n8886 & n9210 ) | ( n8886 & n9211 ) | ( n9210 & n9211 ) ;
  assign n9214 = ( n8886 & n9212 ) | ( n8886 & ~n9213 ) | ( n9212 & ~n9213 ) ;
  assign n9215 = ( x96 & n9209 ) | ( x96 & ~n9214 ) | ( n9209 & ~n9214 ) ;
  assign n9216 = ( x96 & n8887 ) | ( x96 & ~n9019 ) | ( n8887 & ~n9019 ) ;
  assign n9217 = x96 & n8887 ;
  assign n9218 = ( ~n8892 & n9216 ) | ( ~n8892 & n9217 ) | ( n9216 & n9217 ) ;
  assign n9219 = ( n8892 & n9216 ) | ( n8892 & n9217 ) | ( n9216 & n9217 ) ;
  assign n9220 = ( n8892 & n9218 ) | ( n8892 & ~n9219 ) | ( n9218 & ~n9219 ) ;
  assign n9221 = ( x97 & n9215 ) | ( x97 & ~n9220 ) | ( n9215 & ~n9220 ) ;
  assign n9222 = ( x97 & n8893 ) | ( x97 & ~n9019 ) | ( n8893 & ~n9019 ) ;
  assign n9223 = x97 & n8893 ;
  assign n9224 = ( ~n8898 & n9222 ) | ( ~n8898 & n9223 ) | ( n9222 & n9223 ) ;
  assign n9225 = ( n8898 & n9222 ) | ( n8898 & n9223 ) | ( n9222 & n9223 ) ;
  assign n9226 = ( n8898 & n9224 ) | ( n8898 & ~n9225 ) | ( n9224 & ~n9225 ) ;
  assign n9227 = ( x98 & n9221 ) | ( x98 & ~n9226 ) | ( n9221 & ~n9226 ) ;
  assign n9228 = ( x98 & n8899 ) | ( x98 & ~n9019 ) | ( n8899 & ~n9019 ) ;
  assign n9229 = x98 & n8899 ;
  assign n9230 = ( ~n8904 & n9228 ) | ( ~n8904 & n9229 ) | ( n9228 & n9229 ) ;
  assign n9231 = ( n8904 & n9228 ) | ( n8904 & n9229 ) | ( n9228 & n9229 ) ;
  assign n9232 = ( n8904 & n9230 ) | ( n8904 & ~n9231 ) | ( n9230 & ~n9231 ) ;
  assign n9233 = ( x99 & n9227 ) | ( x99 & ~n9232 ) | ( n9227 & ~n9232 ) ;
  assign n9234 = ( x99 & n8905 ) | ( x99 & ~n9019 ) | ( n8905 & ~n9019 ) ;
  assign n9235 = x99 & n8905 ;
  assign n9236 = ( ~n8910 & n9234 ) | ( ~n8910 & n9235 ) | ( n9234 & n9235 ) ;
  assign n9237 = ( n8910 & n9234 ) | ( n8910 & n9235 ) | ( n9234 & n9235 ) ;
  assign n9238 = ( n8910 & n9236 ) | ( n8910 & ~n9237 ) | ( n9236 & ~n9237 ) ;
  assign n9239 = ( x100 & n9233 ) | ( x100 & ~n9238 ) | ( n9233 & ~n9238 ) ;
  assign n9240 = ( x100 & n8911 ) | ( x100 & ~n9019 ) | ( n8911 & ~n9019 ) ;
  assign n9241 = x100 & n8911 ;
  assign n9242 = ( ~n8916 & n9240 ) | ( ~n8916 & n9241 ) | ( n9240 & n9241 ) ;
  assign n9243 = ( n8916 & n9240 ) | ( n8916 & n9241 ) | ( n9240 & n9241 ) ;
  assign n9244 = ( n8916 & n9242 ) | ( n8916 & ~n9243 ) | ( n9242 & ~n9243 ) ;
  assign n9245 = ( x101 & n9239 ) | ( x101 & ~n9244 ) | ( n9239 & ~n9244 ) ;
  assign n9246 = ( x101 & n8917 ) | ( x101 & ~n9019 ) | ( n8917 & ~n9019 ) ;
  assign n9247 = x101 & n8917 ;
  assign n9248 = ( ~n8922 & n9246 ) | ( ~n8922 & n9247 ) | ( n9246 & n9247 ) ;
  assign n9249 = ( n8922 & n9246 ) | ( n8922 & n9247 ) | ( n9246 & n9247 ) ;
  assign n9250 = ( n8922 & n9248 ) | ( n8922 & ~n9249 ) | ( n9248 & ~n9249 ) ;
  assign n9251 = ( x102 & n9245 ) | ( x102 & ~n9250 ) | ( n9245 & ~n9250 ) ;
  assign n9252 = ( x102 & n8923 ) | ( x102 & ~n9019 ) | ( n8923 & ~n9019 ) ;
  assign n9253 = x102 & n8923 ;
  assign n9254 = ( ~n8928 & n9252 ) | ( ~n8928 & n9253 ) | ( n9252 & n9253 ) ;
  assign n9255 = ( n8928 & n9252 ) | ( n8928 & n9253 ) | ( n9252 & n9253 ) ;
  assign n9256 = ( n8928 & n9254 ) | ( n8928 & ~n9255 ) | ( n9254 & ~n9255 ) ;
  assign n9257 = ( x103 & n9251 ) | ( x103 & ~n9256 ) | ( n9251 & ~n9256 ) ;
  assign n9258 = ( x103 & n8929 ) | ( x103 & ~n9019 ) | ( n8929 & ~n9019 ) ;
  assign n9259 = x103 & n8929 ;
  assign n9260 = ( ~n8934 & n9258 ) | ( ~n8934 & n9259 ) | ( n9258 & n9259 ) ;
  assign n9261 = ( n8934 & n9258 ) | ( n8934 & n9259 ) | ( n9258 & n9259 ) ;
  assign n9262 = ( n8934 & n9260 ) | ( n8934 & ~n9261 ) | ( n9260 & ~n9261 ) ;
  assign n9263 = ( x104 & n9257 ) | ( x104 & ~n9262 ) | ( n9257 & ~n9262 ) ;
  assign n9264 = ( x104 & n8935 ) | ( x104 & ~n9019 ) | ( n8935 & ~n9019 ) ;
  assign n9265 = x104 & n8935 ;
  assign n9266 = ( ~n8940 & n9264 ) | ( ~n8940 & n9265 ) | ( n9264 & n9265 ) ;
  assign n9267 = ( n8940 & n9264 ) | ( n8940 & n9265 ) | ( n9264 & n9265 ) ;
  assign n9268 = ( n8940 & n9266 ) | ( n8940 & ~n9267 ) | ( n9266 & ~n9267 ) ;
  assign n9269 = ( x105 & n9263 ) | ( x105 & ~n9268 ) | ( n9263 & ~n9268 ) ;
  assign n9270 = ( x105 & n8941 ) | ( x105 & ~n9019 ) | ( n8941 & ~n9019 ) ;
  assign n9271 = x105 & n8941 ;
  assign n9272 = ( ~n8946 & n9270 ) | ( ~n8946 & n9271 ) | ( n9270 & n9271 ) ;
  assign n9273 = ( n8946 & n9270 ) | ( n8946 & n9271 ) | ( n9270 & n9271 ) ;
  assign n9274 = ( n8946 & n9272 ) | ( n8946 & ~n9273 ) | ( n9272 & ~n9273 ) ;
  assign n9275 = ( x106 & n9269 ) | ( x106 & ~n9274 ) | ( n9269 & ~n9274 ) ;
  assign n9276 = ( x106 & n8947 ) | ( x106 & ~n9019 ) | ( n8947 & ~n9019 ) ;
  assign n9277 = x106 & n8947 ;
  assign n9278 = ( ~n8952 & n9276 ) | ( ~n8952 & n9277 ) | ( n9276 & n9277 ) ;
  assign n9279 = ( n8952 & n9276 ) | ( n8952 & n9277 ) | ( n9276 & n9277 ) ;
  assign n9280 = ( n8952 & n9278 ) | ( n8952 & ~n9279 ) | ( n9278 & ~n9279 ) ;
  assign n9281 = ( x107 & n9275 ) | ( x107 & ~n9280 ) | ( n9275 & ~n9280 ) ;
  assign n9282 = ( x107 & n8953 ) | ( x107 & ~n9019 ) | ( n8953 & ~n9019 ) ;
  assign n9283 = x107 & n8953 ;
  assign n9284 = ( ~n8958 & n9282 ) | ( ~n8958 & n9283 ) | ( n9282 & n9283 ) ;
  assign n9285 = ( n8958 & n9282 ) | ( n8958 & n9283 ) | ( n9282 & n9283 ) ;
  assign n9286 = ( n8958 & n9284 ) | ( n8958 & ~n9285 ) | ( n9284 & ~n9285 ) ;
  assign n9287 = ( x108 & n9281 ) | ( x108 & ~n9286 ) | ( n9281 & ~n9286 ) ;
  assign n9288 = ( x108 & n8959 ) | ( x108 & ~n9019 ) | ( n8959 & ~n9019 ) ;
  assign n9289 = x108 & n8959 ;
  assign n9290 = ( ~n8964 & n9288 ) | ( ~n8964 & n9289 ) | ( n9288 & n9289 ) ;
  assign n9291 = ( n8964 & n9288 ) | ( n8964 & n9289 ) | ( n9288 & n9289 ) ;
  assign n9292 = ( n8964 & n9290 ) | ( n8964 & ~n9291 ) | ( n9290 & ~n9291 ) ;
  assign n9293 = ( x109 & n9287 ) | ( x109 & ~n9292 ) | ( n9287 & ~n9292 ) ;
  assign n9294 = ( x109 & n8965 ) | ( x109 & ~n9019 ) | ( n8965 & ~n9019 ) ;
  assign n9295 = x109 & n8965 ;
  assign n9296 = ( ~n8970 & n9294 ) | ( ~n8970 & n9295 ) | ( n9294 & n9295 ) ;
  assign n9297 = ( n8970 & n9294 ) | ( n8970 & n9295 ) | ( n9294 & n9295 ) ;
  assign n9298 = ( n8970 & n9296 ) | ( n8970 & ~n9297 ) | ( n9296 & ~n9297 ) ;
  assign n9299 = ( x110 & n9293 ) | ( x110 & ~n9298 ) | ( n9293 & ~n9298 ) ;
  assign n9300 = ( x110 & n8971 ) | ( x110 & ~n9019 ) | ( n8971 & ~n9019 ) ;
  assign n9301 = x110 & n8971 ;
  assign n9302 = ( ~n8976 & n9300 ) | ( ~n8976 & n9301 ) | ( n9300 & n9301 ) ;
  assign n9303 = ( n8976 & n9300 ) | ( n8976 & n9301 ) | ( n9300 & n9301 ) ;
  assign n9304 = ( n8976 & n9302 ) | ( n8976 & ~n9303 ) | ( n9302 & ~n9303 ) ;
  assign n9305 = ( x111 & n9299 ) | ( x111 & ~n9304 ) | ( n9299 & ~n9304 ) ;
  assign n9306 = ( x111 & n8977 ) | ( x111 & ~n9019 ) | ( n8977 & ~n9019 ) ;
  assign n9307 = x111 & n8977 ;
  assign n9308 = ( ~n8982 & n9306 ) | ( ~n8982 & n9307 ) | ( n9306 & n9307 ) ;
  assign n9309 = ( n8982 & n9306 ) | ( n8982 & n9307 ) | ( n9306 & n9307 ) ;
  assign n9310 = ( n8982 & n9308 ) | ( n8982 & ~n9309 ) | ( n9308 & ~n9309 ) ;
  assign n9311 = ( x112 & n9305 ) | ( x112 & ~n9310 ) | ( n9305 & ~n9310 ) ;
  assign n9312 = ( x112 & n8983 ) | ( x112 & ~n9019 ) | ( n8983 & ~n9019 ) ;
  assign n9313 = x112 & n8983 ;
  assign n9314 = ( ~n8988 & n9312 ) | ( ~n8988 & n9313 ) | ( n9312 & n9313 ) ;
  assign n9315 = ( n8988 & n9312 ) | ( n8988 & n9313 ) | ( n9312 & n9313 ) ;
  assign n9316 = ( n8988 & n9314 ) | ( n8988 & ~n9315 ) | ( n9314 & ~n9315 ) ;
  assign n9317 = ( x113 & n9311 ) | ( x113 & ~n9316 ) | ( n9311 & ~n9316 ) ;
  assign n9318 = ( x113 & n8989 ) | ( x113 & ~n9019 ) | ( n8989 & ~n9019 ) ;
  assign n9319 = x113 & n8989 ;
  assign n9320 = ( ~n8994 & n9318 ) | ( ~n8994 & n9319 ) | ( n9318 & n9319 ) ;
  assign n9321 = ( n8994 & n9318 ) | ( n8994 & n9319 ) | ( n9318 & n9319 ) ;
  assign n9322 = ( n8994 & n9320 ) | ( n8994 & ~n9321 ) | ( n9320 & ~n9321 ) ;
  assign n9323 = ( x114 & n9317 ) | ( x114 & ~n9322 ) | ( n9317 & ~n9322 ) ;
  assign n9324 = ( x114 & n8995 ) | ( x114 & ~n9019 ) | ( n8995 & ~n9019 ) ;
  assign n9325 = x114 & n8995 ;
  assign n9326 = ( ~n9000 & n9324 ) | ( ~n9000 & n9325 ) | ( n9324 & n9325 ) ;
  assign n9327 = ( n9000 & n9324 ) | ( n9000 & n9325 ) | ( n9324 & n9325 ) ;
  assign n9328 = ( n9000 & n9326 ) | ( n9000 & ~n9327 ) | ( n9326 & ~n9327 ) ;
  assign n9329 = ( x115 & n9323 ) | ( x115 & ~n9328 ) | ( n9323 & ~n9328 ) ;
  assign n9330 = ( x115 & n9001 ) | ( x115 & ~n9019 ) | ( n9001 & ~n9019 ) ;
  assign n9331 = x115 & n9001 ;
  assign n9332 = ( ~n9006 & n9330 ) | ( ~n9006 & n9331 ) | ( n9330 & n9331 ) ;
  assign n9333 = ( n9006 & n9330 ) | ( n9006 & n9331 ) | ( n9330 & n9331 ) ;
  assign n9334 = ( n9006 & n9332 ) | ( n9006 & ~n9333 ) | ( n9332 & ~n9333 ) ;
  assign n9335 = ( x116 & n9329 ) | ( x116 & ~n9334 ) | ( n9329 & ~n9334 ) ;
  assign n9336 = ( x116 & n9007 ) | ( x116 & ~n9019 ) | ( n9007 & ~n9019 ) ;
  assign n9337 = x116 & n9007 ;
  assign n9338 = ( ~n9012 & n9336 ) | ( ~n9012 & n9337 ) | ( n9336 & n9337 ) ;
  assign n9339 = ( n9012 & n9336 ) | ( n9012 & n9337 ) | ( n9336 & n9337 ) ;
  assign n9340 = ( n9012 & n9338 ) | ( n9012 & ~n9339 ) | ( n9338 & ~n9339 ) ;
  assign n9341 = ( x117 & n9335 ) | ( x117 & ~n9340 ) | ( n9335 & ~n9340 ) ;
  assign n9342 = ( x118 & ~n9024 ) | ( x118 & n9341 ) | ( ~n9024 & n9341 ) ;
  assign n9343 = ( n137 & n138 ) | ( n137 & ~n8695 ) | ( n138 & ~n8695 ) ;
  assign n9344 = ( n138 & n139 ) | ( n138 & ~n9017 ) | ( n139 & ~n9017 ) ;
  assign n9345 = ( x118 & n9016 ) | ( x118 & ~n9017 ) | ( n9016 & ~n9017 ) ;
  assign n9346 = ~n9344 & n9345 ;
  assign n9347 = ( n9342 & n9343 ) | ( n9342 & ~n9346 ) | ( n9343 & ~n9346 ) ;
  assign n9348 = ( x118 & n9341 ) | ( x118 & n9347 ) | ( n9341 & n9347 ) ;
  assign n9349 = x118 | n9341 ;
  assign n9350 = ( ~n9024 & n9348 ) | ( ~n9024 & n9349 ) | ( n9348 & n9349 ) ;
  assign n9351 = ( n9024 & n9348 ) | ( n9024 & n9349 ) | ( n9348 & n9349 ) ;
  assign n9352 = ( n9024 & n9350 ) | ( n9024 & ~n9351 ) | ( n9350 & ~n9351 ) ;
  assign n9353 = ~x7 & x64 ;
  assign n9354 = ~x8 & n9347 ;
  assign n9355 = ( x8 & ~x64 ) | ( x8 & n9347 ) | ( ~x64 & n9347 ) ;
  assign n9356 = ( n9025 & ~n9354 ) | ( n9025 & n9355 ) | ( ~n9354 & n9355 ) ;
  assign n9357 = ( x65 & n9353 ) | ( x65 & ~n9356 ) | ( n9353 & ~n9356 ) ;
  assign n9358 = ( x65 & n9025 ) | ( x65 & n9347 ) | ( n9025 & n9347 ) ;
  assign n9359 = x65 | n9025 ;
  assign n9360 = ( ~n9028 & n9358 ) | ( ~n9028 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9361 = ( n9028 & n9358 ) | ( n9028 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9362 = ( n9028 & n9360 ) | ( n9028 & ~n9361 ) | ( n9360 & ~n9361 ) ;
  assign n9363 = ( x66 & n9357 ) | ( x66 & ~n9362 ) | ( n9357 & ~n9362 ) ;
  assign n9364 = ( x66 & n9029 ) | ( x66 & n9347 ) | ( n9029 & n9347 ) ;
  assign n9365 = x66 | n9029 ;
  assign n9366 = ( ~n9034 & n9364 ) | ( ~n9034 & n9365 ) | ( n9364 & n9365 ) ;
  assign n9367 = ( n9034 & n9364 ) | ( n9034 & n9365 ) | ( n9364 & n9365 ) ;
  assign n9368 = ( n9034 & n9366 ) | ( n9034 & ~n9367 ) | ( n9366 & ~n9367 ) ;
  assign n9369 = ( x67 & n9363 ) | ( x67 & ~n9368 ) | ( n9363 & ~n9368 ) ;
  assign n9370 = ( x67 & n9035 ) | ( x67 & ~n9347 ) | ( n9035 & ~n9347 ) ;
  assign n9371 = x67 & n9035 ;
  assign n9372 = ( ~n9040 & n9370 ) | ( ~n9040 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9373 = ( n9040 & n9370 ) | ( n9040 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9374 = ( n9040 & n9372 ) | ( n9040 & ~n9373 ) | ( n9372 & ~n9373 ) ;
  assign n9375 = ( x68 & n9369 ) | ( x68 & ~n9374 ) | ( n9369 & ~n9374 ) ;
  assign n9376 = ( x68 & n9041 ) | ( x68 & ~n9347 ) | ( n9041 & ~n9347 ) ;
  assign n9377 = x68 & n9041 ;
  assign n9378 = ( ~n9046 & n9376 ) | ( ~n9046 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9379 = ( n9046 & n9376 ) | ( n9046 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9380 = ( n9046 & n9378 ) | ( n9046 & ~n9379 ) | ( n9378 & ~n9379 ) ;
  assign n9381 = ( x69 & n9375 ) | ( x69 & ~n9380 ) | ( n9375 & ~n9380 ) ;
  assign n9382 = ( x69 & n9047 ) | ( x69 & ~n9347 ) | ( n9047 & ~n9347 ) ;
  assign n9383 = x69 & n9047 ;
  assign n9384 = ( ~n9052 & n9382 ) | ( ~n9052 & n9383 ) | ( n9382 & n9383 ) ;
  assign n9385 = ( n9052 & n9382 ) | ( n9052 & n9383 ) | ( n9382 & n9383 ) ;
  assign n9386 = ( n9052 & n9384 ) | ( n9052 & ~n9385 ) | ( n9384 & ~n9385 ) ;
  assign n9387 = ( x70 & n9381 ) | ( x70 & ~n9386 ) | ( n9381 & ~n9386 ) ;
  assign n9388 = ( x70 & n9053 ) | ( x70 & ~n9347 ) | ( n9053 & ~n9347 ) ;
  assign n9389 = x70 & n9053 ;
  assign n9390 = ( ~n9058 & n9388 ) | ( ~n9058 & n9389 ) | ( n9388 & n9389 ) ;
  assign n9391 = ( n9058 & n9388 ) | ( n9058 & n9389 ) | ( n9388 & n9389 ) ;
  assign n9392 = ( n9058 & n9390 ) | ( n9058 & ~n9391 ) | ( n9390 & ~n9391 ) ;
  assign n9393 = ( x71 & n9387 ) | ( x71 & ~n9392 ) | ( n9387 & ~n9392 ) ;
  assign n9394 = ( x71 & n9059 ) | ( x71 & ~n9347 ) | ( n9059 & ~n9347 ) ;
  assign n9395 = x71 & n9059 ;
  assign n9396 = ( ~n9064 & n9394 ) | ( ~n9064 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9397 = ( n9064 & n9394 ) | ( n9064 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9398 = ( n9064 & n9396 ) | ( n9064 & ~n9397 ) | ( n9396 & ~n9397 ) ;
  assign n9399 = ( x72 & n9393 ) | ( x72 & ~n9398 ) | ( n9393 & ~n9398 ) ;
  assign n9400 = ( x72 & n9065 ) | ( x72 & ~n9347 ) | ( n9065 & ~n9347 ) ;
  assign n9401 = x72 & n9065 ;
  assign n9402 = ( ~n9070 & n9400 ) | ( ~n9070 & n9401 ) | ( n9400 & n9401 ) ;
  assign n9403 = ( n9070 & n9400 ) | ( n9070 & n9401 ) | ( n9400 & n9401 ) ;
  assign n9404 = ( n9070 & n9402 ) | ( n9070 & ~n9403 ) | ( n9402 & ~n9403 ) ;
  assign n9405 = ( x73 & n9399 ) | ( x73 & ~n9404 ) | ( n9399 & ~n9404 ) ;
  assign n9406 = ( x73 & n9071 ) | ( x73 & ~n9347 ) | ( n9071 & ~n9347 ) ;
  assign n9407 = x73 & n9071 ;
  assign n9408 = ( ~n9076 & n9406 ) | ( ~n9076 & n9407 ) | ( n9406 & n9407 ) ;
  assign n9409 = ( n9076 & n9406 ) | ( n9076 & n9407 ) | ( n9406 & n9407 ) ;
  assign n9410 = ( n9076 & n9408 ) | ( n9076 & ~n9409 ) | ( n9408 & ~n9409 ) ;
  assign n9411 = ( x74 & n9405 ) | ( x74 & ~n9410 ) | ( n9405 & ~n9410 ) ;
  assign n9412 = ( x74 & n9077 ) | ( x74 & ~n9347 ) | ( n9077 & ~n9347 ) ;
  assign n9413 = x74 & n9077 ;
  assign n9414 = ( ~n9082 & n9412 ) | ( ~n9082 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9415 = ( n9082 & n9412 ) | ( n9082 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9416 = ( n9082 & n9414 ) | ( n9082 & ~n9415 ) | ( n9414 & ~n9415 ) ;
  assign n9417 = ( x75 & n9411 ) | ( x75 & ~n9416 ) | ( n9411 & ~n9416 ) ;
  assign n9418 = ( x75 & n9083 ) | ( x75 & ~n9347 ) | ( n9083 & ~n9347 ) ;
  assign n9419 = x75 & n9083 ;
  assign n9420 = ( ~n9088 & n9418 ) | ( ~n9088 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = ( n9088 & n9418 ) | ( n9088 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9422 = ( n9088 & n9420 ) | ( n9088 & ~n9421 ) | ( n9420 & ~n9421 ) ;
  assign n9423 = ( x76 & n9417 ) | ( x76 & ~n9422 ) | ( n9417 & ~n9422 ) ;
  assign n9424 = ( x76 & n9089 ) | ( x76 & ~n9347 ) | ( n9089 & ~n9347 ) ;
  assign n9425 = x76 & n9089 ;
  assign n9426 = ( ~n9094 & n9424 ) | ( ~n9094 & n9425 ) | ( n9424 & n9425 ) ;
  assign n9427 = ( n9094 & n9424 ) | ( n9094 & n9425 ) | ( n9424 & n9425 ) ;
  assign n9428 = ( n9094 & n9426 ) | ( n9094 & ~n9427 ) | ( n9426 & ~n9427 ) ;
  assign n9429 = ( x77 & n9423 ) | ( x77 & ~n9428 ) | ( n9423 & ~n9428 ) ;
  assign n9430 = ( x77 & n9095 ) | ( x77 & ~n9347 ) | ( n9095 & ~n9347 ) ;
  assign n9431 = x77 & n9095 ;
  assign n9432 = ( ~n9100 & n9430 ) | ( ~n9100 & n9431 ) | ( n9430 & n9431 ) ;
  assign n9433 = ( n9100 & n9430 ) | ( n9100 & n9431 ) | ( n9430 & n9431 ) ;
  assign n9434 = ( n9100 & n9432 ) | ( n9100 & ~n9433 ) | ( n9432 & ~n9433 ) ;
  assign n9435 = ( x78 & n9429 ) | ( x78 & ~n9434 ) | ( n9429 & ~n9434 ) ;
  assign n9436 = ( x78 & n9101 ) | ( x78 & ~n9347 ) | ( n9101 & ~n9347 ) ;
  assign n9437 = x78 & n9101 ;
  assign n9438 = ( ~n9106 & n9436 ) | ( ~n9106 & n9437 ) | ( n9436 & n9437 ) ;
  assign n9439 = ( n9106 & n9436 ) | ( n9106 & n9437 ) | ( n9436 & n9437 ) ;
  assign n9440 = ( n9106 & n9438 ) | ( n9106 & ~n9439 ) | ( n9438 & ~n9439 ) ;
  assign n9441 = ( x79 & n9435 ) | ( x79 & ~n9440 ) | ( n9435 & ~n9440 ) ;
  assign n9442 = ( x79 & n9107 ) | ( x79 & ~n9347 ) | ( n9107 & ~n9347 ) ;
  assign n9443 = x79 & n9107 ;
  assign n9444 = ( ~n9112 & n9442 ) | ( ~n9112 & n9443 ) | ( n9442 & n9443 ) ;
  assign n9445 = ( n9112 & n9442 ) | ( n9112 & n9443 ) | ( n9442 & n9443 ) ;
  assign n9446 = ( n9112 & n9444 ) | ( n9112 & ~n9445 ) | ( n9444 & ~n9445 ) ;
  assign n9447 = ( x80 & n9441 ) | ( x80 & ~n9446 ) | ( n9441 & ~n9446 ) ;
  assign n9448 = ( x80 & n9113 ) | ( x80 & ~n9347 ) | ( n9113 & ~n9347 ) ;
  assign n9449 = x80 & n9113 ;
  assign n9450 = ( ~n9118 & n9448 ) | ( ~n9118 & n9449 ) | ( n9448 & n9449 ) ;
  assign n9451 = ( n9118 & n9448 ) | ( n9118 & n9449 ) | ( n9448 & n9449 ) ;
  assign n9452 = ( n9118 & n9450 ) | ( n9118 & ~n9451 ) | ( n9450 & ~n9451 ) ;
  assign n9453 = ( x81 & n9447 ) | ( x81 & ~n9452 ) | ( n9447 & ~n9452 ) ;
  assign n9454 = ( x81 & n9119 ) | ( x81 & ~n9347 ) | ( n9119 & ~n9347 ) ;
  assign n9455 = x81 & n9119 ;
  assign n9456 = ( ~n9124 & n9454 ) | ( ~n9124 & n9455 ) | ( n9454 & n9455 ) ;
  assign n9457 = ( n9124 & n9454 ) | ( n9124 & n9455 ) | ( n9454 & n9455 ) ;
  assign n9458 = ( n9124 & n9456 ) | ( n9124 & ~n9457 ) | ( n9456 & ~n9457 ) ;
  assign n9459 = ( x82 & n9453 ) | ( x82 & ~n9458 ) | ( n9453 & ~n9458 ) ;
  assign n9460 = ( x82 & n9125 ) | ( x82 & ~n9347 ) | ( n9125 & ~n9347 ) ;
  assign n9461 = x82 & n9125 ;
  assign n9462 = ( ~n9130 & n9460 ) | ( ~n9130 & n9461 ) | ( n9460 & n9461 ) ;
  assign n9463 = ( n9130 & n9460 ) | ( n9130 & n9461 ) | ( n9460 & n9461 ) ;
  assign n9464 = ( n9130 & n9462 ) | ( n9130 & ~n9463 ) | ( n9462 & ~n9463 ) ;
  assign n9465 = ( x83 & n9459 ) | ( x83 & ~n9464 ) | ( n9459 & ~n9464 ) ;
  assign n9466 = ( x83 & n9131 ) | ( x83 & ~n9347 ) | ( n9131 & ~n9347 ) ;
  assign n9467 = x83 & n9131 ;
  assign n9468 = ( ~n9136 & n9466 ) | ( ~n9136 & n9467 ) | ( n9466 & n9467 ) ;
  assign n9469 = ( n9136 & n9466 ) | ( n9136 & n9467 ) | ( n9466 & n9467 ) ;
  assign n9470 = ( n9136 & n9468 ) | ( n9136 & ~n9469 ) | ( n9468 & ~n9469 ) ;
  assign n9471 = ( x84 & n9465 ) | ( x84 & ~n9470 ) | ( n9465 & ~n9470 ) ;
  assign n9472 = ( x84 & n9137 ) | ( x84 & ~n9347 ) | ( n9137 & ~n9347 ) ;
  assign n9473 = x84 & n9137 ;
  assign n9474 = ( ~n9142 & n9472 ) | ( ~n9142 & n9473 ) | ( n9472 & n9473 ) ;
  assign n9475 = ( n9142 & n9472 ) | ( n9142 & n9473 ) | ( n9472 & n9473 ) ;
  assign n9476 = ( n9142 & n9474 ) | ( n9142 & ~n9475 ) | ( n9474 & ~n9475 ) ;
  assign n9477 = ( x85 & n9471 ) | ( x85 & ~n9476 ) | ( n9471 & ~n9476 ) ;
  assign n9478 = ( x85 & n9143 ) | ( x85 & ~n9347 ) | ( n9143 & ~n9347 ) ;
  assign n9479 = x85 & n9143 ;
  assign n9480 = ( ~n9148 & n9478 ) | ( ~n9148 & n9479 ) | ( n9478 & n9479 ) ;
  assign n9481 = ( n9148 & n9478 ) | ( n9148 & n9479 ) | ( n9478 & n9479 ) ;
  assign n9482 = ( n9148 & n9480 ) | ( n9148 & ~n9481 ) | ( n9480 & ~n9481 ) ;
  assign n9483 = ( x86 & n9477 ) | ( x86 & ~n9482 ) | ( n9477 & ~n9482 ) ;
  assign n9484 = ( x86 & n9149 ) | ( x86 & ~n9347 ) | ( n9149 & ~n9347 ) ;
  assign n9485 = x86 & n9149 ;
  assign n9486 = ( ~n9154 & n9484 ) | ( ~n9154 & n9485 ) | ( n9484 & n9485 ) ;
  assign n9487 = ( n9154 & n9484 ) | ( n9154 & n9485 ) | ( n9484 & n9485 ) ;
  assign n9488 = ( n9154 & n9486 ) | ( n9154 & ~n9487 ) | ( n9486 & ~n9487 ) ;
  assign n9489 = ( x87 & n9483 ) | ( x87 & ~n9488 ) | ( n9483 & ~n9488 ) ;
  assign n9490 = ( x87 & n9155 ) | ( x87 & ~n9347 ) | ( n9155 & ~n9347 ) ;
  assign n9491 = x87 & n9155 ;
  assign n9492 = ( ~n9160 & n9490 ) | ( ~n9160 & n9491 ) | ( n9490 & n9491 ) ;
  assign n9493 = ( n9160 & n9490 ) | ( n9160 & n9491 ) | ( n9490 & n9491 ) ;
  assign n9494 = ( n9160 & n9492 ) | ( n9160 & ~n9493 ) | ( n9492 & ~n9493 ) ;
  assign n9495 = ( x88 & n9489 ) | ( x88 & ~n9494 ) | ( n9489 & ~n9494 ) ;
  assign n9496 = ( x88 & n9161 ) | ( x88 & ~n9347 ) | ( n9161 & ~n9347 ) ;
  assign n9497 = x88 & n9161 ;
  assign n9498 = ( ~n9166 & n9496 ) | ( ~n9166 & n9497 ) | ( n9496 & n9497 ) ;
  assign n9499 = ( n9166 & n9496 ) | ( n9166 & n9497 ) | ( n9496 & n9497 ) ;
  assign n9500 = ( n9166 & n9498 ) | ( n9166 & ~n9499 ) | ( n9498 & ~n9499 ) ;
  assign n9501 = ( x89 & n9495 ) | ( x89 & ~n9500 ) | ( n9495 & ~n9500 ) ;
  assign n9502 = ( x89 & n9167 ) | ( x89 & ~n9347 ) | ( n9167 & ~n9347 ) ;
  assign n9503 = x89 & n9167 ;
  assign n9504 = ( ~n9172 & n9502 ) | ( ~n9172 & n9503 ) | ( n9502 & n9503 ) ;
  assign n9505 = ( n9172 & n9502 ) | ( n9172 & n9503 ) | ( n9502 & n9503 ) ;
  assign n9506 = ( n9172 & n9504 ) | ( n9172 & ~n9505 ) | ( n9504 & ~n9505 ) ;
  assign n9507 = ( x90 & n9501 ) | ( x90 & ~n9506 ) | ( n9501 & ~n9506 ) ;
  assign n9508 = ( x90 & n9173 ) | ( x90 & ~n9347 ) | ( n9173 & ~n9347 ) ;
  assign n9509 = x90 & n9173 ;
  assign n9510 = ( ~n9178 & n9508 ) | ( ~n9178 & n9509 ) | ( n9508 & n9509 ) ;
  assign n9511 = ( n9178 & n9508 ) | ( n9178 & n9509 ) | ( n9508 & n9509 ) ;
  assign n9512 = ( n9178 & n9510 ) | ( n9178 & ~n9511 ) | ( n9510 & ~n9511 ) ;
  assign n9513 = ( x91 & n9507 ) | ( x91 & ~n9512 ) | ( n9507 & ~n9512 ) ;
  assign n9514 = ( x91 & n9179 ) | ( x91 & ~n9347 ) | ( n9179 & ~n9347 ) ;
  assign n9515 = x91 & n9179 ;
  assign n9516 = ( ~n9184 & n9514 ) | ( ~n9184 & n9515 ) | ( n9514 & n9515 ) ;
  assign n9517 = ( n9184 & n9514 ) | ( n9184 & n9515 ) | ( n9514 & n9515 ) ;
  assign n9518 = ( n9184 & n9516 ) | ( n9184 & ~n9517 ) | ( n9516 & ~n9517 ) ;
  assign n9519 = ( x92 & n9513 ) | ( x92 & ~n9518 ) | ( n9513 & ~n9518 ) ;
  assign n9520 = ( x92 & n9185 ) | ( x92 & ~n9347 ) | ( n9185 & ~n9347 ) ;
  assign n9521 = x92 & n9185 ;
  assign n9522 = ( ~n9190 & n9520 ) | ( ~n9190 & n9521 ) | ( n9520 & n9521 ) ;
  assign n9523 = ( n9190 & n9520 ) | ( n9190 & n9521 ) | ( n9520 & n9521 ) ;
  assign n9524 = ( n9190 & n9522 ) | ( n9190 & ~n9523 ) | ( n9522 & ~n9523 ) ;
  assign n9525 = ( x93 & n9519 ) | ( x93 & ~n9524 ) | ( n9519 & ~n9524 ) ;
  assign n9526 = ( x93 & n9191 ) | ( x93 & ~n9347 ) | ( n9191 & ~n9347 ) ;
  assign n9527 = x93 & n9191 ;
  assign n9528 = ( ~n9196 & n9526 ) | ( ~n9196 & n9527 ) | ( n9526 & n9527 ) ;
  assign n9529 = ( n9196 & n9526 ) | ( n9196 & n9527 ) | ( n9526 & n9527 ) ;
  assign n9530 = ( n9196 & n9528 ) | ( n9196 & ~n9529 ) | ( n9528 & ~n9529 ) ;
  assign n9531 = ( x94 & n9525 ) | ( x94 & ~n9530 ) | ( n9525 & ~n9530 ) ;
  assign n9532 = ( x94 & n9197 ) | ( x94 & ~n9347 ) | ( n9197 & ~n9347 ) ;
  assign n9533 = x94 & n9197 ;
  assign n9534 = ( ~n9202 & n9532 ) | ( ~n9202 & n9533 ) | ( n9532 & n9533 ) ;
  assign n9535 = ( n9202 & n9532 ) | ( n9202 & n9533 ) | ( n9532 & n9533 ) ;
  assign n9536 = ( n9202 & n9534 ) | ( n9202 & ~n9535 ) | ( n9534 & ~n9535 ) ;
  assign n9537 = ( x95 & n9531 ) | ( x95 & ~n9536 ) | ( n9531 & ~n9536 ) ;
  assign n9538 = ( x95 & n9203 ) | ( x95 & ~n9347 ) | ( n9203 & ~n9347 ) ;
  assign n9539 = x95 & n9203 ;
  assign n9540 = ( ~n9208 & n9538 ) | ( ~n9208 & n9539 ) | ( n9538 & n9539 ) ;
  assign n9541 = ( n9208 & n9538 ) | ( n9208 & n9539 ) | ( n9538 & n9539 ) ;
  assign n9542 = ( n9208 & n9540 ) | ( n9208 & ~n9541 ) | ( n9540 & ~n9541 ) ;
  assign n9543 = ( x96 & n9537 ) | ( x96 & ~n9542 ) | ( n9537 & ~n9542 ) ;
  assign n9544 = ( x96 & n9209 ) | ( x96 & ~n9347 ) | ( n9209 & ~n9347 ) ;
  assign n9545 = x96 & n9209 ;
  assign n9546 = ( ~n9214 & n9544 ) | ( ~n9214 & n9545 ) | ( n9544 & n9545 ) ;
  assign n9547 = ( n9214 & n9544 ) | ( n9214 & n9545 ) | ( n9544 & n9545 ) ;
  assign n9548 = ( n9214 & n9546 ) | ( n9214 & ~n9547 ) | ( n9546 & ~n9547 ) ;
  assign n9549 = ( x97 & n9543 ) | ( x97 & ~n9548 ) | ( n9543 & ~n9548 ) ;
  assign n9550 = ( x97 & n9215 ) | ( x97 & ~n9347 ) | ( n9215 & ~n9347 ) ;
  assign n9551 = x97 & n9215 ;
  assign n9552 = ( ~n9220 & n9550 ) | ( ~n9220 & n9551 ) | ( n9550 & n9551 ) ;
  assign n9553 = ( n9220 & n9550 ) | ( n9220 & n9551 ) | ( n9550 & n9551 ) ;
  assign n9554 = ( n9220 & n9552 ) | ( n9220 & ~n9553 ) | ( n9552 & ~n9553 ) ;
  assign n9555 = ( x98 & n9549 ) | ( x98 & ~n9554 ) | ( n9549 & ~n9554 ) ;
  assign n9556 = ( x98 & n9221 ) | ( x98 & ~n9347 ) | ( n9221 & ~n9347 ) ;
  assign n9557 = x98 & n9221 ;
  assign n9558 = ( ~n9226 & n9556 ) | ( ~n9226 & n9557 ) | ( n9556 & n9557 ) ;
  assign n9559 = ( n9226 & n9556 ) | ( n9226 & n9557 ) | ( n9556 & n9557 ) ;
  assign n9560 = ( n9226 & n9558 ) | ( n9226 & ~n9559 ) | ( n9558 & ~n9559 ) ;
  assign n9561 = ( x99 & n9555 ) | ( x99 & ~n9560 ) | ( n9555 & ~n9560 ) ;
  assign n9562 = ( x99 & n9227 ) | ( x99 & ~n9347 ) | ( n9227 & ~n9347 ) ;
  assign n9563 = x99 & n9227 ;
  assign n9564 = ( ~n9232 & n9562 ) | ( ~n9232 & n9563 ) | ( n9562 & n9563 ) ;
  assign n9565 = ( n9232 & n9562 ) | ( n9232 & n9563 ) | ( n9562 & n9563 ) ;
  assign n9566 = ( n9232 & n9564 ) | ( n9232 & ~n9565 ) | ( n9564 & ~n9565 ) ;
  assign n9567 = ( x100 & n9561 ) | ( x100 & ~n9566 ) | ( n9561 & ~n9566 ) ;
  assign n9568 = ( x100 & n9233 ) | ( x100 & ~n9347 ) | ( n9233 & ~n9347 ) ;
  assign n9569 = x100 & n9233 ;
  assign n9570 = ( ~n9238 & n9568 ) | ( ~n9238 & n9569 ) | ( n9568 & n9569 ) ;
  assign n9571 = ( n9238 & n9568 ) | ( n9238 & n9569 ) | ( n9568 & n9569 ) ;
  assign n9572 = ( n9238 & n9570 ) | ( n9238 & ~n9571 ) | ( n9570 & ~n9571 ) ;
  assign n9573 = ( x101 & n9567 ) | ( x101 & ~n9572 ) | ( n9567 & ~n9572 ) ;
  assign n9574 = ( x101 & n9239 ) | ( x101 & ~n9347 ) | ( n9239 & ~n9347 ) ;
  assign n9575 = x101 & n9239 ;
  assign n9576 = ( ~n9244 & n9574 ) | ( ~n9244 & n9575 ) | ( n9574 & n9575 ) ;
  assign n9577 = ( n9244 & n9574 ) | ( n9244 & n9575 ) | ( n9574 & n9575 ) ;
  assign n9578 = ( n9244 & n9576 ) | ( n9244 & ~n9577 ) | ( n9576 & ~n9577 ) ;
  assign n9579 = ( x102 & n9573 ) | ( x102 & ~n9578 ) | ( n9573 & ~n9578 ) ;
  assign n9580 = ( x102 & n9245 ) | ( x102 & ~n9347 ) | ( n9245 & ~n9347 ) ;
  assign n9581 = x102 & n9245 ;
  assign n9582 = ( ~n9250 & n9580 ) | ( ~n9250 & n9581 ) | ( n9580 & n9581 ) ;
  assign n9583 = ( n9250 & n9580 ) | ( n9250 & n9581 ) | ( n9580 & n9581 ) ;
  assign n9584 = ( n9250 & n9582 ) | ( n9250 & ~n9583 ) | ( n9582 & ~n9583 ) ;
  assign n9585 = ( x103 & n9579 ) | ( x103 & ~n9584 ) | ( n9579 & ~n9584 ) ;
  assign n9586 = ( x103 & n9251 ) | ( x103 & ~n9347 ) | ( n9251 & ~n9347 ) ;
  assign n9587 = x103 & n9251 ;
  assign n9588 = ( ~n9256 & n9586 ) | ( ~n9256 & n9587 ) | ( n9586 & n9587 ) ;
  assign n9589 = ( n9256 & n9586 ) | ( n9256 & n9587 ) | ( n9586 & n9587 ) ;
  assign n9590 = ( n9256 & n9588 ) | ( n9256 & ~n9589 ) | ( n9588 & ~n9589 ) ;
  assign n9591 = ( x104 & n9585 ) | ( x104 & ~n9590 ) | ( n9585 & ~n9590 ) ;
  assign n9592 = ( x104 & n9257 ) | ( x104 & ~n9347 ) | ( n9257 & ~n9347 ) ;
  assign n9593 = x104 & n9257 ;
  assign n9594 = ( ~n9262 & n9592 ) | ( ~n9262 & n9593 ) | ( n9592 & n9593 ) ;
  assign n9595 = ( n9262 & n9592 ) | ( n9262 & n9593 ) | ( n9592 & n9593 ) ;
  assign n9596 = ( n9262 & n9594 ) | ( n9262 & ~n9595 ) | ( n9594 & ~n9595 ) ;
  assign n9597 = ( x105 & n9591 ) | ( x105 & ~n9596 ) | ( n9591 & ~n9596 ) ;
  assign n9598 = ( x105 & n9263 ) | ( x105 & ~n9347 ) | ( n9263 & ~n9347 ) ;
  assign n9599 = x105 & n9263 ;
  assign n9600 = ( ~n9268 & n9598 ) | ( ~n9268 & n9599 ) | ( n9598 & n9599 ) ;
  assign n9601 = ( n9268 & n9598 ) | ( n9268 & n9599 ) | ( n9598 & n9599 ) ;
  assign n9602 = ( n9268 & n9600 ) | ( n9268 & ~n9601 ) | ( n9600 & ~n9601 ) ;
  assign n9603 = ( x106 & n9597 ) | ( x106 & ~n9602 ) | ( n9597 & ~n9602 ) ;
  assign n9604 = ( x106 & n9269 ) | ( x106 & ~n9347 ) | ( n9269 & ~n9347 ) ;
  assign n9605 = x106 & n9269 ;
  assign n9606 = ( ~n9274 & n9604 ) | ( ~n9274 & n9605 ) | ( n9604 & n9605 ) ;
  assign n9607 = ( n9274 & n9604 ) | ( n9274 & n9605 ) | ( n9604 & n9605 ) ;
  assign n9608 = ( n9274 & n9606 ) | ( n9274 & ~n9607 ) | ( n9606 & ~n9607 ) ;
  assign n9609 = ( x107 & n9603 ) | ( x107 & ~n9608 ) | ( n9603 & ~n9608 ) ;
  assign n9610 = ( x107 & n9275 ) | ( x107 & ~n9347 ) | ( n9275 & ~n9347 ) ;
  assign n9611 = x107 & n9275 ;
  assign n9612 = ( ~n9280 & n9610 ) | ( ~n9280 & n9611 ) | ( n9610 & n9611 ) ;
  assign n9613 = ( n9280 & n9610 ) | ( n9280 & n9611 ) | ( n9610 & n9611 ) ;
  assign n9614 = ( n9280 & n9612 ) | ( n9280 & ~n9613 ) | ( n9612 & ~n9613 ) ;
  assign n9615 = ( x108 & n9609 ) | ( x108 & ~n9614 ) | ( n9609 & ~n9614 ) ;
  assign n9616 = ( x108 & n9281 ) | ( x108 & ~n9347 ) | ( n9281 & ~n9347 ) ;
  assign n9617 = x108 & n9281 ;
  assign n9618 = ( ~n9286 & n9616 ) | ( ~n9286 & n9617 ) | ( n9616 & n9617 ) ;
  assign n9619 = ( n9286 & n9616 ) | ( n9286 & n9617 ) | ( n9616 & n9617 ) ;
  assign n9620 = ( n9286 & n9618 ) | ( n9286 & ~n9619 ) | ( n9618 & ~n9619 ) ;
  assign n9621 = ( x109 & n9615 ) | ( x109 & ~n9620 ) | ( n9615 & ~n9620 ) ;
  assign n9622 = ( x109 & n9287 ) | ( x109 & ~n9347 ) | ( n9287 & ~n9347 ) ;
  assign n9623 = x109 & n9287 ;
  assign n9624 = ( ~n9292 & n9622 ) | ( ~n9292 & n9623 ) | ( n9622 & n9623 ) ;
  assign n9625 = ( n9292 & n9622 ) | ( n9292 & n9623 ) | ( n9622 & n9623 ) ;
  assign n9626 = ( n9292 & n9624 ) | ( n9292 & ~n9625 ) | ( n9624 & ~n9625 ) ;
  assign n9627 = ( x110 & n9621 ) | ( x110 & ~n9626 ) | ( n9621 & ~n9626 ) ;
  assign n9628 = ( x110 & n9293 ) | ( x110 & ~n9347 ) | ( n9293 & ~n9347 ) ;
  assign n9629 = x110 & n9293 ;
  assign n9630 = ( ~n9298 & n9628 ) | ( ~n9298 & n9629 ) | ( n9628 & n9629 ) ;
  assign n9631 = ( n9298 & n9628 ) | ( n9298 & n9629 ) | ( n9628 & n9629 ) ;
  assign n9632 = ( n9298 & n9630 ) | ( n9298 & ~n9631 ) | ( n9630 & ~n9631 ) ;
  assign n9633 = ( x111 & n9627 ) | ( x111 & ~n9632 ) | ( n9627 & ~n9632 ) ;
  assign n9634 = ( x111 & n9299 ) | ( x111 & ~n9347 ) | ( n9299 & ~n9347 ) ;
  assign n9635 = x111 & n9299 ;
  assign n9636 = ( ~n9304 & n9634 ) | ( ~n9304 & n9635 ) | ( n9634 & n9635 ) ;
  assign n9637 = ( n9304 & n9634 ) | ( n9304 & n9635 ) | ( n9634 & n9635 ) ;
  assign n9638 = ( n9304 & n9636 ) | ( n9304 & ~n9637 ) | ( n9636 & ~n9637 ) ;
  assign n9639 = ( x112 & n9633 ) | ( x112 & ~n9638 ) | ( n9633 & ~n9638 ) ;
  assign n9640 = ( x112 & n9305 ) | ( x112 & ~n9347 ) | ( n9305 & ~n9347 ) ;
  assign n9641 = x112 & n9305 ;
  assign n9642 = ( ~n9310 & n9640 ) | ( ~n9310 & n9641 ) | ( n9640 & n9641 ) ;
  assign n9643 = ( n9310 & n9640 ) | ( n9310 & n9641 ) | ( n9640 & n9641 ) ;
  assign n9644 = ( n9310 & n9642 ) | ( n9310 & ~n9643 ) | ( n9642 & ~n9643 ) ;
  assign n9645 = ( x113 & n9639 ) | ( x113 & ~n9644 ) | ( n9639 & ~n9644 ) ;
  assign n9646 = ( x113 & n9311 ) | ( x113 & ~n9347 ) | ( n9311 & ~n9347 ) ;
  assign n9647 = x113 & n9311 ;
  assign n9648 = ( ~n9316 & n9646 ) | ( ~n9316 & n9647 ) | ( n9646 & n9647 ) ;
  assign n9649 = ( n9316 & n9646 ) | ( n9316 & n9647 ) | ( n9646 & n9647 ) ;
  assign n9650 = ( n9316 & n9648 ) | ( n9316 & ~n9649 ) | ( n9648 & ~n9649 ) ;
  assign n9651 = ( x114 & n9645 ) | ( x114 & ~n9650 ) | ( n9645 & ~n9650 ) ;
  assign n9652 = ( x114 & n9317 ) | ( x114 & ~n9347 ) | ( n9317 & ~n9347 ) ;
  assign n9653 = x114 & n9317 ;
  assign n9654 = ( ~n9322 & n9652 ) | ( ~n9322 & n9653 ) | ( n9652 & n9653 ) ;
  assign n9655 = ( n9322 & n9652 ) | ( n9322 & n9653 ) | ( n9652 & n9653 ) ;
  assign n9656 = ( n9322 & n9654 ) | ( n9322 & ~n9655 ) | ( n9654 & ~n9655 ) ;
  assign n9657 = ( x115 & n9651 ) | ( x115 & ~n9656 ) | ( n9651 & ~n9656 ) ;
  assign n9658 = ( x115 & n9323 ) | ( x115 & ~n9347 ) | ( n9323 & ~n9347 ) ;
  assign n9659 = x115 & n9323 ;
  assign n9660 = ( ~n9328 & n9658 ) | ( ~n9328 & n9659 ) | ( n9658 & n9659 ) ;
  assign n9661 = ( n9328 & n9658 ) | ( n9328 & n9659 ) | ( n9658 & n9659 ) ;
  assign n9662 = ( n9328 & n9660 ) | ( n9328 & ~n9661 ) | ( n9660 & ~n9661 ) ;
  assign n9663 = ( x116 & n9657 ) | ( x116 & ~n9662 ) | ( n9657 & ~n9662 ) ;
  assign n9664 = ( x116 & n9329 ) | ( x116 & ~n9347 ) | ( n9329 & ~n9347 ) ;
  assign n9665 = x116 & n9329 ;
  assign n9666 = ( ~n9334 & n9664 ) | ( ~n9334 & n9665 ) | ( n9664 & n9665 ) ;
  assign n9667 = ( n9334 & n9664 ) | ( n9334 & n9665 ) | ( n9664 & n9665 ) ;
  assign n9668 = ( n9334 & n9666 ) | ( n9334 & ~n9667 ) | ( n9666 & ~n9667 ) ;
  assign n9669 = ( x117 & n9663 ) | ( x117 & ~n9668 ) | ( n9663 & ~n9668 ) ;
  assign n9670 = ( x117 & n9335 ) | ( x117 & ~n9347 ) | ( n9335 & ~n9347 ) ;
  assign n9671 = x117 & n9335 ;
  assign n9672 = ( ~n9340 & n9670 ) | ( ~n9340 & n9671 ) | ( n9670 & n9671 ) ;
  assign n9673 = ( n9340 & n9670 ) | ( n9340 & n9671 ) | ( n9670 & n9671 ) ;
  assign n9674 = ( n9340 & n9672 ) | ( n9340 & ~n9673 ) | ( n9672 & ~n9673 ) ;
  assign n9675 = ( x118 & n9669 ) | ( x118 & ~n9674 ) | ( n9669 & ~n9674 ) ;
  assign n9676 = ( x119 & ~n9352 ) | ( x119 & n9675 ) | ( ~n9352 & n9675 ) ;
  assign n9677 = ( n137 & n138 ) | ( n137 & n9342 ) | ( n138 & n9342 ) ;
  assign n9678 = n9016 & n9677 ;
  assign n9679 = n389 | n9678 ;
  assign n9680 = ( x120 & n9676 ) | ( x120 & ~n9679 ) | ( n9676 & ~n9679 ) ;
  assign n9681 = n136 | n9680 ;
  assign n9682 = ( x119 & n9675 ) | ( x119 & n9681 ) | ( n9675 & n9681 ) ;
  assign n9683 = x119 | n9675 ;
  assign n9684 = ( ~n9352 & n9682 ) | ( ~n9352 & n9683 ) | ( n9682 & n9683 ) ;
  assign n9685 = ( n9352 & n9682 ) | ( n9352 & n9683 ) | ( n9682 & n9683 ) ;
  assign n9686 = ( n9352 & n9684 ) | ( n9352 & ~n9685 ) | ( n9684 & ~n9685 ) ;
  assign n9687 = ~x6 & x64 ;
  assign n9688 = ~x7 & n9681 ;
  assign n9689 = ( x7 & ~x64 ) | ( x7 & n9681 ) | ( ~x64 & n9681 ) ;
  assign n9690 = ( n9353 & ~n9688 ) | ( n9353 & n9689 ) | ( ~n9688 & n9689 ) ;
  assign n9691 = ( x65 & n9687 ) | ( x65 & ~n9690 ) | ( n9687 & ~n9690 ) ;
  assign n9692 = ( x65 & n9353 ) | ( x65 & n9681 ) | ( n9353 & n9681 ) ;
  assign n9693 = x65 | n9353 ;
  assign n9694 = ( ~n9356 & n9692 ) | ( ~n9356 & n9693 ) | ( n9692 & n9693 ) ;
  assign n9695 = ( n9356 & n9692 ) | ( n9356 & n9693 ) | ( n9692 & n9693 ) ;
  assign n9696 = ( n9356 & n9694 ) | ( n9356 & ~n9695 ) | ( n9694 & ~n9695 ) ;
  assign n9697 = ( x66 & n9691 ) | ( x66 & ~n9696 ) | ( n9691 & ~n9696 ) ;
  assign n9698 = ( x66 & n9357 ) | ( x66 & n9681 ) | ( n9357 & n9681 ) ;
  assign n9699 = x66 | n9357 ;
  assign n9700 = ( ~n9362 & n9698 ) | ( ~n9362 & n9699 ) | ( n9698 & n9699 ) ;
  assign n9701 = ( n9362 & n9698 ) | ( n9362 & n9699 ) | ( n9698 & n9699 ) ;
  assign n9702 = ( n9362 & n9700 ) | ( n9362 & ~n9701 ) | ( n9700 & ~n9701 ) ;
  assign n9703 = ( x67 & n9697 ) | ( x67 & ~n9702 ) | ( n9697 & ~n9702 ) ;
  assign n9704 = ( x67 & n9363 ) | ( x67 & ~n9681 ) | ( n9363 & ~n9681 ) ;
  assign n9705 = x67 & n9363 ;
  assign n9706 = ( ~n9368 & n9704 ) | ( ~n9368 & n9705 ) | ( n9704 & n9705 ) ;
  assign n9707 = ( n9368 & n9704 ) | ( n9368 & n9705 ) | ( n9704 & n9705 ) ;
  assign n9708 = ( n9368 & n9706 ) | ( n9368 & ~n9707 ) | ( n9706 & ~n9707 ) ;
  assign n9709 = ( x68 & n9703 ) | ( x68 & ~n9708 ) | ( n9703 & ~n9708 ) ;
  assign n9710 = ( x68 & n9369 ) | ( x68 & ~n9681 ) | ( n9369 & ~n9681 ) ;
  assign n9711 = x68 & n9369 ;
  assign n9712 = ( ~n9374 & n9710 ) | ( ~n9374 & n9711 ) | ( n9710 & n9711 ) ;
  assign n9713 = ( n9374 & n9710 ) | ( n9374 & n9711 ) | ( n9710 & n9711 ) ;
  assign n9714 = ( n9374 & n9712 ) | ( n9374 & ~n9713 ) | ( n9712 & ~n9713 ) ;
  assign n9715 = ( x69 & n9709 ) | ( x69 & ~n9714 ) | ( n9709 & ~n9714 ) ;
  assign n9716 = ( x69 & n9375 ) | ( x69 & ~n9681 ) | ( n9375 & ~n9681 ) ;
  assign n9717 = x69 & n9375 ;
  assign n9718 = ( ~n9380 & n9716 ) | ( ~n9380 & n9717 ) | ( n9716 & n9717 ) ;
  assign n9719 = ( n9380 & n9716 ) | ( n9380 & n9717 ) | ( n9716 & n9717 ) ;
  assign n9720 = ( n9380 & n9718 ) | ( n9380 & ~n9719 ) | ( n9718 & ~n9719 ) ;
  assign n9721 = ( x70 & n9715 ) | ( x70 & ~n9720 ) | ( n9715 & ~n9720 ) ;
  assign n9722 = ( x70 & n9381 ) | ( x70 & ~n9681 ) | ( n9381 & ~n9681 ) ;
  assign n9723 = x70 & n9381 ;
  assign n9724 = ( ~n9386 & n9722 ) | ( ~n9386 & n9723 ) | ( n9722 & n9723 ) ;
  assign n9725 = ( n9386 & n9722 ) | ( n9386 & n9723 ) | ( n9722 & n9723 ) ;
  assign n9726 = ( n9386 & n9724 ) | ( n9386 & ~n9725 ) | ( n9724 & ~n9725 ) ;
  assign n9727 = ( x71 & n9721 ) | ( x71 & ~n9726 ) | ( n9721 & ~n9726 ) ;
  assign n9728 = ( x71 & n9387 ) | ( x71 & ~n9681 ) | ( n9387 & ~n9681 ) ;
  assign n9729 = x71 & n9387 ;
  assign n9730 = ( ~n9392 & n9728 ) | ( ~n9392 & n9729 ) | ( n9728 & n9729 ) ;
  assign n9731 = ( n9392 & n9728 ) | ( n9392 & n9729 ) | ( n9728 & n9729 ) ;
  assign n9732 = ( n9392 & n9730 ) | ( n9392 & ~n9731 ) | ( n9730 & ~n9731 ) ;
  assign n9733 = ( x72 & n9727 ) | ( x72 & ~n9732 ) | ( n9727 & ~n9732 ) ;
  assign n9734 = ( x72 & n9393 ) | ( x72 & ~n9681 ) | ( n9393 & ~n9681 ) ;
  assign n9735 = x72 & n9393 ;
  assign n9736 = ( ~n9398 & n9734 ) | ( ~n9398 & n9735 ) | ( n9734 & n9735 ) ;
  assign n9737 = ( n9398 & n9734 ) | ( n9398 & n9735 ) | ( n9734 & n9735 ) ;
  assign n9738 = ( n9398 & n9736 ) | ( n9398 & ~n9737 ) | ( n9736 & ~n9737 ) ;
  assign n9739 = ( x73 & n9733 ) | ( x73 & ~n9738 ) | ( n9733 & ~n9738 ) ;
  assign n9740 = ( x73 & n9399 ) | ( x73 & ~n9681 ) | ( n9399 & ~n9681 ) ;
  assign n9741 = x73 & n9399 ;
  assign n9742 = ( ~n9404 & n9740 ) | ( ~n9404 & n9741 ) | ( n9740 & n9741 ) ;
  assign n9743 = ( n9404 & n9740 ) | ( n9404 & n9741 ) | ( n9740 & n9741 ) ;
  assign n9744 = ( n9404 & n9742 ) | ( n9404 & ~n9743 ) | ( n9742 & ~n9743 ) ;
  assign n9745 = ( x74 & n9739 ) | ( x74 & ~n9744 ) | ( n9739 & ~n9744 ) ;
  assign n9746 = ( x74 & n9405 ) | ( x74 & ~n9681 ) | ( n9405 & ~n9681 ) ;
  assign n9747 = x74 & n9405 ;
  assign n9748 = ( ~n9410 & n9746 ) | ( ~n9410 & n9747 ) | ( n9746 & n9747 ) ;
  assign n9749 = ( n9410 & n9746 ) | ( n9410 & n9747 ) | ( n9746 & n9747 ) ;
  assign n9750 = ( n9410 & n9748 ) | ( n9410 & ~n9749 ) | ( n9748 & ~n9749 ) ;
  assign n9751 = ( x75 & n9745 ) | ( x75 & ~n9750 ) | ( n9745 & ~n9750 ) ;
  assign n9752 = ( x75 & n9411 ) | ( x75 & ~n9681 ) | ( n9411 & ~n9681 ) ;
  assign n9753 = x75 & n9411 ;
  assign n9754 = ( ~n9416 & n9752 ) | ( ~n9416 & n9753 ) | ( n9752 & n9753 ) ;
  assign n9755 = ( n9416 & n9752 ) | ( n9416 & n9753 ) | ( n9752 & n9753 ) ;
  assign n9756 = ( n9416 & n9754 ) | ( n9416 & ~n9755 ) | ( n9754 & ~n9755 ) ;
  assign n9757 = ( x76 & n9751 ) | ( x76 & ~n9756 ) | ( n9751 & ~n9756 ) ;
  assign n9758 = ( x76 & n9417 ) | ( x76 & ~n9681 ) | ( n9417 & ~n9681 ) ;
  assign n9759 = x76 & n9417 ;
  assign n9760 = ( ~n9422 & n9758 ) | ( ~n9422 & n9759 ) | ( n9758 & n9759 ) ;
  assign n9761 = ( n9422 & n9758 ) | ( n9422 & n9759 ) | ( n9758 & n9759 ) ;
  assign n9762 = ( n9422 & n9760 ) | ( n9422 & ~n9761 ) | ( n9760 & ~n9761 ) ;
  assign n9763 = ( x77 & n9757 ) | ( x77 & ~n9762 ) | ( n9757 & ~n9762 ) ;
  assign n9764 = ( x77 & n9423 ) | ( x77 & ~n9681 ) | ( n9423 & ~n9681 ) ;
  assign n9765 = x77 & n9423 ;
  assign n9766 = ( ~n9428 & n9764 ) | ( ~n9428 & n9765 ) | ( n9764 & n9765 ) ;
  assign n9767 = ( n9428 & n9764 ) | ( n9428 & n9765 ) | ( n9764 & n9765 ) ;
  assign n9768 = ( n9428 & n9766 ) | ( n9428 & ~n9767 ) | ( n9766 & ~n9767 ) ;
  assign n9769 = ( x78 & n9763 ) | ( x78 & ~n9768 ) | ( n9763 & ~n9768 ) ;
  assign n9770 = ( x78 & n9429 ) | ( x78 & ~n9681 ) | ( n9429 & ~n9681 ) ;
  assign n9771 = x78 & n9429 ;
  assign n9772 = ( ~n9434 & n9770 ) | ( ~n9434 & n9771 ) | ( n9770 & n9771 ) ;
  assign n9773 = ( n9434 & n9770 ) | ( n9434 & n9771 ) | ( n9770 & n9771 ) ;
  assign n9774 = ( n9434 & n9772 ) | ( n9434 & ~n9773 ) | ( n9772 & ~n9773 ) ;
  assign n9775 = ( x79 & n9769 ) | ( x79 & ~n9774 ) | ( n9769 & ~n9774 ) ;
  assign n9776 = ( x79 & n9435 ) | ( x79 & ~n9681 ) | ( n9435 & ~n9681 ) ;
  assign n9777 = x79 & n9435 ;
  assign n9778 = ( ~n9440 & n9776 ) | ( ~n9440 & n9777 ) | ( n9776 & n9777 ) ;
  assign n9779 = ( n9440 & n9776 ) | ( n9440 & n9777 ) | ( n9776 & n9777 ) ;
  assign n9780 = ( n9440 & n9778 ) | ( n9440 & ~n9779 ) | ( n9778 & ~n9779 ) ;
  assign n9781 = ( x80 & n9775 ) | ( x80 & ~n9780 ) | ( n9775 & ~n9780 ) ;
  assign n9782 = ( x80 & n9441 ) | ( x80 & ~n9681 ) | ( n9441 & ~n9681 ) ;
  assign n9783 = x80 & n9441 ;
  assign n9784 = ( ~n9446 & n9782 ) | ( ~n9446 & n9783 ) | ( n9782 & n9783 ) ;
  assign n9785 = ( n9446 & n9782 ) | ( n9446 & n9783 ) | ( n9782 & n9783 ) ;
  assign n9786 = ( n9446 & n9784 ) | ( n9446 & ~n9785 ) | ( n9784 & ~n9785 ) ;
  assign n9787 = ( x81 & n9781 ) | ( x81 & ~n9786 ) | ( n9781 & ~n9786 ) ;
  assign n9788 = ( x81 & n9447 ) | ( x81 & ~n9681 ) | ( n9447 & ~n9681 ) ;
  assign n9789 = x81 & n9447 ;
  assign n9790 = ( ~n9452 & n9788 ) | ( ~n9452 & n9789 ) | ( n9788 & n9789 ) ;
  assign n9791 = ( n9452 & n9788 ) | ( n9452 & n9789 ) | ( n9788 & n9789 ) ;
  assign n9792 = ( n9452 & n9790 ) | ( n9452 & ~n9791 ) | ( n9790 & ~n9791 ) ;
  assign n9793 = ( x82 & n9787 ) | ( x82 & ~n9792 ) | ( n9787 & ~n9792 ) ;
  assign n9794 = ( x82 & n9453 ) | ( x82 & ~n9681 ) | ( n9453 & ~n9681 ) ;
  assign n9795 = x82 & n9453 ;
  assign n9796 = ( ~n9458 & n9794 ) | ( ~n9458 & n9795 ) | ( n9794 & n9795 ) ;
  assign n9797 = ( n9458 & n9794 ) | ( n9458 & n9795 ) | ( n9794 & n9795 ) ;
  assign n9798 = ( n9458 & n9796 ) | ( n9458 & ~n9797 ) | ( n9796 & ~n9797 ) ;
  assign n9799 = ( x83 & n9793 ) | ( x83 & ~n9798 ) | ( n9793 & ~n9798 ) ;
  assign n9800 = ( x83 & n9459 ) | ( x83 & ~n9681 ) | ( n9459 & ~n9681 ) ;
  assign n9801 = x83 & n9459 ;
  assign n9802 = ( ~n9464 & n9800 ) | ( ~n9464 & n9801 ) | ( n9800 & n9801 ) ;
  assign n9803 = ( n9464 & n9800 ) | ( n9464 & n9801 ) | ( n9800 & n9801 ) ;
  assign n9804 = ( n9464 & n9802 ) | ( n9464 & ~n9803 ) | ( n9802 & ~n9803 ) ;
  assign n9805 = ( x84 & n9799 ) | ( x84 & ~n9804 ) | ( n9799 & ~n9804 ) ;
  assign n9806 = ( x84 & n9465 ) | ( x84 & ~n9681 ) | ( n9465 & ~n9681 ) ;
  assign n9807 = x84 & n9465 ;
  assign n9808 = ( ~n9470 & n9806 ) | ( ~n9470 & n9807 ) | ( n9806 & n9807 ) ;
  assign n9809 = ( n9470 & n9806 ) | ( n9470 & n9807 ) | ( n9806 & n9807 ) ;
  assign n9810 = ( n9470 & n9808 ) | ( n9470 & ~n9809 ) | ( n9808 & ~n9809 ) ;
  assign n9811 = ( x85 & n9805 ) | ( x85 & ~n9810 ) | ( n9805 & ~n9810 ) ;
  assign n9812 = ( x85 & n9471 ) | ( x85 & ~n9681 ) | ( n9471 & ~n9681 ) ;
  assign n9813 = x85 & n9471 ;
  assign n9814 = ( ~n9476 & n9812 ) | ( ~n9476 & n9813 ) | ( n9812 & n9813 ) ;
  assign n9815 = ( n9476 & n9812 ) | ( n9476 & n9813 ) | ( n9812 & n9813 ) ;
  assign n9816 = ( n9476 & n9814 ) | ( n9476 & ~n9815 ) | ( n9814 & ~n9815 ) ;
  assign n9817 = ( x86 & n9811 ) | ( x86 & ~n9816 ) | ( n9811 & ~n9816 ) ;
  assign n9818 = ( x86 & n9477 ) | ( x86 & ~n9681 ) | ( n9477 & ~n9681 ) ;
  assign n9819 = x86 & n9477 ;
  assign n9820 = ( ~n9482 & n9818 ) | ( ~n9482 & n9819 ) | ( n9818 & n9819 ) ;
  assign n9821 = ( n9482 & n9818 ) | ( n9482 & n9819 ) | ( n9818 & n9819 ) ;
  assign n9822 = ( n9482 & n9820 ) | ( n9482 & ~n9821 ) | ( n9820 & ~n9821 ) ;
  assign n9823 = ( x87 & n9817 ) | ( x87 & ~n9822 ) | ( n9817 & ~n9822 ) ;
  assign n9824 = ( x87 & n9483 ) | ( x87 & ~n9681 ) | ( n9483 & ~n9681 ) ;
  assign n9825 = x87 & n9483 ;
  assign n9826 = ( ~n9488 & n9824 ) | ( ~n9488 & n9825 ) | ( n9824 & n9825 ) ;
  assign n9827 = ( n9488 & n9824 ) | ( n9488 & n9825 ) | ( n9824 & n9825 ) ;
  assign n9828 = ( n9488 & n9826 ) | ( n9488 & ~n9827 ) | ( n9826 & ~n9827 ) ;
  assign n9829 = ( x88 & n9823 ) | ( x88 & ~n9828 ) | ( n9823 & ~n9828 ) ;
  assign n9830 = ( x88 & n9489 ) | ( x88 & ~n9681 ) | ( n9489 & ~n9681 ) ;
  assign n9831 = x88 & n9489 ;
  assign n9832 = ( ~n9494 & n9830 ) | ( ~n9494 & n9831 ) | ( n9830 & n9831 ) ;
  assign n9833 = ( n9494 & n9830 ) | ( n9494 & n9831 ) | ( n9830 & n9831 ) ;
  assign n9834 = ( n9494 & n9832 ) | ( n9494 & ~n9833 ) | ( n9832 & ~n9833 ) ;
  assign n9835 = ( x89 & n9829 ) | ( x89 & ~n9834 ) | ( n9829 & ~n9834 ) ;
  assign n9836 = ( x89 & n9495 ) | ( x89 & ~n9681 ) | ( n9495 & ~n9681 ) ;
  assign n9837 = x89 & n9495 ;
  assign n9838 = ( ~n9500 & n9836 ) | ( ~n9500 & n9837 ) | ( n9836 & n9837 ) ;
  assign n9839 = ( n9500 & n9836 ) | ( n9500 & n9837 ) | ( n9836 & n9837 ) ;
  assign n9840 = ( n9500 & n9838 ) | ( n9500 & ~n9839 ) | ( n9838 & ~n9839 ) ;
  assign n9841 = ( x90 & n9835 ) | ( x90 & ~n9840 ) | ( n9835 & ~n9840 ) ;
  assign n9842 = ( x90 & n9501 ) | ( x90 & ~n9681 ) | ( n9501 & ~n9681 ) ;
  assign n9843 = x90 & n9501 ;
  assign n9844 = ( ~n9506 & n9842 ) | ( ~n9506 & n9843 ) | ( n9842 & n9843 ) ;
  assign n9845 = ( n9506 & n9842 ) | ( n9506 & n9843 ) | ( n9842 & n9843 ) ;
  assign n9846 = ( n9506 & n9844 ) | ( n9506 & ~n9845 ) | ( n9844 & ~n9845 ) ;
  assign n9847 = ( x91 & n9841 ) | ( x91 & ~n9846 ) | ( n9841 & ~n9846 ) ;
  assign n9848 = ( x91 & n9507 ) | ( x91 & ~n9681 ) | ( n9507 & ~n9681 ) ;
  assign n9849 = x91 & n9507 ;
  assign n9850 = ( ~n9512 & n9848 ) | ( ~n9512 & n9849 ) | ( n9848 & n9849 ) ;
  assign n9851 = ( n9512 & n9848 ) | ( n9512 & n9849 ) | ( n9848 & n9849 ) ;
  assign n9852 = ( n9512 & n9850 ) | ( n9512 & ~n9851 ) | ( n9850 & ~n9851 ) ;
  assign n9853 = ( x92 & n9847 ) | ( x92 & ~n9852 ) | ( n9847 & ~n9852 ) ;
  assign n9854 = ( x92 & n9513 ) | ( x92 & ~n9681 ) | ( n9513 & ~n9681 ) ;
  assign n9855 = x92 & n9513 ;
  assign n9856 = ( ~n9518 & n9854 ) | ( ~n9518 & n9855 ) | ( n9854 & n9855 ) ;
  assign n9857 = ( n9518 & n9854 ) | ( n9518 & n9855 ) | ( n9854 & n9855 ) ;
  assign n9858 = ( n9518 & n9856 ) | ( n9518 & ~n9857 ) | ( n9856 & ~n9857 ) ;
  assign n9859 = ( x93 & n9853 ) | ( x93 & ~n9858 ) | ( n9853 & ~n9858 ) ;
  assign n9860 = ( x93 & n9519 ) | ( x93 & ~n9681 ) | ( n9519 & ~n9681 ) ;
  assign n9861 = x93 & n9519 ;
  assign n9862 = ( ~n9524 & n9860 ) | ( ~n9524 & n9861 ) | ( n9860 & n9861 ) ;
  assign n9863 = ( n9524 & n9860 ) | ( n9524 & n9861 ) | ( n9860 & n9861 ) ;
  assign n9864 = ( n9524 & n9862 ) | ( n9524 & ~n9863 ) | ( n9862 & ~n9863 ) ;
  assign n9865 = ( x94 & n9859 ) | ( x94 & ~n9864 ) | ( n9859 & ~n9864 ) ;
  assign n9866 = ( x94 & n9525 ) | ( x94 & ~n9681 ) | ( n9525 & ~n9681 ) ;
  assign n9867 = x94 & n9525 ;
  assign n9868 = ( ~n9530 & n9866 ) | ( ~n9530 & n9867 ) | ( n9866 & n9867 ) ;
  assign n9869 = ( n9530 & n9866 ) | ( n9530 & n9867 ) | ( n9866 & n9867 ) ;
  assign n9870 = ( n9530 & n9868 ) | ( n9530 & ~n9869 ) | ( n9868 & ~n9869 ) ;
  assign n9871 = ( x95 & n9865 ) | ( x95 & ~n9870 ) | ( n9865 & ~n9870 ) ;
  assign n9872 = ( x95 & n9531 ) | ( x95 & ~n9681 ) | ( n9531 & ~n9681 ) ;
  assign n9873 = x95 & n9531 ;
  assign n9874 = ( ~n9536 & n9872 ) | ( ~n9536 & n9873 ) | ( n9872 & n9873 ) ;
  assign n9875 = ( n9536 & n9872 ) | ( n9536 & n9873 ) | ( n9872 & n9873 ) ;
  assign n9876 = ( n9536 & n9874 ) | ( n9536 & ~n9875 ) | ( n9874 & ~n9875 ) ;
  assign n9877 = ( x96 & n9871 ) | ( x96 & ~n9876 ) | ( n9871 & ~n9876 ) ;
  assign n9878 = ( x96 & n9537 ) | ( x96 & ~n9681 ) | ( n9537 & ~n9681 ) ;
  assign n9879 = x96 & n9537 ;
  assign n9880 = ( ~n9542 & n9878 ) | ( ~n9542 & n9879 ) | ( n9878 & n9879 ) ;
  assign n9881 = ( n9542 & n9878 ) | ( n9542 & n9879 ) | ( n9878 & n9879 ) ;
  assign n9882 = ( n9542 & n9880 ) | ( n9542 & ~n9881 ) | ( n9880 & ~n9881 ) ;
  assign n9883 = ( x97 & n9877 ) | ( x97 & ~n9882 ) | ( n9877 & ~n9882 ) ;
  assign n9884 = ( x97 & n9543 ) | ( x97 & ~n9681 ) | ( n9543 & ~n9681 ) ;
  assign n9885 = x97 & n9543 ;
  assign n9886 = ( ~n9548 & n9884 ) | ( ~n9548 & n9885 ) | ( n9884 & n9885 ) ;
  assign n9887 = ( n9548 & n9884 ) | ( n9548 & n9885 ) | ( n9884 & n9885 ) ;
  assign n9888 = ( n9548 & n9886 ) | ( n9548 & ~n9887 ) | ( n9886 & ~n9887 ) ;
  assign n9889 = ( x98 & n9883 ) | ( x98 & ~n9888 ) | ( n9883 & ~n9888 ) ;
  assign n9890 = ( x98 & n9549 ) | ( x98 & ~n9681 ) | ( n9549 & ~n9681 ) ;
  assign n9891 = x98 & n9549 ;
  assign n9892 = ( ~n9554 & n9890 ) | ( ~n9554 & n9891 ) | ( n9890 & n9891 ) ;
  assign n9893 = ( n9554 & n9890 ) | ( n9554 & n9891 ) | ( n9890 & n9891 ) ;
  assign n9894 = ( n9554 & n9892 ) | ( n9554 & ~n9893 ) | ( n9892 & ~n9893 ) ;
  assign n9895 = ( x99 & n9889 ) | ( x99 & ~n9894 ) | ( n9889 & ~n9894 ) ;
  assign n9896 = ( x99 & n9555 ) | ( x99 & ~n9681 ) | ( n9555 & ~n9681 ) ;
  assign n9897 = x99 & n9555 ;
  assign n9898 = ( ~n9560 & n9896 ) | ( ~n9560 & n9897 ) | ( n9896 & n9897 ) ;
  assign n9899 = ( n9560 & n9896 ) | ( n9560 & n9897 ) | ( n9896 & n9897 ) ;
  assign n9900 = ( n9560 & n9898 ) | ( n9560 & ~n9899 ) | ( n9898 & ~n9899 ) ;
  assign n9901 = ( x100 & n9895 ) | ( x100 & ~n9900 ) | ( n9895 & ~n9900 ) ;
  assign n9902 = ( x100 & n9561 ) | ( x100 & ~n9681 ) | ( n9561 & ~n9681 ) ;
  assign n9903 = x100 & n9561 ;
  assign n9904 = ( ~n9566 & n9902 ) | ( ~n9566 & n9903 ) | ( n9902 & n9903 ) ;
  assign n9905 = ( n9566 & n9902 ) | ( n9566 & n9903 ) | ( n9902 & n9903 ) ;
  assign n9906 = ( n9566 & n9904 ) | ( n9566 & ~n9905 ) | ( n9904 & ~n9905 ) ;
  assign n9907 = ( x101 & n9901 ) | ( x101 & ~n9906 ) | ( n9901 & ~n9906 ) ;
  assign n9908 = ( x101 & n9567 ) | ( x101 & ~n9681 ) | ( n9567 & ~n9681 ) ;
  assign n9909 = x101 & n9567 ;
  assign n9910 = ( ~n9572 & n9908 ) | ( ~n9572 & n9909 ) | ( n9908 & n9909 ) ;
  assign n9911 = ( n9572 & n9908 ) | ( n9572 & n9909 ) | ( n9908 & n9909 ) ;
  assign n9912 = ( n9572 & n9910 ) | ( n9572 & ~n9911 ) | ( n9910 & ~n9911 ) ;
  assign n9913 = ( x102 & n9907 ) | ( x102 & ~n9912 ) | ( n9907 & ~n9912 ) ;
  assign n9914 = ( x102 & n9573 ) | ( x102 & ~n9681 ) | ( n9573 & ~n9681 ) ;
  assign n9915 = x102 & n9573 ;
  assign n9916 = ( ~n9578 & n9914 ) | ( ~n9578 & n9915 ) | ( n9914 & n9915 ) ;
  assign n9917 = ( n9578 & n9914 ) | ( n9578 & n9915 ) | ( n9914 & n9915 ) ;
  assign n9918 = ( n9578 & n9916 ) | ( n9578 & ~n9917 ) | ( n9916 & ~n9917 ) ;
  assign n9919 = ( x103 & n9913 ) | ( x103 & ~n9918 ) | ( n9913 & ~n9918 ) ;
  assign n9920 = ( x103 & n9579 ) | ( x103 & ~n9681 ) | ( n9579 & ~n9681 ) ;
  assign n9921 = x103 & n9579 ;
  assign n9922 = ( ~n9584 & n9920 ) | ( ~n9584 & n9921 ) | ( n9920 & n9921 ) ;
  assign n9923 = ( n9584 & n9920 ) | ( n9584 & n9921 ) | ( n9920 & n9921 ) ;
  assign n9924 = ( n9584 & n9922 ) | ( n9584 & ~n9923 ) | ( n9922 & ~n9923 ) ;
  assign n9925 = ( x104 & n9919 ) | ( x104 & ~n9924 ) | ( n9919 & ~n9924 ) ;
  assign n9926 = ( x104 & n9585 ) | ( x104 & ~n9681 ) | ( n9585 & ~n9681 ) ;
  assign n9927 = x104 & n9585 ;
  assign n9928 = ( ~n9590 & n9926 ) | ( ~n9590 & n9927 ) | ( n9926 & n9927 ) ;
  assign n9929 = ( n9590 & n9926 ) | ( n9590 & n9927 ) | ( n9926 & n9927 ) ;
  assign n9930 = ( n9590 & n9928 ) | ( n9590 & ~n9929 ) | ( n9928 & ~n9929 ) ;
  assign n9931 = ( x105 & n9925 ) | ( x105 & ~n9930 ) | ( n9925 & ~n9930 ) ;
  assign n9932 = ( x105 & n9591 ) | ( x105 & ~n9681 ) | ( n9591 & ~n9681 ) ;
  assign n9933 = x105 & n9591 ;
  assign n9934 = ( ~n9596 & n9932 ) | ( ~n9596 & n9933 ) | ( n9932 & n9933 ) ;
  assign n9935 = ( n9596 & n9932 ) | ( n9596 & n9933 ) | ( n9932 & n9933 ) ;
  assign n9936 = ( n9596 & n9934 ) | ( n9596 & ~n9935 ) | ( n9934 & ~n9935 ) ;
  assign n9937 = ( x106 & n9931 ) | ( x106 & ~n9936 ) | ( n9931 & ~n9936 ) ;
  assign n9938 = ( x106 & n9597 ) | ( x106 & ~n9681 ) | ( n9597 & ~n9681 ) ;
  assign n9939 = x106 & n9597 ;
  assign n9940 = ( ~n9602 & n9938 ) | ( ~n9602 & n9939 ) | ( n9938 & n9939 ) ;
  assign n9941 = ( n9602 & n9938 ) | ( n9602 & n9939 ) | ( n9938 & n9939 ) ;
  assign n9942 = ( n9602 & n9940 ) | ( n9602 & ~n9941 ) | ( n9940 & ~n9941 ) ;
  assign n9943 = ( x107 & n9937 ) | ( x107 & ~n9942 ) | ( n9937 & ~n9942 ) ;
  assign n9944 = ( x107 & n9603 ) | ( x107 & ~n9681 ) | ( n9603 & ~n9681 ) ;
  assign n9945 = x107 & n9603 ;
  assign n9946 = ( ~n9608 & n9944 ) | ( ~n9608 & n9945 ) | ( n9944 & n9945 ) ;
  assign n9947 = ( n9608 & n9944 ) | ( n9608 & n9945 ) | ( n9944 & n9945 ) ;
  assign n9948 = ( n9608 & n9946 ) | ( n9608 & ~n9947 ) | ( n9946 & ~n9947 ) ;
  assign n9949 = ( x108 & n9943 ) | ( x108 & ~n9948 ) | ( n9943 & ~n9948 ) ;
  assign n9950 = ( x108 & n9609 ) | ( x108 & ~n9681 ) | ( n9609 & ~n9681 ) ;
  assign n9951 = x108 & n9609 ;
  assign n9952 = ( ~n9614 & n9950 ) | ( ~n9614 & n9951 ) | ( n9950 & n9951 ) ;
  assign n9953 = ( n9614 & n9950 ) | ( n9614 & n9951 ) | ( n9950 & n9951 ) ;
  assign n9954 = ( n9614 & n9952 ) | ( n9614 & ~n9953 ) | ( n9952 & ~n9953 ) ;
  assign n9955 = ( x109 & n9949 ) | ( x109 & ~n9954 ) | ( n9949 & ~n9954 ) ;
  assign n9956 = ( x109 & n9615 ) | ( x109 & ~n9681 ) | ( n9615 & ~n9681 ) ;
  assign n9957 = x109 & n9615 ;
  assign n9958 = ( ~n9620 & n9956 ) | ( ~n9620 & n9957 ) | ( n9956 & n9957 ) ;
  assign n9959 = ( n9620 & n9956 ) | ( n9620 & n9957 ) | ( n9956 & n9957 ) ;
  assign n9960 = ( n9620 & n9958 ) | ( n9620 & ~n9959 ) | ( n9958 & ~n9959 ) ;
  assign n9961 = ( x110 & n9955 ) | ( x110 & ~n9960 ) | ( n9955 & ~n9960 ) ;
  assign n9962 = ( x110 & n9621 ) | ( x110 & ~n9681 ) | ( n9621 & ~n9681 ) ;
  assign n9963 = x110 & n9621 ;
  assign n9964 = ( ~n9626 & n9962 ) | ( ~n9626 & n9963 ) | ( n9962 & n9963 ) ;
  assign n9965 = ( n9626 & n9962 ) | ( n9626 & n9963 ) | ( n9962 & n9963 ) ;
  assign n9966 = ( n9626 & n9964 ) | ( n9626 & ~n9965 ) | ( n9964 & ~n9965 ) ;
  assign n9967 = ( x111 & n9961 ) | ( x111 & ~n9966 ) | ( n9961 & ~n9966 ) ;
  assign n9968 = ( x111 & n9627 ) | ( x111 & ~n9681 ) | ( n9627 & ~n9681 ) ;
  assign n9969 = x111 & n9627 ;
  assign n9970 = ( ~n9632 & n9968 ) | ( ~n9632 & n9969 ) | ( n9968 & n9969 ) ;
  assign n9971 = ( n9632 & n9968 ) | ( n9632 & n9969 ) | ( n9968 & n9969 ) ;
  assign n9972 = ( n9632 & n9970 ) | ( n9632 & ~n9971 ) | ( n9970 & ~n9971 ) ;
  assign n9973 = ( x112 & n9967 ) | ( x112 & ~n9972 ) | ( n9967 & ~n9972 ) ;
  assign n9974 = ( x112 & n9633 ) | ( x112 & ~n9681 ) | ( n9633 & ~n9681 ) ;
  assign n9975 = x112 & n9633 ;
  assign n9976 = ( ~n9638 & n9974 ) | ( ~n9638 & n9975 ) | ( n9974 & n9975 ) ;
  assign n9977 = ( n9638 & n9974 ) | ( n9638 & n9975 ) | ( n9974 & n9975 ) ;
  assign n9978 = ( n9638 & n9976 ) | ( n9638 & ~n9977 ) | ( n9976 & ~n9977 ) ;
  assign n9979 = ( x113 & n9973 ) | ( x113 & ~n9978 ) | ( n9973 & ~n9978 ) ;
  assign n9980 = ( x113 & n9639 ) | ( x113 & ~n9681 ) | ( n9639 & ~n9681 ) ;
  assign n9981 = x113 & n9639 ;
  assign n9982 = ( ~n9644 & n9980 ) | ( ~n9644 & n9981 ) | ( n9980 & n9981 ) ;
  assign n9983 = ( n9644 & n9980 ) | ( n9644 & n9981 ) | ( n9980 & n9981 ) ;
  assign n9984 = ( n9644 & n9982 ) | ( n9644 & ~n9983 ) | ( n9982 & ~n9983 ) ;
  assign n9985 = ( x114 & n9979 ) | ( x114 & ~n9984 ) | ( n9979 & ~n9984 ) ;
  assign n9986 = ( x114 & n9645 ) | ( x114 & ~n9681 ) | ( n9645 & ~n9681 ) ;
  assign n9987 = x114 & n9645 ;
  assign n9988 = ( ~n9650 & n9986 ) | ( ~n9650 & n9987 ) | ( n9986 & n9987 ) ;
  assign n9989 = ( n9650 & n9986 ) | ( n9650 & n9987 ) | ( n9986 & n9987 ) ;
  assign n9990 = ( n9650 & n9988 ) | ( n9650 & ~n9989 ) | ( n9988 & ~n9989 ) ;
  assign n9991 = ( x115 & n9985 ) | ( x115 & ~n9990 ) | ( n9985 & ~n9990 ) ;
  assign n9992 = ( x115 & n9651 ) | ( x115 & ~n9681 ) | ( n9651 & ~n9681 ) ;
  assign n9993 = x115 & n9651 ;
  assign n9994 = ( ~n9656 & n9992 ) | ( ~n9656 & n9993 ) | ( n9992 & n9993 ) ;
  assign n9995 = ( n9656 & n9992 ) | ( n9656 & n9993 ) | ( n9992 & n9993 ) ;
  assign n9996 = ( n9656 & n9994 ) | ( n9656 & ~n9995 ) | ( n9994 & ~n9995 ) ;
  assign n9997 = ( x116 & n9991 ) | ( x116 & ~n9996 ) | ( n9991 & ~n9996 ) ;
  assign n9998 = ( x116 & n9657 ) | ( x116 & ~n9681 ) | ( n9657 & ~n9681 ) ;
  assign n9999 = x116 & n9657 ;
  assign n10000 = ( ~n9662 & n9998 ) | ( ~n9662 & n9999 ) | ( n9998 & n9999 ) ;
  assign n10001 = ( n9662 & n9998 ) | ( n9662 & n9999 ) | ( n9998 & n9999 ) ;
  assign n10002 = ( n9662 & n10000 ) | ( n9662 & ~n10001 ) | ( n10000 & ~n10001 ) ;
  assign n10003 = ( x117 & n9997 ) | ( x117 & ~n10002 ) | ( n9997 & ~n10002 ) ;
  assign n10004 = ( x117 & n9663 ) | ( x117 & ~n9681 ) | ( n9663 & ~n9681 ) ;
  assign n10005 = x117 & n9663 ;
  assign n10006 = ( ~n9668 & n10004 ) | ( ~n9668 & n10005 ) | ( n10004 & n10005 ) ;
  assign n10007 = ( n9668 & n10004 ) | ( n9668 & n10005 ) | ( n10004 & n10005 ) ;
  assign n10008 = ( n9668 & n10006 ) | ( n9668 & ~n10007 ) | ( n10006 & ~n10007 ) ;
  assign n10009 = ( x118 & n10003 ) | ( x118 & ~n10008 ) | ( n10003 & ~n10008 ) ;
  assign n10010 = ( x118 & n9669 ) | ( x118 & ~n9681 ) | ( n9669 & ~n9681 ) ;
  assign n10011 = x118 & n9669 ;
  assign n10012 = ( ~n9674 & n10010 ) | ( ~n9674 & n10011 ) | ( n10010 & n10011 ) ;
  assign n10013 = ( n9674 & n10010 ) | ( n9674 & n10011 ) | ( n10010 & n10011 ) ;
  assign n10014 = ( n9674 & n10012 ) | ( n9674 & ~n10013 ) | ( n10012 & ~n10013 ) ;
  assign n10015 = ( x119 & n10009 ) | ( x119 & ~n10014 ) | ( n10009 & ~n10014 ) ;
  assign n10016 = ( x120 & ~n9686 ) | ( x120 & n10015 ) | ( ~n9686 & n10015 ) ;
  assign n10017 = ( x120 & n136 ) | ( x120 & n9676 ) | ( n136 & n9676 ) ;
  assign n10018 = x120 | n9676 ;
  assign n10019 = ( n9679 & n10017 ) | ( n9679 & ~n10018 ) | ( n10017 & ~n10018 ) ;
  assign n10020 = ~n136 & n10019 ;
  assign n10021 = ~n134 & n9679 ;
  assign n10022 = ~x122 & n10021 ;
  assign n10023 = n136 & ~n10022 ;
  assign n10024 = ( n10016 & ~n10020 ) | ( n10016 & n10023 ) | ( ~n10020 & n10023 ) ;
  assign n10025 = ( x120 & n10015 ) | ( x120 & n10024 ) | ( n10015 & n10024 ) ;
  assign n10026 = x120 | n10015 ;
  assign n10027 = ( ~n9686 & n10025 ) | ( ~n9686 & n10026 ) | ( n10025 & n10026 ) ;
  assign n10028 = ( n9686 & n10025 ) | ( n9686 & n10026 ) | ( n10025 & n10026 ) ;
  assign n10029 = ( n9686 & n10027 ) | ( n9686 & ~n10028 ) | ( n10027 & ~n10028 ) ;
  assign n10030 = ~x5 & x64 ;
  assign n10031 = ~x6 & n10024 ;
  assign n10032 = ( x6 & ~x64 ) | ( x6 & n10024 ) | ( ~x64 & n10024 ) ;
  assign n10033 = ( n9687 & ~n10031 ) | ( n9687 & n10032 ) | ( ~n10031 & n10032 ) ;
  assign n10034 = ( x65 & n10030 ) | ( x65 & ~n10033 ) | ( n10030 & ~n10033 ) ;
  assign n10035 = ( x65 & n9687 ) | ( x65 & n10024 ) | ( n9687 & n10024 ) ;
  assign n10036 = x65 | n9687 ;
  assign n10037 = ( ~n9690 & n10035 ) | ( ~n9690 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10038 = ( n9690 & n10035 ) | ( n9690 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10039 = ( n9690 & n10037 ) | ( n9690 & ~n10038 ) | ( n10037 & ~n10038 ) ;
  assign n10040 = ( x66 & n10034 ) | ( x66 & ~n10039 ) | ( n10034 & ~n10039 ) ;
  assign n10041 = ( x66 & n9691 ) | ( x66 & n10024 ) | ( n9691 & n10024 ) ;
  assign n10042 = x66 | n9691 ;
  assign n10043 = ( ~n9696 & n10041 ) | ( ~n9696 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10044 = ( n9696 & n10041 ) | ( n9696 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10045 = ( n9696 & n10043 ) | ( n9696 & ~n10044 ) | ( n10043 & ~n10044 ) ;
  assign n10046 = ( x67 & n10040 ) | ( x67 & ~n10045 ) | ( n10040 & ~n10045 ) ;
  assign n10047 = ( x67 & n9697 ) | ( x67 & ~n10024 ) | ( n9697 & ~n10024 ) ;
  assign n10048 = x67 & n9697 ;
  assign n10049 = ( ~n9702 & n10047 ) | ( ~n9702 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10050 = ( n9702 & n10047 ) | ( n9702 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10051 = ( n9702 & n10049 ) | ( n9702 & ~n10050 ) | ( n10049 & ~n10050 ) ;
  assign n10052 = ( x68 & n10046 ) | ( x68 & ~n10051 ) | ( n10046 & ~n10051 ) ;
  assign n10053 = ( x68 & n9703 ) | ( x68 & ~n10024 ) | ( n9703 & ~n10024 ) ;
  assign n10054 = x68 & n9703 ;
  assign n10055 = ( ~n9708 & n10053 ) | ( ~n9708 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10056 = ( n9708 & n10053 ) | ( n9708 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10057 = ( n9708 & n10055 ) | ( n9708 & ~n10056 ) | ( n10055 & ~n10056 ) ;
  assign n10058 = ( x69 & n10052 ) | ( x69 & ~n10057 ) | ( n10052 & ~n10057 ) ;
  assign n10059 = ( x69 & n9709 ) | ( x69 & ~n10024 ) | ( n9709 & ~n10024 ) ;
  assign n10060 = x69 & n9709 ;
  assign n10061 = ( ~n9714 & n10059 ) | ( ~n9714 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10062 = ( n9714 & n10059 ) | ( n9714 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10063 = ( n9714 & n10061 ) | ( n9714 & ~n10062 ) | ( n10061 & ~n10062 ) ;
  assign n10064 = ( x70 & n10058 ) | ( x70 & ~n10063 ) | ( n10058 & ~n10063 ) ;
  assign n10065 = ( x70 & n9715 ) | ( x70 & ~n10024 ) | ( n9715 & ~n10024 ) ;
  assign n10066 = x70 & n9715 ;
  assign n10067 = ( ~n9720 & n10065 ) | ( ~n9720 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10068 = ( n9720 & n10065 ) | ( n9720 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10069 = ( n9720 & n10067 ) | ( n9720 & ~n10068 ) | ( n10067 & ~n10068 ) ;
  assign n10070 = ( x71 & n10064 ) | ( x71 & ~n10069 ) | ( n10064 & ~n10069 ) ;
  assign n10071 = ( x71 & n9721 ) | ( x71 & ~n10024 ) | ( n9721 & ~n10024 ) ;
  assign n10072 = x71 & n9721 ;
  assign n10073 = ( ~n9726 & n10071 ) | ( ~n9726 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10074 = ( n9726 & n10071 ) | ( n9726 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10075 = ( n9726 & n10073 ) | ( n9726 & ~n10074 ) | ( n10073 & ~n10074 ) ;
  assign n10076 = ( x72 & n10070 ) | ( x72 & ~n10075 ) | ( n10070 & ~n10075 ) ;
  assign n10077 = ( x72 & n9727 ) | ( x72 & ~n10024 ) | ( n9727 & ~n10024 ) ;
  assign n10078 = x72 & n9727 ;
  assign n10079 = ( ~n9732 & n10077 ) | ( ~n9732 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10080 = ( n9732 & n10077 ) | ( n9732 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10081 = ( n9732 & n10079 ) | ( n9732 & ~n10080 ) | ( n10079 & ~n10080 ) ;
  assign n10082 = ( x73 & n10076 ) | ( x73 & ~n10081 ) | ( n10076 & ~n10081 ) ;
  assign n10083 = ( x73 & n9733 ) | ( x73 & ~n10024 ) | ( n9733 & ~n10024 ) ;
  assign n10084 = x73 & n9733 ;
  assign n10085 = ( ~n9738 & n10083 ) | ( ~n9738 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10086 = ( n9738 & n10083 ) | ( n9738 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10087 = ( n9738 & n10085 ) | ( n9738 & ~n10086 ) | ( n10085 & ~n10086 ) ;
  assign n10088 = ( x74 & n10082 ) | ( x74 & ~n10087 ) | ( n10082 & ~n10087 ) ;
  assign n10089 = ( x74 & n9739 ) | ( x74 & ~n10024 ) | ( n9739 & ~n10024 ) ;
  assign n10090 = x74 & n9739 ;
  assign n10091 = ( ~n9744 & n10089 ) | ( ~n9744 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10092 = ( n9744 & n10089 ) | ( n9744 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10093 = ( n9744 & n10091 ) | ( n9744 & ~n10092 ) | ( n10091 & ~n10092 ) ;
  assign n10094 = ( x75 & n10088 ) | ( x75 & ~n10093 ) | ( n10088 & ~n10093 ) ;
  assign n10095 = ( x75 & n9745 ) | ( x75 & ~n10024 ) | ( n9745 & ~n10024 ) ;
  assign n10096 = x75 & n9745 ;
  assign n10097 = ( ~n9750 & n10095 ) | ( ~n9750 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10098 = ( n9750 & n10095 ) | ( n9750 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10099 = ( n9750 & n10097 ) | ( n9750 & ~n10098 ) | ( n10097 & ~n10098 ) ;
  assign n10100 = ( x76 & n10094 ) | ( x76 & ~n10099 ) | ( n10094 & ~n10099 ) ;
  assign n10101 = ( x76 & n9751 ) | ( x76 & ~n10024 ) | ( n9751 & ~n10024 ) ;
  assign n10102 = x76 & n9751 ;
  assign n10103 = ( ~n9756 & n10101 ) | ( ~n9756 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10104 = ( n9756 & n10101 ) | ( n9756 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10105 = ( n9756 & n10103 ) | ( n9756 & ~n10104 ) | ( n10103 & ~n10104 ) ;
  assign n10106 = ( x77 & n10100 ) | ( x77 & ~n10105 ) | ( n10100 & ~n10105 ) ;
  assign n10107 = ( x77 & n9757 ) | ( x77 & ~n10024 ) | ( n9757 & ~n10024 ) ;
  assign n10108 = x77 & n9757 ;
  assign n10109 = ( ~n9762 & n10107 ) | ( ~n9762 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10110 = ( n9762 & n10107 ) | ( n9762 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10111 = ( n9762 & n10109 ) | ( n9762 & ~n10110 ) | ( n10109 & ~n10110 ) ;
  assign n10112 = ( x78 & n10106 ) | ( x78 & ~n10111 ) | ( n10106 & ~n10111 ) ;
  assign n10113 = ( x78 & n9763 ) | ( x78 & ~n10024 ) | ( n9763 & ~n10024 ) ;
  assign n10114 = x78 & n9763 ;
  assign n10115 = ( ~n9768 & n10113 ) | ( ~n9768 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10116 = ( n9768 & n10113 ) | ( n9768 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10117 = ( n9768 & n10115 ) | ( n9768 & ~n10116 ) | ( n10115 & ~n10116 ) ;
  assign n10118 = ( x79 & n10112 ) | ( x79 & ~n10117 ) | ( n10112 & ~n10117 ) ;
  assign n10119 = ( x79 & n9769 ) | ( x79 & ~n10024 ) | ( n9769 & ~n10024 ) ;
  assign n10120 = x79 & n9769 ;
  assign n10121 = ( ~n9774 & n10119 ) | ( ~n9774 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10122 = ( n9774 & n10119 ) | ( n9774 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10123 = ( n9774 & n10121 ) | ( n9774 & ~n10122 ) | ( n10121 & ~n10122 ) ;
  assign n10124 = ( x80 & n10118 ) | ( x80 & ~n10123 ) | ( n10118 & ~n10123 ) ;
  assign n10125 = ( x80 & n9775 ) | ( x80 & ~n10024 ) | ( n9775 & ~n10024 ) ;
  assign n10126 = x80 & n9775 ;
  assign n10127 = ( ~n9780 & n10125 ) | ( ~n9780 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10128 = ( n9780 & n10125 ) | ( n9780 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10129 = ( n9780 & n10127 ) | ( n9780 & ~n10128 ) | ( n10127 & ~n10128 ) ;
  assign n10130 = ( x81 & n10124 ) | ( x81 & ~n10129 ) | ( n10124 & ~n10129 ) ;
  assign n10131 = ( x81 & n9781 ) | ( x81 & ~n10024 ) | ( n9781 & ~n10024 ) ;
  assign n10132 = x81 & n9781 ;
  assign n10133 = ( ~n9786 & n10131 ) | ( ~n9786 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10134 = ( n9786 & n10131 ) | ( n9786 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10135 = ( n9786 & n10133 ) | ( n9786 & ~n10134 ) | ( n10133 & ~n10134 ) ;
  assign n10136 = ( x82 & n10130 ) | ( x82 & ~n10135 ) | ( n10130 & ~n10135 ) ;
  assign n10137 = ( x82 & n9787 ) | ( x82 & ~n10024 ) | ( n9787 & ~n10024 ) ;
  assign n10138 = x82 & n9787 ;
  assign n10139 = ( ~n9792 & n10137 ) | ( ~n9792 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10140 = ( n9792 & n10137 ) | ( n9792 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10141 = ( n9792 & n10139 ) | ( n9792 & ~n10140 ) | ( n10139 & ~n10140 ) ;
  assign n10142 = ( x83 & n10136 ) | ( x83 & ~n10141 ) | ( n10136 & ~n10141 ) ;
  assign n10143 = ( x83 & n9793 ) | ( x83 & ~n10024 ) | ( n9793 & ~n10024 ) ;
  assign n10144 = x83 & n9793 ;
  assign n10145 = ( ~n9798 & n10143 ) | ( ~n9798 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10146 = ( n9798 & n10143 ) | ( n9798 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10147 = ( n9798 & n10145 ) | ( n9798 & ~n10146 ) | ( n10145 & ~n10146 ) ;
  assign n10148 = ( x84 & n10142 ) | ( x84 & ~n10147 ) | ( n10142 & ~n10147 ) ;
  assign n10149 = ( x84 & n9799 ) | ( x84 & ~n10024 ) | ( n9799 & ~n10024 ) ;
  assign n10150 = x84 & n9799 ;
  assign n10151 = ( ~n9804 & n10149 ) | ( ~n9804 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = ( n9804 & n10149 ) | ( n9804 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10153 = ( n9804 & n10151 ) | ( n9804 & ~n10152 ) | ( n10151 & ~n10152 ) ;
  assign n10154 = ( x85 & n10148 ) | ( x85 & ~n10153 ) | ( n10148 & ~n10153 ) ;
  assign n10155 = ( x85 & n9805 ) | ( x85 & ~n10024 ) | ( n9805 & ~n10024 ) ;
  assign n10156 = x85 & n9805 ;
  assign n10157 = ( ~n9810 & n10155 ) | ( ~n9810 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = ( n9810 & n10155 ) | ( n9810 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10159 = ( n9810 & n10157 ) | ( n9810 & ~n10158 ) | ( n10157 & ~n10158 ) ;
  assign n10160 = ( x86 & n10154 ) | ( x86 & ~n10159 ) | ( n10154 & ~n10159 ) ;
  assign n10161 = ( x86 & n9811 ) | ( x86 & ~n10024 ) | ( n9811 & ~n10024 ) ;
  assign n10162 = x86 & n9811 ;
  assign n10163 = ( ~n9816 & n10161 ) | ( ~n9816 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10164 = ( n9816 & n10161 ) | ( n9816 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10165 = ( n9816 & n10163 ) | ( n9816 & ~n10164 ) | ( n10163 & ~n10164 ) ;
  assign n10166 = ( x87 & n10160 ) | ( x87 & ~n10165 ) | ( n10160 & ~n10165 ) ;
  assign n10167 = ( x87 & n9817 ) | ( x87 & ~n10024 ) | ( n9817 & ~n10024 ) ;
  assign n10168 = x87 & n9817 ;
  assign n10169 = ( ~n9822 & n10167 ) | ( ~n9822 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10170 = ( n9822 & n10167 ) | ( n9822 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10171 = ( n9822 & n10169 ) | ( n9822 & ~n10170 ) | ( n10169 & ~n10170 ) ;
  assign n10172 = ( x88 & n10166 ) | ( x88 & ~n10171 ) | ( n10166 & ~n10171 ) ;
  assign n10173 = ( x88 & n9823 ) | ( x88 & ~n10024 ) | ( n9823 & ~n10024 ) ;
  assign n10174 = x88 & n9823 ;
  assign n10175 = ( ~n9828 & n10173 ) | ( ~n9828 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10176 = ( n9828 & n10173 ) | ( n9828 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10177 = ( n9828 & n10175 ) | ( n9828 & ~n10176 ) | ( n10175 & ~n10176 ) ;
  assign n10178 = ( x89 & n10172 ) | ( x89 & ~n10177 ) | ( n10172 & ~n10177 ) ;
  assign n10179 = ( x89 & n9829 ) | ( x89 & ~n10024 ) | ( n9829 & ~n10024 ) ;
  assign n10180 = x89 & n9829 ;
  assign n10181 = ( ~n9834 & n10179 ) | ( ~n9834 & n10180 ) | ( n10179 & n10180 ) ;
  assign n10182 = ( n9834 & n10179 ) | ( n9834 & n10180 ) | ( n10179 & n10180 ) ;
  assign n10183 = ( n9834 & n10181 ) | ( n9834 & ~n10182 ) | ( n10181 & ~n10182 ) ;
  assign n10184 = ( x90 & n10178 ) | ( x90 & ~n10183 ) | ( n10178 & ~n10183 ) ;
  assign n10185 = ( x90 & n9835 ) | ( x90 & ~n10024 ) | ( n9835 & ~n10024 ) ;
  assign n10186 = x90 & n9835 ;
  assign n10187 = ( ~n9840 & n10185 ) | ( ~n9840 & n10186 ) | ( n10185 & n10186 ) ;
  assign n10188 = ( n9840 & n10185 ) | ( n9840 & n10186 ) | ( n10185 & n10186 ) ;
  assign n10189 = ( n9840 & n10187 ) | ( n9840 & ~n10188 ) | ( n10187 & ~n10188 ) ;
  assign n10190 = ( x91 & n10184 ) | ( x91 & ~n10189 ) | ( n10184 & ~n10189 ) ;
  assign n10191 = ( x91 & n9841 ) | ( x91 & ~n10024 ) | ( n9841 & ~n10024 ) ;
  assign n10192 = x91 & n9841 ;
  assign n10193 = ( ~n9846 & n10191 ) | ( ~n9846 & n10192 ) | ( n10191 & n10192 ) ;
  assign n10194 = ( n9846 & n10191 ) | ( n9846 & n10192 ) | ( n10191 & n10192 ) ;
  assign n10195 = ( n9846 & n10193 ) | ( n9846 & ~n10194 ) | ( n10193 & ~n10194 ) ;
  assign n10196 = ( x92 & n10190 ) | ( x92 & ~n10195 ) | ( n10190 & ~n10195 ) ;
  assign n10197 = ( x92 & n9847 ) | ( x92 & ~n10024 ) | ( n9847 & ~n10024 ) ;
  assign n10198 = x92 & n9847 ;
  assign n10199 = ( ~n9852 & n10197 ) | ( ~n9852 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10200 = ( n9852 & n10197 ) | ( n9852 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10201 = ( n9852 & n10199 ) | ( n9852 & ~n10200 ) | ( n10199 & ~n10200 ) ;
  assign n10202 = ( x93 & n10196 ) | ( x93 & ~n10201 ) | ( n10196 & ~n10201 ) ;
  assign n10203 = ( x93 & n9853 ) | ( x93 & ~n10024 ) | ( n9853 & ~n10024 ) ;
  assign n10204 = x93 & n9853 ;
  assign n10205 = ( ~n9858 & n10203 ) | ( ~n9858 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10206 = ( n9858 & n10203 ) | ( n9858 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10207 = ( n9858 & n10205 ) | ( n9858 & ~n10206 ) | ( n10205 & ~n10206 ) ;
  assign n10208 = ( x94 & n10202 ) | ( x94 & ~n10207 ) | ( n10202 & ~n10207 ) ;
  assign n10209 = ( x94 & n9859 ) | ( x94 & ~n10024 ) | ( n9859 & ~n10024 ) ;
  assign n10210 = x94 & n9859 ;
  assign n10211 = ( ~n9864 & n10209 ) | ( ~n9864 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10212 = ( n9864 & n10209 ) | ( n9864 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10213 = ( n9864 & n10211 ) | ( n9864 & ~n10212 ) | ( n10211 & ~n10212 ) ;
  assign n10214 = ( x95 & n10208 ) | ( x95 & ~n10213 ) | ( n10208 & ~n10213 ) ;
  assign n10215 = ( x95 & n9865 ) | ( x95 & ~n10024 ) | ( n9865 & ~n10024 ) ;
  assign n10216 = x95 & n9865 ;
  assign n10217 = ( ~n9870 & n10215 ) | ( ~n9870 & n10216 ) | ( n10215 & n10216 ) ;
  assign n10218 = ( n9870 & n10215 ) | ( n9870 & n10216 ) | ( n10215 & n10216 ) ;
  assign n10219 = ( n9870 & n10217 ) | ( n9870 & ~n10218 ) | ( n10217 & ~n10218 ) ;
  assign n10220 = ( x96 & n10214 ) | ( x96 & ~n10219 ) | ( n10214 & ~n10219 ) ;
  assign n10221 = ( x96 & n9871 ) | ( x96 & ~n10024 ) | ( n9871 & ~n10024 ) ;
  assign n10222 = x96 & n9871 ;
  assign n10223 = ( ~n9876 & n10221 ) | ( ~n9876 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10224 = ( n9876 & n10221 ) | ( n9876 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10225 = ( n9876 & n10223 ) | ( n9876 & ~n10224 ) | ( n10223 & ~n10224 ) ;
  assign n10226 = ( x97 & n10220 ) | ( x97 & ~n10225 ) | ( n10220 & ~n10225 ) ;
  assign n10227 = ( x97 & n9877 ) | ( x97 & ~n10024 ) | ( n9877 & ~n10024 ) ;
  assign n10228 = x97 & n9877 ;
  assign n10229 = ( ~n9882 & n10227 ) | ( ~n9882 & n10228 ) | ( n10227 & n10228 ) ;
  assign n10230 = ( n9882 & n10227 ) | ( n9882 & n10228 ) | ( n10227 & n10228 ) ;
  assign n10231 = ( n9882 & n10229 ) | ( n9882 & ~n10230 ) | ( n10229 & ~n10230 ) ;
  assign n10232 = ( x98 & n10226 ) | ( x98 & ~n10231 ) | ( n10226 & ~n10231 ) ;
  assign n10233 = ( x98 & n9883 ) | ( x98 & ~n10024 ) | ( n9883 & ~n10024 ) ;
  assign n10234 = x98 & n9883 ;
  assign n10235 = ( ~n9888 & n10233 ) | ( ~n9888 & n10234 ) | ( n10233 & n10234 ) ;
  assign n10236 = ( n9888 & n10233 ) | ( n9888 & n10234 ) | ( n10233 & n10234 ) ;
  assign n10237 = ( n9888 & n10235 ) | ( n9888 & ~n10236 ) | ( n10235 & ~n10236 ) ;
  assign n10238 = ( x99 & n10232 ) | ( x99 & ~n10237 ) | ( n10232 & ~n10237 ) ;
  assign n10239 = ( x99 & n9889 ) | ( x99 & ~n10024 ) | ( n9889 & ~n10024 ) ;
  assign n10240 = x99 & n9889 ;
  assign n10241 = ( ~n9894 & n10239 ) | ( ~n9894 & n10240 ) | ( n10239 & n10240 ) ;
  assign n10242 = ( n9894 & n10239 ) | ( n9894 & n10240 ) | ( n10239 & n10240 ) ;
  assign n10243 = ( n9894 & n10241 ) | ( n9894 & ~n10242 ) | ( n10241 & ~n10242 ) ;
  assign n10244 = ( x100 & n10238 ) | ( x100 & ~n10243 ) | ( n10238 & ~n10243 ) ;
  assign n10245 = ( x100 & n9895 ) | ( x100 & ~n10024 ) | ( n9895 & ~n10024 ) ;
  assign n10246 = x100 & n9895 ;
  assign n10247 = ( ~n9900 & n10245 ) | ( ~n9900 & n10246 ) | ( n10245 & n10246 ) ;
  assign n10248 = ( n9900 & n10245 ) | ( n9900 & n10246 ) | ( n10245 & n10246 ) ;
  assign n10249 = ( n9900 & n10247 ) | ( n9900 & ~n10248 ) | ( n10247 & ~n10248 ) ;
  assign n10250 = ( x101 & n10244 ) | ( x101 & ~n10249 ) | ( n10244 & ~n10249 ) ;
  assign n10251 = ( x101 & n9901 ) | ( x101 & ~n10024 ) | ( n9901 & ~n10024 ) ;
  assign n10252 = x101 & n9901 ;
  assign n10253 = ( ~n9906 & n10251 ) | ( ~n9906 & n10252 ) | ( n10251 & n10252 ) ;
  assign n10254 = ( n9906 & n10251 ) | ( n9906 & n10252 ) | ( n10251 & n10252 ) ;
  assign n10255 = ( n9906 & n10253 ) | ( n9906 & ~n10254 ) | ( n10253 & ~n10254 ) ;
  assign n10256 = ( x102 & n10250 ) | ( x102 & ~n10255 ) | ( n10250 & ~n10255 ) ;
  assign n10257 = ( x102 & n9907 ) | ( x102 & ~n10024 ) | ( n9907 & ~n10024 ) ;
  assign n10258 = x102 & n9907 ;
  assign n10259 = ( ~n9912 & n10257 ) | ( ~n9912 & n10258 ) | ( n10257 & n10258 ) ;
  assign n10260 = ( n9912 & n10257 ) | ( n9912 & n10258 ) | ( n10257 & n10258 ) ;
  assign n10261 = ( n9912 & n10259 ) | ( n9912 & ~n10260 ) | ( n10259 & ~n10260 ) ;
  assign n10262 = ( x103 & n10256 ) | ( x103 & ~n10261 ) | ( n10256 & ~n10261 ) ;
  assign n10263 = ( x103 & n9913 ) | ( x103 & ~n10024 ) | ( n9913 & ~n10024 ) ;
  assign n10264 = x103 & n9913 ;
  assign n10265 = ( ~n9918 & n10263 ) | ( ~n9918 & n10264 ) | ( n10263 & n10264 ) ;
  assign n10266 = ( n9918 & n10263 ) | ( n9918 & n10264 ) | ( n10263 & n10264 ) ;
  assign n10267 = ( n9918 & n10265 ) | ( n9918 & ~n10266 ) | ( n10265 & ~n10266 ) ;
  assign n10268 = ( x104 & n10262 ) | ( x104 & ~n10267 ) | ( n10262 & ~n10267 ) ;
  assign n10269 = ( x104 & n9919 ) | ( x104 & ~n10024 ) | ( n9919 & ~n10024 ) ;
  assign n10270 = x104 & n9919 ;
  assign n10271 = ( ~n9924 & n10269 ) | ( ~n9924 & n10270 ) | ( n10269 & n10270 ) ;
  assign n10272 = ( n9924 & n10269 ) | ( n9924 & n10270 ) | ( n10269 & n10270 ) ;
  assign n10273 = ( n9924 & n10271 ) | ( n9924 & ~n10272 ) | ( n10271 & ~n10272 ) ;
  assign n10274 = ( x105 & n10268 ) | ( x105 & ~n10273 ) | ( n10268 & ~n10273 ) ;
  assign n10275 = ( x105 & n9925 ) | ( x105 & ~n10024 ) | ( n9925 & ~n10024 ) ;
  assign n10276 = x105 & n9925 ;
  assign n10277 = ( ~n9930 & n10275 ) | ( ~n9930 & n10276 ) | ( n10275 & n10276 ) ;
  assign n10278 = ( n9930 & n10275 ) | ( n9930 & n10276 ) | ( n10275 & n10276 ) ;
  assign n10279 = ( n9930 & n10277 ) | ( n9930 & ~n10278 ) | ( n10277 & ~n10278 ) ;
  assign n10280 = ( x106 & n10274 ) | ( x106 & ~n10279 ) | ( n10274 & ~n10279 ) ;
  assign n10281 = ( x106 & n9931 ) | ( x106 & ~n10024 ) | ( n9931 & ~n10024 ) ;
  assign n10282 = x106 & n9931 ;
  assign n10283 = ( ~n9936 & n10281 ) | ( ~n9936 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10284 = ( n9936 & n10281 ) | ( n9936 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10285 = ( n9936 & n10283 ) | ( n9936 & ~n10284 ) | ( n10283 & ~n10284 ) ;
  assign n10286 = ( x107 & n10280 ) | ( x107 & ~n10285 ) | ( n10280 & ~n10285 ) ;
  assign n10287 = ( x107 & n9937 ) | ( x107 & ~n10024 ) | ( n9937 & ~n10024 ) ;
  assign n10288 = x107 & n9937 ;
  assign n10289 = ( ~n9942 & n10287 ) | ( ~n9942 & n10288 ) | ( n10287 & n10288 ) ;
  assign n10290 = ( n9942 & n10287 ) | ( n9942 & n10288 ) | ( n10287 & n10288 ) ;
  assign n10291 = ( n9942 & n10289 ) | ( n9942 & ~n10290 ) | ( n10289 & ~n10290 ) ;
  assign n10292 = ( x108 & n10286 ) | ( x108 & ~n10291 ) | ( n10286 & ~n10291 ) ;
  assign n10293 = ( x108 & n9943 ) | ( x108 & ~n10024 ) | ( n9943 & ~n10024 ) ;
  assign n10294 = x108 & n9943 ;
  assign n10295 = ( ~n9948 & n10293 ) | ( ~n9948 & n10294 ) | ( n10293 & n10294 ) ;
  assign n10296 = ( n9948 & n10293 ) | ( n9948 & n10294 ) | ( n10293 & n10294 ) ;
  assign n10297 = ( n9948 & n10295 ) | ( n9948 & ~n10296 ) | ( n10295 & ~n10296 ) ;
  assign n10298 = ( x109 & n10292 ) | ( x109 & ~n10297 ) | ( n10292 & ~n10297 ) ;
  assign n10299 = ( x109 & n9949 ) | ( x109 & ~n10024 ) | ( n9949 & ~n10024 ) ;
  assign n10300 = x109 & n9949 ;
  assign n10301 = ( ~n9954 & n10299 ) | ( ~n9954 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10302 = ( n9954 & n10299 ) | ( n9954 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10303 = ( n9954 & n10301 ) | ( n9954 & ~n10302 ) | ( n10301 & ~n10302 ) ;
  assign n10304 = ( x110 & n10298 ) | ( x110 & ~n10303 ) | ( n10298 & ~n10303 ) ;
  assign n10305 = ( x110 & n9955 ) | ( x110 & ~n10024 ) | ( n9955 & ~n10024 ) ;
  assign n10306 = x110 & n9955 ;
  assign n10307 = ( ~n9960 & n10305 ) | ( ~n9960 & n10306 ) | ( n10305 & n10306 ) ;
  assign n10308 = ( n9960 & n10305 ) | ( n9960 & n10306 ) | ( n10305 & n10306 ) ;
  assign n10309 = ( n9960 & n10307 ) | ( n9960 & ~n10308 ) | ( n10307 & ~n10308 ) ;
  assign n10310 = ( x111 & n10304 ) | ( x111 & ~n10309 ) | ( n10304 & ~n10309 ) ;
  assign n10311 = ( x111 & n9961 ) | ( x111 & ~n10024 ) | ( n9961 & ~n10024 ) ;
  assign n10312 = x111 & n9961 ;
  assign n10313 = ( ~n9966 & n10311 ) | ( ~n9966 & n10312 ) | ( n10311 & n10312 ) ;
  assign n10314 = ( n9966 & n10311 ) | ( n9966 & n10312 ) | ( n10311 & n10312 ) ;
  assign n10315 = ( n9966 & n10313 ) | ( n9966 & ~n10314 ) | ( n10313 & ~n10314 ) ;
  assign n10316 = ( x112 & n10310 ) | ( x112 & ~n10315 ) | ( n10310 & ~n10315 ) ;
  assign n10317 = ( x112 & n9967 ) | ( x112 & ~n10024 ) | ( n9967 & ~n10024 ) ;
  assign n10318 = x112 & n9967 ;
  assign n10319 = ( ~n9972 & n10317 ) | ( ~n9972 & n10318 ) | ( n10317 & n10318 ) ;
  assign n10320 = ( n9972 & n10317 ) | ( n9972 & n10318 ) | ( n10317 & n10318 ) ;
  assign n10321 = ( n9972 & n10319 ) | ( n9972 & ~n10320 ) | ( n10319 & ~n10320 ) ;
  assign n10322 = ( x113 & n10316 ) | ( x113 & ~n10321 ) | ( n10316 & ~n10321 ) ;
  assign n10323 = ( x113 & n9973 ) | ( x113 & ~n10024 ) | ( n9973 & ~n10024 ) ;
  assign n10324 = x113 & n9973 ;
  assign n10325 = ( ~n9978 & n10323 ) | ( ~n9978 & n10324 ) | ( n10323 & n10324 ) ;
  assign n10326 = ( n9978 & n10323 ) | ( n9978 & n10324 ) | ( n10323 & n10324 ) ;
  assign n10327 = ( n9978 & n10325 ) | ( n9978 & ~n10326 ) | ( n10325 & ~n10326 ) ;
  assign n10328 = ( x114 & n10322 ) | ( x114 & ~n10327 ) | ( n10322 & ~n10327 ) ;
  assign n10329 = ( x114 & n9979 ) | ( x114 & ~n10024 ) | ( n9979 & ~n10024 ) ;
  assign n10330 = x114 & n9979 ;
  assign n10331 = ( ~n9984 & n10329 ) | ( ~n9984 & n10330 ) | ( n10329 & n10330 ) ;
  assign n10332 = ( n9984 & n10329 ) | ( n9984 & n10330 ) | ( n10329 & n10330 ) ;
  assign n10333 = ( n9984 & n10331 ) | ( n9984 & ~n10332 ) | ( n10331 & ~n10332 ) ;
  assign n10334 = ( x115 & n10328 ) | ( x115 & ~n10333 ) | ( n10328 & ~n10333 ) ;
  assign n10335 = ( x115 & n9985 ) | ( x115 & ~n10024 ) | ( n9985 & ~n10024 ) ;
  assign n10336 = x115 & n9985 ;
  assign n10337 = ( ~n9990 & n10335 ) | ( ~n9990 & n10336 ) | ( n10335 & n10336 ) ;
  assign n10338 = ( n9990 & n10335 ) | ( n9990 & n10336 ) | ( n10335 & n10336 ) ;
  assign n10339 = ( n9990 & n10337 ) | ( n9990 & ~n10338 ) | ( n10337 & ~n10338 ) ;
  assign n10340 = ( x116 & n10334 ) | ( x116 & ~n10339 ) | ( n10334 & ~n10339 ) ;
  assign n10341 = ( x116 & n9991 ) | ( x116 & ~n10024 ) | ( n9991 & ~n10024 ) ;
  assign n10342 = x116 & n9991 ;
  assign n10343 = ( ~n9996 & n10341 ) | ( ~n9996 & n10342 ) | ( n10341 & n10342 ) ;
  assign n10344 = ( n9996 & n10341 ) | ( n9996 & n10342 ) | ( n10341 & n10342 ) ;
  assign n10345 = ( n9996 & n10343 ) | ( n9996 & ~n10344 ) | ( n10343 & ~n10344 ) ;
  assign n10346 = ( x117 & n10340 ) | ( x117 & ~n10345 ) | ( n10340 & ~n10345 ) ;
  assign n10347 = ( x117 & n9997 ) | ( x117 & ~n10024 ) | ( n9997 & ~n10024 ) ;
  assign n10348 = x117 & n9997 ;
  assign n10349 = ( ~n10002 & n10347 ) | ( ~n10002 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10350 = ( n10002 & n10347 ) | ( n10002 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10351 = ( n10002 & n10349 ) | ( n10002 & ~n10350 ) | ( n10349 & ~n10350 ) ;
  assign n10352 = ( x118 & n10346 ) | ( x118 & ~n10351 ) | ( n10346 & ~n10351 ) ;
  assign n10353 = ( x118 & n10003 ) | ( x118 & ~n10024 ) | ( n10003 & ~n10024 ) ;
  assign n10354 = x118 & n10003 ;
  assign n10355 = ( ~n10008 & n10353 ) | ( ~n10008 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10356 = ( n10008 & n10353 ) | ( n10008 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10357 = ( n10008 & n10355 ) | ( n10008 & ~n10356 ) | ( n10355 & ~n10356 ) ;
  assign n10358 = ( x119 & n10352 ) | ( x119 & ~n10357 ) | ( n10352 & ~n10357 ) ;
  assign n10359 = ( x119 & n10009 ) | ( x119 & ~n10024 ) | ( n10009 & ~n10024 ) ;
  assign n10360 = x119 & n10009 ;
  assign n10361 = ( ~n10014 & n10359 ) | ( ~n10014 & n10360 ) | ( n10359 & n10360 ) ;
  assign n10362 = ( n10014 & n10359 ) | ( n10014 & n10360 ) | ( n10359 & n10360 ) ;
  assign n10363 = ( n10014 & n10361 ) | ( n10014 & ~n10362 ) | ( n10361 & ~n10362 ) ;
  assign n10364 = ( x120 & n10358 ) | ( x120 & ~n10363 ) | ( n10358 & ~n10363 ) ;
  assign n10365 = ( x121 & ~n10029 ) | ( x121 & n10364 ) | ( ~n10029 & n10364 ) ;
  assign n10366 = n135 & ~n10021 ;
  assign n10367 = x121 & n10022 ;
  assign n10368 = n389 | n10367 ;
  assign n10369 = ( n389 & n10016 ) | ( n389 & n10368 ) | ( n10016 & n10368 ) ;
  assign n10370 = ~n10366 & n10369 ;
  assign n10371 = ( n10365 & n10366 ) | ( n10365 & ~n10370 ) | ( n10366 & ~n10370 ) ;
  assign n10372 = ( x121 & n10364 ) | ( x121 & n10371 ) | ( n10364 & n10371 ) ;
  assign n10373 = x121 | n10364 ;
  assign n10374 = ( ~n10029 & n10372 ) | ( ~n10029 & n10373 ) | ( n10372 & n10373 ) ;
  assign n10375 = ( n10029 & n10372 ) | ( n10029 & n10373 ) | ( n10372 & n10373 ) ;
  assign n10376 = ( n10029 & n10374 ) | ( n10029 & ~n10375 ) | ( n10374 & ~n10375 ) ;
  assign n10377 = ~x4 & x64 ;
  assign n10378 = ~x5 & n10371 ;
  assign n10379 = ( x5 & ~x64 ) | ( x5 & n10371 ) | ( ~x64 & n10371 ) ;
  assign n10380 = ( n10030 & ~n10378 ) | ( n10030 & n10379 ) | ( ~n10378 & n10379 ) ;
  assign n10381 = ( x65 & n10377 ) | ( x65 & ~n10380 ) | ( n10377 & ~n10380 ) ;
  assign n10382 = ( x65 & n10030 ) | ( x65 & n10371 ) | ( n10030 & n10371 ) ;
  assign n10383 = x65 | n10030 ;
  assign n10384 = ( ~n10033 & n10382 ) | ( ~n10033 & n10383 ) | ( n10382 & n10383 ) ;
  assign n10385 = ( n10033 & n10382 ) | ( n10033 & n10383 ) | ( n10382 & n10383 ) ;
  assign n10386 = ( n10033 & n10384 ) | ( n10033 & ~n10385 ) | ( n10384 & ~n10385 ) ;
  assign n10387 = ( x66 & n10381 ) | ( x66 & ~n10386 ) | ( n10381 & ~n10386 ) ;
  assign n10388 = ( x66 & n10034 ) | ( x66 & n10371 ) | ( n10034 & n10371 ) ;
  assign n10389 = x66 | n10034 ;
  assign n10390 = ( ~n10039 & n10388 ) | ( ~n10039 & n10389 ) | ( n10388 & n10389 ) ;
  assign n10391 = ( n10039 & n10388 ) | ( n10039 & n10389 ) | ( n10388 & n10389 ) ;
  assign n10392 = ( n10039 & n10390 ) | ( n10039 & ~n10391 ) | ( n10390 & ~n10391 ) ;
  assign n10393 = ( x67 & n10387 ) | ( x67 & ~n10392 ) | ( n10387 & ~n10392 ) ;
  assign n10394 = ( x67 & n10040 ) | ( x67 & ~n10371 ) | ( n10040 & ~n10371 ) ;
  assign n10395 = x67 & n10040 ;
  assign n10396 = ( ~n10045 & n10394 ) | ( ~n10045 & n10395 ) | ( n10394 & n10395 ) ;
  assign n10397 = ( n10045 & n10394 ) | ( n10045 & n10395 ) | ( n10394 & n10395 ) ;
  assign n10398 = ( n10045 & n10396 ) | ( n10045 & ~n10397 ) | ( n10396 & ~n10397 ) ;
  assign n10399 = ( x68 & n10393 ) | ( x68 & ~n10398 ) | ( n10393 & ~n10398 ) ;
  assign n10400 = ( x68 & n10046 ) | ( x68 & ~n10371 ) | ( n10046 & ~n10371 ) ;
  assign n10401 = x68 & n10046 ;
  assign n10402 = ( ~n10051 & n10400 ) | ( ~n10051 & n10401 ) | ( n10400 & n10401 ) ;
  assign n10403 = ( n10051 & n10400 ) | ( n10051 & n10401 ) | ( n10400 & n10401 ) ;
  assign n10404 = ( n10051 & n10402 ) | ( n10051 & ~n10403 ) | ( n10402 & ~n10403 ) ;
  assign n10405 = ( x69 & n10399 ) | ( x69 & ~n10404 ) | ( n10399 & ~n10404 ) ;
  assign n10406 = ( x69 & n10052 ) | ( x69 & ~n10371 ) | ( n10052 & ~n10371 ) ;
  assign n10407 = x69 & n10052 ;
  assign n10408 = ( ~n10057 & n10406 ) | ( ~n10057 & n10407 ) | ( n10406 & n10407 ) ;
  assign n10409 = ( n10057 & n10406 ) | ( n10057 & n10407 ) | ( n10406 & n10407 ) ;
  assign n10410 = ( n10057 & n10408 ) | ( n10057 & ~n10409 ) | ( n10408 & ~n10409 ) ;
  assign n10411 = ( x70 & n10405 ) | ( x70 & ~n10410 ) | ( n10405 & ~n10410 ) ;
  assign n10412 = ( x70 & n10058 ) | ( x70 & ~n10371 ) | ( n10058 & ~n10371 ) ;
  assign n10413 = x70 & n10058 ;
  assign n10414 = ( ~n10063 & n10412 ) | ( ~n10063 & n10413 ) | ( n10412 & n10413 ) ;
  assign n10415 = ( n10063 & n10412 ) | ( n10063 & n10413 ) | ( n10412 & n10413 ) ;
  assign n10416 = ( n10063 & n10414 ) | ( n10063 & ~n10415 ) | ( n10414 & ~n10415 ) ;
  assign n10417 = ( x71 & n10411 ) | ( x71 & ~n10416 ) | ( n10411 & ~n10416 ) ;
  assign n10418 = ( x71 & n10064 ) | ( x71 & ~n10371 ) | ( n10064 & ~n10371 ) ;
  assign n10419 = x71 & n10064 ;
  assign n10420 = ( ~n10069 & n10418 ) | ( ~n10069 & n10419 ) | ( n10418 & n10419 ) ;
  assign n10421 = ( n10069 & n10418 ) | ( n10069 & n10419 ) | ( n10418 & n10419 ) ;
  assign n10422 = ( n10069 & n10420 ) | ( n10069 & ~n10421 ) | ( n10420 & ~n10421 ) ;
  assign n10423 = ( x72 & n10417 ) | ( x72 & ~n10422 ) | ( n10417 & ~n10422 ) ;
  assign n10424 = ( x72 & n10070 ) | ( x72 & ~n10371 ) | ( n10070 & ~n10371 ) ;
  assign n10425 = x72 & n10070 ;
  assign n10426 = ( ~n10075 & n10424 ) | ( ~n10075 & n10425 ) | ( n10424 & n10425 ) ;
  assign n10427 = ( n10075 & n10424 ) | ( n10075 & n10425 ) | ( n10424 & n10425 ) ;
  assign n10428 = ( n10075 & n10426 ) | ( n10075 & ~n10427 ) | ( n10426 & ~n10427 ) ;
  assign n10429 = ( x73 & n10423 ) | ( x73 & ~n10428 ) | ( n10423 & ~n10428 ) ;
  assign n10430 = ( x73 & n10076 ) | ( x73 & ~n10371 ) | ( n10076 & ~n10371 ) ;
  assign n10431 = x73 & n10076 ;
  assign n10432 = ( ~n10081 & n10430 ) | ( ~n10081 & n10431 ) | ( n10430 & n10431 ) ;
  assign n10433 = ( n10081 & n10430 ) | ( n10081 & n10431 ) | ( n10430 & n10431 ) ;
  assign n10434 = ( n10081 & n10432 ) | ( n10081 & ~n10433 ) | ( n10432 & ~n10433 ) ;
  assign n10435 = ( x74 & n10429 ) | ( x74 & ~n10434 ) | ( n10429 & ~n10434 ) ;
  assign n10436 = ( x74 & n10082 ) | ( x74 & ~n10371 ) | ( n10082 & ~n10371 ) ;
  assign n10437 = x74 & n10082 ;
  assign n10438 = ( ~n10087 & n10436 ) | ( ~n10087 & n10437 ) | ( n10436 & n10437 ) ;
  assign n10439 = ( n10087 & n10436 ) | ( n10087 & n10437 ) | ( n10436 & n10437 ) ;
  assign n10440 = ( n10087 & n10438 ) | ( n10087 & ~n10439 ) | ( n10438 & ~n10439 ) ;
  assign n10441 = ( x75 & n10435 ) | ( x75 & ~n10440 ) | ( n10435 & ~n10440 ) ;
  assign n10442 = ( x75 & n10088 ) | ( x75 & ~n10371 ) | ( n10088 & ~n10371 ) ;
  assign n10443 = x75 & n10088 ;
  assign n10444 = ( ~n10093 & n10442 ) | ( ~n10093 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10445 = ( n10093 & n10442 ) | ( n10093 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10446 = ( n10093 & n10444 ) | ( n10093 & ~n10445 ) | ( n10444 & ~n10445 ) ;
  assign n10447 = ( x76 & n10441 ) | ( x76 & ~n10446 ) | ( n10441 & ~n10446 ) ;
  assign n10448 = ( x76 & n10094 ) | ( x76 & ~n10371 ) | ( n10094 & ~n10371 ) ;
  assign n10449 = x76 & n10094 ;
  assign n10450 = ( ~n10099 & n10448 ) | ( ~n10099 & n10449 ) | ( n10448 & n10449 ) ;
  assign n10451 = ( n10099 & n10448 ) | ( n10099 & n10449 ) | ( n10448 & n10449 ) ;
  assign n10452 = ( n10099 & n10450 ) | ( n10099 & ~n10451 ) | ( n10450 & ~n10451 ) ;
  assign n10453 = ( x77 & n10447 ) | ( x77 & ~n10452 ) | ( n10447 & ~n10452 ) ;
  assign n10454 = ( x77 & n10100 ) | ( x77 & ~n10371 ) | ( n10100 & ~n10371 ) ;
  assign n10455 = x77 & n10100 ;
  assign n10456 = ( ~n10105 & n10454 ) | ( ~n10105 & n10455 ) | ( n10454 & n10455 ) ;
  assign n10457 = ( n10105 & n10454 ) | ( n10105 & n10455 ) | ( n10454 & n10455 ) ;
  assign n10458 = ( n10105 & n10456 ) | ( n10105 & ~n10457 ) | ( n10456 & ~n10457 ) ;
  assign n10459 = ( x78 & n10453 ) | ( x78 & ~n10458 ) | ( n10453 & ~n10458 ) ;
  assign n10460 = ( x78 & n10106 ) | ( x78 & ~n10371 ) | ( n10106 & ~n10371 ) ;
  assign n10461 = x78 & n10106 ;
  assign n10462 = ( ~n10111 & n10460 ) | ( ~n10111 & n10461 ) | ( n10460 & n10461 ) ;
  assign n10463 = ( n10111 & n10460 ) | ( n10111 & n10461 ) | ( n10460 & n10461 ) ;
  assign n10464 = ( n10111 & n10462 ) | ( n10111 & ~n10463 ) | ( n10462 & ~n10463 ) ;
  assign n10465 = ( x79 & n10459 ) | ( x79 & ~n10464 ) | ( n10459 & ~n10464 ) ;
  assign n10466 = ( x79 & n10112 ) | ( x79 & ~n10371 ) | ( n10112 & ~n10371 ) ;
  assign n10467 = x79 & n10112 ;
  assign n10468 = ( ~n10117 & n10466 ) | ( ~n10117 & n10467 ) | ( n10466 & n10467 ) ;
  assign n10469 = ( n10117 & n10466 ) | ( n10117 & n10467 ) | ( n10466 & n10467 ) ;
  assign n10470 = ( n10117 & n10468 ) | ( n10117 & ~n10469 ) | ( n10468 & ~n10469 ) ;
  assign n10471 = ( x80 & n10465 ) | ( x80 & ~n10470 ) | ( n10465 & ~n10470 ) ;
  assign n10472 = ( x80 & n10118 ) | ( x80 & ~n10371 ) | ( n10118 & ~n10371 ) ;
  assign n10473 = x80 & n10118 ;
  assign n10474 = ( ~n10123 & n10472 ) | ( ~n10123 & n10473 ) | ( n10472 & n10473 ) ;
  assign n10475 = ( n10123 & n10472 ) | ( n10123 & n10473 ) | ( n10472 & n10473 ) ;
  assign n10476 = ( n10123 & n10474 ) | ( n10123 & ~n10475 ) | ( n10474 & ~n10475 ) ;
  assign n10477 = ( x81 & n10471 ) | ( x81 & ~n10476 ) | ( n10471 & ~n10476 ) ;
  assign n10478 = ( x81 & n10124 ) | ( x81 & ~n10371 ) | ( n10124 & ~n10371 ) ;
  assign n10479 = x81 & n10124 ;
  assign n10480 = ( ~n10129 & n10478 ) | ( ~n10129 & n10479 ) | ( n10478 & n10479 ) ;
  assign n10481 = ( n10129 & n10478 ) | ( n10129 & n10479 ) | ( n10478 & n10479 ) ;
  assign n10482 = ( n10129 & n10480 ) | ( n10129 & ~n10481 ) | ( n10480 & ~n10481 ) ;
  assign n10483 = ( x82 & n10477 ) | ( x82 & ~n10482 ) | ( n10477 & ~n10482 ) ;
  assign n10484 = ( x82 & n10130 ) | ( x82 & ~n10371 ) | ( n10130 & ~n10371 ) ;
  assign n10485 = x82 & n10130 ;
  assign n10486 = ( ~n10135 & n10484 ) | ( ~n10135 & n10485 ) | ( n10484 & n10485 ) ;
  assign n10487 = ( n10135 & n10484 ) | ( n10135 & n10485 ) | ( n10484 & n10485 ) ;
  assign n10488 = ( n10135 & n10486 ) | ( n10135 & ~n10487 ) | ( n10486 & ~n10487 ) ;
  assign n10489 = ( x83 & n10483 ) | ( x83 & ~n10488 ) | ( n10483 & ~n10488 ) ;
  assign n10490 = ( x83 & n10136 ) | ( x83 & ~n10371 ) | ( n10136 & ~n10371 ) ;
  assign n10491 = x83 & n10136 ;
  assign n10492 = ( ~n10141 & n10490 ) | ( ~n10141 & n10491 ) | ( n10490 & n10491 ) ;
  assign n10493 = ( n10141 & n10490 ) | ( n10141 & n10491 ) | ( n10490 & n10491 ) ;
  assign n10494 = ( n10141 & n10492 ) | ( n10141 & ~n10493 ) | ( n10492 & ~n10493 ) ;
  assign n10495 = ( x84 & n10489 ) | ( x84 & ~n10494 ) | ( n10489 & ~n10494 ) ;
  assign n10496 = ( x84 & n10142 ) | ( x84 & ~n10371 ) | ( n10142 & ~n10371 ) ;
  assign n10497 = x84 & n10142 ;
  assign n10498 = ( ~n10147 & n10496 ) | ( ~n10147 & n10497 ) | ( n10496 & n10497 ) ;
  assign n10499 = ( n10147 & n10496 ) | ( n10147 & n10497 ) | ( n10496 & n10497 ) ;
  assign n10500 = ( n10147 & n10498 ) | ( n10147 & ~n10499 ) | ( n10498 & ~n10499 ) ;
  assign n10501 = ( x85 & n10495 ) | ( x85 & ~n10500 ) | ( n10495 & ~n10500 ) ;
  assign n10502 = ( x85 & n10148 ) | ( x85 & ~n10371 ) | ( n10148 & ~n10371 ) ;
  assign n10503 = x85 & n10148 ;
  assign n10504 = ( ~n10153 & n10502 ) | ( ~n10153 & n10503 ) | ( n10502 & n10503 ) ;
  assign n10505 = ( n10153 & n10502 ) | ( n10153 & n10503 ) | ( n10502 & n10503 ) ;
  assign n10506 = ( n10153 & n10504 ) | ( n10153 & ~n10505 ) | ( n10504 & ~n10505 ) ;
  assign n10507 = ( x86 & n10501 ) | ( x86 & ~n10506 ) | ( n10501 & ~n10506 ) ;
  assign n10508 = ( x86 & n10154 ) | ( x86 & ~n10371 ) | ( n10154 & ~n10371 ) ;
  assign n10509 = x86 & n10154 ;
  assign n10510 = ( ~n10159 & n10508 ) | ( ~n10159 & n10509 ) | ( n10508 & n10509 ) ;
  assign n10511 = ( n10159 & n10508 ) | ( n10159 & n10509 ) | ( n10508 & n10509 ) ;
  assign n10512 = ( n10159 & n10510 ) | ( n10159 & ~n10511 ) | ( n10510 & ~n10511 ) ;
  assign n10513 = ( x87 & n10507 ) | ( x87 & ~n10512 ) | ( n10507 & ~n10512 ) ;
  assign n10514 = ( x87 & n10160 ) | ( x87 & ~n10371 ) | ( n10160 & ~n10371 ) ;
  assign n10515 = x87 & n10160 ;
  assign n10516 = ( ~n10165 & n10514 ) | ( ~n10165 & n10515 ) | ( n10514 & n10515 ) ;
  assign n10517 = ( n10165 & n10514 ) | ( n10165 & n10515 ) | ( n10514 & n10515 ) ;
  assign n10518 = ( n10165 & n10516 ) | ( n10165 & ~n10517 ) | ( n10516 & ~n10517 ) ;
  assign n10519 = ( x88 & n10513 ) | ( x88 & ~n10518 ) | ( n10513 & ~n10518 ) ;
  assign n10520 = ( x88 & n10166 ) | ( x88 & ~n10371 ) | ( n10166 & ~n10371 ) ;
  assign n10521 = x88 & n10166 ;
  assign n10522 = ( ~n10171 & n10520 ) | ( ~n10171 & n10521 ) | ( n10520 & n10521 ) ;
  assign n10523 = ( n10171 & n10520 ) | ( n10171 & n10521 ) | ( n10520 & n10521 ) ;
  assign n10524 = ( n10171 & n10522 ) | ( n10171 & ~n10523 ) | ( n10522 & ~n10523 ) ;
  assign n10525 = ( x89 & n10519 ) | ( x89 & ~n10524 ) | ( n10519 & ~n10524 ) ;
  assign n10526 = ( x89 & n10172 ) | ( x89 & ~n10371 ) | ( n10172 & ~n10371 ) ;
  assign n10527 = x89 & n10172 ;
  assign n10528 = ( ~n10177 & n10526 ) | ( ~n10177 & n10527 ) | ( n10526 & n10527 ) ;
  assign n10529 = ( n10177 & n10526 ) | ( n10177 & n10527 ) | ( n10526 & n10527 ) ;
  assign n10530 = ( n10177 & n10528 ) | ( n10177 & ~n10529 ) | ( n10528 & ~n10529 ) ;
  assign n10531 = ( x90 & n10525 ) | ( x90 & ~n10530 ) | ( n10525 & ~n10530 ) ;
  assign n10532 = ( x90 & n10178 ) | ( x90 & ~n10371 ) | ( n10178 & ~n10371 ) ;
  assign n10533 = x90 & n10178 ;
  assign n10534 = ( ~n10183 & n10532 ) | ( ~n10183 & n10533 ) | ( n10532 & n10533 ) ;
  assign n10535 = ( n10183 & n10532 ) | ( n10183 & n10533 ) | ( n10532 & n10533 ) ;
  assign n10536 = ( n10183 & n10534 ) | ( n10183 & ~n10535 ) | ( n10534 & ~n10535 ) ;
  assign n10537 = ( x91 & n10531 ) | ( x91 & ~n10536 ) | ( n10531 & ~n10536 ) ;
  assign n10538 = ( x91 & n10184 ) | ( x91 & ~n10371 ) | ( n10184 & ~n10371 ) ;
  assign n10539 = x91 & n10184 ;
  assign n10540 = ( ~n10189 & n10538 ) | ( ~n10189 & n10539 ) | ( n10538 & n10539 ) ;
  assign n10541 = ( n10189 & n10538 ) | ( n10189 & n10539 ) | ( n10538 & n10539 ) ;
  assign n10542 = ( n10189 & n10540 ) | ( n10189 & ~n10541 ) | ( n10540 & ~n10541 ) ;
  assign n10543 = ( x92 & n10537 ) | ( x92 & ~n10542 ) | ( n10537 & ~n10542 ) ;
  assign n10544 = ( x92 & n10190 ) | ( x92 & ~n10371 ) | ( n10190 & ~n10371 ) ;
  assign n10545 = x92 & n10190 ;
  assign n10546 = ( ~n10195 & n10544 ) | ( ~n10195 & n10545 ) | ( n10544 & n10545 ) ;
  assign n10547 = ( n10195 & n10544 ) | ( n10195 & n10545 ) | ( n10544 & n10545 ) ;
  assign n10548 = ( n10195 & n10546 ) | ( n10195 & ~n10547 ) | ( n10546 & ~n10547 ) ;
  assign n10549 = ( x93 & n10543 ) | ( x93 & ~n10548 ) | ( n10543 & ~n10548 ) ;
  assign n10550 = ( x93 & n10196 ) | ( x93 & ~n10371 ) | ( n10196 & ~n10371 ) ;
  assign n10551 = x93 & n10196 ;
  assign n10552 = ( ~n10201 & n10550 ) | ( ~n10201 & n10551 ) | ( n10550 & n10551 ) ;
  assign n10553 = ( n10201 & n10550 ) | ( n10201 & n10551 ) | ( n10550 & n10551 ) ;
  assign n10554 = ( n10201 & n10552 ) | ( n10201 & ~n10553 ) | ( n10552 & ~n10553 ) ;
  assign n10555 = ( x94 & n10549 ) | ( x94 & ~n10554 ) | ( n10549 & ~n10554 ) ;
  assign n10556 = ( x94 & n10202 ) | ( x94 & ~n10371 ) | ( n10202 & ~n10371 ) ;
  assign n10557 = x94 & n10202 ;
  assign n10558 = ( ~n10207 & n10556 ) | ( ~n10207 & n10557 ) | ( n10556 & n10557 ) ;
  assign n10559 = ( n10207 & n10556 ) | ( n10207 & n10557 ) | ( n10556 & n10557 ) ;
  assign n10560 = ( n10207 & n10558 ) | ( n10207 & ~n10559 ) | ( n10558 & ~n10559 ) ;
  assign n10561 = ( x95 & n10555 ) | ( x95 & ~n10560 ) | ( n10555 & ~n10560 ) ;
  assign n10562 = ( x95 & n10208 ) | ( x95 & ~n10371 ) | ( n10208 & ~n10371 ) ;
  assign n10563 = x95 & n10208 ;
  assign n10564 = ( ~n10213 & n10562 ) | ( ~n10213 & n10563 ) | ( n10562 & n10563 ) ;
  assign n10565 = ( n10213 & n10562 ) | ( n10213 & n10563 ) | ( n10562 & n10563 ) ;
  assign n10566 = ( n10213 & n10564 ) | ( n10213 & ~n10565 ) | ( n10564 & ~n10565 ) ;
  assign n10567 = ( x96 & n10561 ) | ( x96 & ~n10566 ) | ( n10561 & ~n10566 ) ;
  assign n10568 = ( x96 & n10214 ) | ( x96 & ~n10371 ) | ( n10214 & ~n10371 ) ;
  assign n10569 = x96 & n10214 ;
  assign n10570 = ( ~n10219 & n10568 ) | ( ~n10219 & n10569 ) | ( n10568 & n10569 ) ;
  assign n10571 = ( n10219 & n10568 ) | ( n10219 & n10569 ) | ( n10568 & n10569 ) ;
  assign n10572 = ( n10219 & n10570 ) | ( n10219 & ~n10571 ) | ( n10570 & ~n10571 ) ;
  assign n10573 = ( x97 & n10567 ) | ( x97 & ~n10572 ) | ( n10567 & ~n10572 ) ;
  assign n10574 = ( x97 & n10220 ) | ( x97 & ~n10371 ) | ( n10220 & ~n10371 ) ;
  assign n10575 = x97 & n10220 ;
  assign n10576 = ( ~n10225 & n10574 ) | ( ~n10225 & n10575 ) | ( n10574 & n10575 ) ;
  assign n10577 = ( n10225 & n10574 ) | ( n10225 & n10575 ) | ( n10574 & n10575 ) ;
  assign n10578 = ( n10225 & n10576 ) | ( n10225 & ~n10577 ) | ( n10576 & ~n10577 ) ;
  assign n10579 = ( x98 & n10573 ) | ( x98 & ~n10578 ) | ( n10573 & ~n10578 ) ;
  assign n10580 = ( x98 & n10226 ) | ( x98 & ~n10371 ) | ( n10226 & ~n10371 ) ;
  assign n10581 = x98 & n10226 ;
  assign n10582 = ( ~n10231 & n10580 ) | ( ~n10231 & n10581 ) | ( n10580 & n10581 ) ;
  assign n10583 = ( n10231 & n10580 ) | ( n10231 & n10581 ) | ( n10580 & n10581 ) ;
  assign n10584 = ( n10231 & n10582 ) | ( n10231 & ~n10583 ) | ( n10582 & ~n10583 ) ;
  assign n10585 = ( x99 & n10579 ) | ( x99 & ~n10584 ) | ( n10579 & ~n10584 ) ;
  assign n10586 = ( x99 & n10232 ) | ( x99 & ~n10371 ) | ( n10232 & ~n10371 ) ;
  assign n10587 = x99 & n10232 ;
  assign n10588 = ( ~n10237 & n10586 ) | ( ~n10237 & n10587 ) | ( n10586 & n10587 ) ;
  assign n10589 = ( n10237 & n10586 ) | ( n10237 & n10587 ) | ( n10586 & n10587 ) ;
  assign n10590 = ( n10237 & n10588 ) | ( n10237 & ~n10589 ) | ( n10588 & ~n10589 ) ;
  assign n10591 = ( x100 & n10585 ) | ( x100 & ~n10590 ) | ( n10585 & ~n10590 ) ;
  assign n10592 = ( x100 & n10238 ) | ( x100 & ~n10371 ) | ( n10238 & ~n10371 ) ;
  assign n10593 = x100 & n10238 ;
  assign n10594 = ( ~n10243 & n10592 ) | ( ~n10243 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10595 = ( n10243 & n10592 ) | ( n10243 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10596 = ( n10243 & n10594 ) | ( n10243 & ~n10595 ) | ( n10594 & ~n10595 ) ;
  assign n10597 = ( x101 & n10591 ) | ( x101 & ~n10596 ) | ( n10591 & ~n10596 ) ;
  assign n10598 = ( x101 & n10244 ) | ( x101 & ~n10371 ) | ( n10244 & ~n10371 ) ;
  assign n10599 = x101 & n10244 ;
  assign n10600 = ( ~n10249 & n10598 ) | ( ~n10249 & n10599 ) | ( n10598 & n10599 ) ;
  assign n10601 = ( n10249 & n10598 ) | ( n10249 & n10599 ) | ( n10598 & n10599 ) ;
  assign n10602 = ( n10249 & n10600 ) | ( n10249 & ~n10601 ) | ( n10600 & ~n10601 ) ;
  assign n10603 = ( x102 & n10597 ) | ( x102 & ~n10602 ) | ( n10597 & ~n10602 ) ;
  assign n10604 = ( x102 & n10250 ) | ( x102 & ~n10371 ) | ( n10250 & ~n10371 ) ;
  assign n10605 = x102 & n10250 ;
  assign n10606 = ( ~n10255 & n10604 ) | ( ~n10255 & n10605 ) | ( n10604 & n10605 ) ;
  assign n10607 = ( n10255 & n10604 ) | ( n10255 & n10605 ) | ( n10604 & n10605 ) ;
  assign n10608 = ( n10255 & n10606 ) | ( n10255 & ~n10607 ) | ( n10606 & ~n10607 ) ;
  assign n10609 = ( x103 & n10603 ) | ( x103 & ~n10608 ) | ( n10603 & ~n10608 ) ;
  assign n10610 = ( x103 & n10256 ) | ( x103 & ~n10371 ) | ( n10256 & ~n10371 ) ;
  assign n10611 = x103 & n10256 ;
  assign n10612 = ( ~n10261 & n10610 ) | ( ~n10261 & n10611 ) | ( n10610 & n10611 ) ;
  assign n10613 = ( n10261 & n10610 ) | ( n10261 & n10611 ) | ( n10610 & n10611 ) ;
  assign n10614 = ( n10261 & n10612 ) | ( n10261 & ~n10613 ) | ( n10612 & ~n10613 ) ;
  assign n10615 = ( x104 & n10609 ) | ( x104 & ~n10614 ) | ( n10609 & ~n10614 ) ;
  assign n10616 = ( x104 & n10262 ) | ( x104 & ~n10371 ) | ( n10262 & ~n10371 ) ;
  assign n10617 = x104 & n10262 ;
  assign n10618 = ( ~n10267 & n10616 ) | ( ~n10267 & n10617 ) | ( n10616 & n10617 ) ;
  assign n10619 = ( n10267 & n10616 ) | ( n10267 & n10617 ) | ( n10616 & n10617 ) ;
  assign n10620 = ( n10267 & n10618 ) | ( n10267 & ~n10619 ) | ( n10618 & ~n10619 ) ;
  assign n10621 = ( x105 & n10615 ) | ( x105 & ~n10620 ) | ( n10615 & ~n10620 ) ;
  assign n10622 = ( x105 & n10268 ) | ( x105 & ~n10371 ) | ( n10268 & ~n10371 ) ;
  assign n10623 = x105 & n10268 ;
  assign n10624 = ( ~n10273 & n10622 ) | ( ~n10273 & n10623 ) | ( n10622 & n10623 ) ;
  assign n10625 = ( n10273 & n10622 ) | ( n10273 & n10623 ) | ( n10622 & n10623 ) ;
  assign n10626 = ( n10273 & n10624 ) | ( n10273 & ~n10625 ) | ( n10624 & ~n10625 ) ;
  assign n10627 = ( x106 & n10621 ) | ( x106 & ~n10626 ) | ( n10621 & ~n10626 ) ;
  assign n10628 = ( x106 & n10274 ) | ( x106 & ~n10371 ) | ( n10274 & ~n10371 ) ;
  assign n10629 = x106 & n10274 ;
  assign n10630 = ( ~n10279 & n10628 ) | ( ~n10279 & n10629 ) | ( n10628 & n10629 ) ;
  assign n10631 = ( n10279 & n10628 ) | ( n10279 & n10629 ) | ( n10628 & n10629 ) ;
  assign n10632 = ( n10279 & n10630 ) | ( n10279 & ~n10631 ) | ( n10630 & ~n10631 ) ;
  assign n10633 = ( x107 & n10627 ) | ( x107 & ~n10632 ) | ( n10627 & ~n10632 ) ;
  assign n10634 = ( x107 & n10280 ) | ( x107 & ~n10371 ) | ( n10280 & ~n10371 ) ;
  assign n10635 = x107 & n10280 ;
  assign n10636 = ( ~n10285 & n10634 ) | ( ~n10285 & n10635 ) | ( n10634 & n10635 ) ;
  assign n10637 = ( n10285 & n10634 ) | ( n10285 & n10635 ) | ( n10634 & n10635 ) ;
  assign n10638 = ( n10285 & n10636 ) | ( n10285 & ~n10637 ) | ( n10636 & ~n10637 ) ;
  assign n10639 = ( x108 & n10633 ) | ( x108 & ~n10638 ) | ( n10633 & ~n10638 ) ;
  assign n10640 = ( x108 & n10286 ) | ( x108 & ~n10371 ) | ( n10286 & ~n10371 ) ;
  assign n10641 = x108 & n10286 ;
  assign n10642 = ( ~n10291 & n10640 ) | ( ~n10291 & n10641 ) | ( n10640 & n10641 ) ;
  assign n10643 = ( n10291 & n10640 ) | ( n10291 & n10641 ) | ( n10640 & n10641 ) ;
  assign n10644 = ( n10291 & n10642 ) | ( n10291 & ~n10643 ) | ( n10642 & ~n10643 ) ;
  assign n10645 = ( x109 & n10639 ) | ( x109 & ~n10644 ) | ( n10639 & ~n10644 ) ;
  assign n10646 = ( x109 & n10292 ) | ( x109 & ~n10371 ) | ( n10292 & ~n10371 ) ;
  assign n10647 = x109 & n10292 ;
  assign n10648 = ( ~n10297 & n10646 ) | ( ~n10297 & n10647 ) | ( n10646 & n10647 ) ;
  assign n10649 = ( n10297 & n10646 ) | ( n10297 & n10647 ) | ( n10646 & n10647 ) ;
  assign n10650 = ( n10297 & n10648 ) | ( n10297 & ~n10649 ) | ( n10648 & ~n10649 ) ;
  assign n10651 = ( x110 & n10645 ) | ( x110 & ~n10650 ) | ( n10645 & ~n10650 ) ;
  assign n10652 = ( x110 & n10298 ) | ( x110 & ~n10371 ) | ( n10298 & ~n10371 ) ;
  assign n10653 = x110 & n10298 ;
  assign n10654 = ( ~n10303 & n10652 ) | ( ~n10303 & n10653 ) | ( n10652 & n10653 ) ;
  assign n10655 = ( n10303 & n10652 ) | ( n10303 & n10653 ) | ( n10652 & n10653 ) ;
  assign n10656 = ( n10303 & n10654 ) | ( n10303 & ~n10655 ) | ( n10654 & ~n10655 ) ;
  assign n10657 = ( x111 & n10651 ) | ( x111 & ~n10656 ) | ( n10651 & ~n10656 ) ;
  assign n10658 = ( x111 & n10304 ) | ( x111 & ~n10371 ) | ( n10304 & ~n10371 ) ;
  assign n10659 = x111 & n10304 ;
  assign n10660 = ( ~n10309 & n10658 ) | ( ~n10309 & n10659 ) | ( n10658 & n10659 ) ;
  assign n10661 = ( n10309 & n10658 ) | ( n10309 & n10659 ) | ( n10658 & n10659 ) ;
  assign n10662 = ( n10309 & n10660 ) | ( n10309 & ~n10661 ) | ( n10660 & ~n10661 ) ;
  assign n10663 = ( x112 & n10657 ) | ( x112 & ~n10662 ) | ( n10657 & ~n10662 ) ;
  assign n10664 = ( x112 & n10310 ) | ( x112 & ~n10371 ) | ( n10310 & ~n10371 ) ;
  assign n10665 = x112 & n10310 ;
  assign n10666 = ( ~n10315 & n10664 ) | ( ~n10315 & n10665 ) | ( n10664 & n10665 ) ;
  assign n10667 = ( n10315 & n10664 ) | ( n10315 & n10665 ) | ( n10664 & n10665 ) ;
  assign n10668 = ( n10315 & n10666 ) | ( n10315 & ~n10667 ) | ( n10666 & ~n10667 ) ;
  assign n10669 = ( x113 & n10663 ) | ( x113 & ~n10668 ) | ( n10663 & ~n10668 ) ;
  assign n10670 = ( x113 & n10316 ) | ( x113 & ~n10371 ) | ( n10316 & ~n10371 ) ;
  assign n10671 = x113 & n10316 ;
  assign n10672 = ( ~n10321 & n10670 ) | ( ~n10321 & n10671 ) | ( n10670 & n10671 ) ;
  assign n10673 = ( n10321 & n10670 ) | ( n10321 & n10671 ) | ( n10670 & n10671 ) ;
  assign n10674 = ( n10321 & n10672 ) | ( n10321 & ~n10673 ) | ( n10672 & ~n10673 ) ;
  assign n10675 = ( x114 & n10669 ) | ( x114 & ~n10674 ) | ( n10669 & ~n10674 ) ;
  assign n10676 = ( x114 & n10322 ) | ( x114 & ~n10371 ) | ( n10322 & ~n10371 ) ;
  assign n10677 = x114 & n10322 ;
  assign n10678 = ( ~n10327 & n10676 ) | ( ~n10327 & n10677 ) | ( n10676 & n10677 ) ;
  assign n10679 = ( n10327 & n10676 ) | ( n10327 & n10677 ) | ( n10676 & n10677 ) ;
  assign n10680 = ( n10327 & n10678 ) | ( n10327 & ~n10679 ) | ( n10678 & ~n10679 ) ;
  assign n10681 = ( x115 & n10675 ) | ( x115 & ~n10680 ) | ( n10675 & ~n10680 ) ;
  assign n10682 = ( x115 & n10328 ) | ( x115 & ~n10371 ) | ( n10328 & ~n10371 ) ;
  assign n10683 = x115 & n10328 ;
  assign n10684 = ( ~n10333 & n10682 ) | ( ~n10333 & n10683 ) | ( n10682 & n10683 ) ;
  assign n10685 = ( n10333 & n10682 ) | ( n10333 & n10683 ) | ( n10682 & n10683 ) ;
  assign n10686 = ( n10333 & n10684 ) | ( n10333 & ~n10685 ) | ( n10684 & ~n10685 ) ;
  assign n10687 = ( x116 & n10681 ) | ( x116 & ~n10686 ) | ( n10681 & ~n10686 ) ;
  assign n10688 = ( x116 & n10334 ) | ( x116 & ~n10371 ) | ( n10334 & ~n10371 ) ;
  assign n10689 = x116 & n10334 ;
  assign n10690 = ( ~n10339 & n10688 ) | ( ~n10339 & n10689 ) | ( n10688 & n10689 ) ;
  assign n10691 = ( n10339 & n10688 ) | ( n10339 & n10689 ) | ( n10688 & n10689 ) ;
  assign n10692 = ( n10339 & n10690 ) | ( n10339 & ~n10691 ) | ( n10690 & ~n10691 ) ;
  assign n10693 = ( x117 & n10687 ) | ( x117 & ~n10692 ) | ( n10687 & ~n10692 ) ;
  assign n10694 = ( x117 & n10340 ) | ( x117 & ~n10371 ) | ( n10340 & ~n10371 ) ;
  assign n10695 = x117 & n10340 ;
  assign n10696 = ( ~n10345 & n10694 ) | ( ~n10345 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = ( n10345 & n10694 ) | ( n10345 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10698 = ( n10345 & n10696 ) | ( n10345 & ~n10697 ) | ( n10696 & ~n10697 ) ;
  assign n10699 = ( x118 & n10693 ) | ( x118 & ~n10698 ) | ( n10693 & ~n10698 ) ;
  assign n10700 = ( x118 & n10346 ) | ( x118 & ~n10371 ) | ( n10346 & ~n10371 ) ;
  assign n10701 = x118 & n10346 ;
  assign n10702 = ( ~n10351 & n10700 ) | ( ~n10351 & n10701 ) | ( n10700 & n10701 ) ;
  assign n10703 = ( n10351 & n10700 ) | ( n10351 & n10701 ) | ( n10700 & n10701 ) ;
  assign n10704 = ( n10351 & n10702 ) | ( n10351 & ~n10703 ) | ( n10702 & ~n10703 ) ;
  assign n10705 = ( x119 & n10699 ) | ( x119 & ~n10704 ) | ( n10699 & ~n10704 ) ;
  assign n10706 = ( x119 & n10352 ) | ( x119 & ~n10371 ) | ( n10352 & ~n10371 ) ;
  assign n10707 = x119 & n10352 ;
  assign n10708 = ( ~n10357 & n10706 ) | ( ~n10357 & n10707 ) | ( n10706 & n10707 ) ;
  assign n10709 = ( n10357 & n10706 ) | ( n10357 & n10707 ) | ( n10706 & n10707 ) ;
  assign n10710 = ( n10357 & n10708 ) | ( n10357 & ~n10709 ) | ( n10708 & ~n10709 ) ;
  assign n10711 = ( x120 & n10705 ) | ( x120 & ~n10710 ) | ( n10705 & ~n10710 ) ;
  assign n10712 = ( x120 & n10358 ) | ( x120 & ~n10371 ) | ( n10358 & ~n10371 ) ;
  assign n10713 = x120 & n10358 ;
  assign n10714 = ( ~n10363 & n10712 ) | ( ~n10363 & n10713 ) | ( n10712 & n10713 ) ;
  assign n10715 = ( n10363 & n10712 ) | ( n10363 & n10713 ) | ( n10712 & n10713 ) ;
  assign n10716 = ( n10363 & n10714 ) | ( n10363 & ~n10715 ) | ( n10714 & ~n10715 ) ;
  assign n10717 = ( x121 & n10711 ) | ( x121 & ~n10716 ) | ( n10711 & ~n10716 ) ;
  assign n10718 = n134 | n389 ;
  assign n10719 = x122 | n10718 ;
  assign n10720 = ( n10365 & n10718 ) | ( n10365 & n10719 ) | ( n10718 & n10719 ) ;
  assign n10721 = n9679 & n10720 ;
  assign n10722 = ( x122 & ~n10376 ) | ( x122 & n10717 ) | ( ~n10376 & n10717 ) ;
  assign n10723 = ( x123 & ~n10721 ) | ( x123 & n10722 ) | ( ~n10721 & n10722 ) ;
  assign n10724 = n133 | n10723 ;
  assign n10725 = ( x122 & n10717 ) | ( x122 & n10724 ) | ( n10717 & n10724 ) ;
  assign n10726 = x122 | n10717 ;
  assign n10727 = ( ~n10376 & n10725 ) | ( ~n10376 & n10726 ) | ( n10725 & n10726 ) ;
  assign n10728 = ( n10376 & n10725 ) | ( n10376 & n10726 ) | ( n10725 & n10726 ) ;
  assign n10729 = ( n10376 & n10727 ) | ( n10376 & ~n10728 ) | ( n10727 & ~n10728 ) ;
  assign n10730 = ~x3 & x64 ;
  assign n10731 = ~x4 & n10724 ;
  assign n10732 = ( x4 & ~x64 ) | ( x4 & n10724 ) | ( ~x64 & n10724 ) ;
  assign n10733 = ( n10377 & ~n10731 ) | ( n10377 & n10732 ) | ( ~n10731 & n10732 ) ;
  assign n10734 = ( x65 & n10730 ) | ( x65 & ~n10733 ) | ( n10730 & ~n10733 ) ;
  assign n10735 = ( x65 & n10377 ) | ( x65 & n10724 ) | ( n10377 & n10724 ) ;
  assign n10736 = x65 | n10377 ;
  assign n10737 = ( ~n10380 & n10735 ) | ( ~n10380 & n10736 ) | ( n10735 & n10736 ) ;
  assign n10738 = ( n10380 & n10735 ) | ( n10380 & n10736 ) | ( n10735 & n10736 ) ;
  assign n10739 = ( n10380 & n10737 ) | ( n10380 & ~n10738 ) | ( n10737 & ~n10738 ) ;
  assign n10740 = ( x66 & n10734 ) | ( x66 & ~n10739 ) | ( n10734 & ~n10739 ) ;
  assign n10741 = ( x66 & n10381 ) | ( x66 & n10724 ) | ( n10381 & n10724 ) ;
  assign n10742 = x66 | n10381 ;
  assign n10743 = ( ~n10386 & n10741 ) | ( ~n10386 & n10742 ) | ( n10741 & n10742 ) ;
  assign n10744 = ( n10386 & n10741 ) | ( n10386 & n10742 ) | ( n10741 & n10742 ) ;
  assign n10745 = ( n10386 & n10743 ) | ( n10386 & ~n10744 ) | ( n10743 & ~n10744 ) ;
  assign n10746 = ( x67 & n10740 ) | ( x67 & ~n10745 ) | ( n10740 & ~n10745 ) ;
  assign n10747 = ( x67 & n10387 ) | ( x67 & ~n10724 ) | ( n10387 & ~n10724 ) ;
  assign n10748 = x67 & n10387 ;
  assign n10749 = ( ~n10392 & n10747 ) | ( ~n10392 & n10748 ) | ( n10747 & n10748 ) ;
  assign n10750 = ( n10392 & n10747 ) | ( n10392 & n10748 ) | ( n10747 & n10748 ) ;
  assign n10751 = ( n10392 & n10749 ) | ( n10392 & ~n10750 ) | ( n10749 & ~n10750 ) ;
  assign n10752 = ( x68 & n10746 ) | ( x68 & ~n10751 ) | ( n10746 & ~n10751 ) ;
  assign n10753 = ( x68 & n10393 ) | ( x68 & ~n10724 ) | ( n10393 & ~n10724 ) ;
  assign n10754 = x68 & n10393 ;
  assign n10755 = ( ~n10398 & n10753 ) | ( ~n10398 & n10754 ) | ( n10753 & n10754 ) ;
  assign n10756 = ( n10398 & n10753 ) | ( n10398 & n10754 ) | ( n10753 & n10754 ) ;
  assign n10757 = ( n10398 & n10755 ) | ( n10398 & ~n10756 ) | ( n10755 & ~n10756 ) ;
  assign n10758 = ( x69 & n10752 ) | ( x69 & ~n10757 ) | ( n10752 & ~n10757 ) ;
  assign n10759 = ( x69 & n10399 ) | ( x69 & ~n10724 ) | ( n10399 & ~n10724 ) ;
  assign n10760 = x69 & n10399 ;
  assign n10761 = ( ~n10404 & n10759 ) | ( ~n10404 & n10760 ) | ( n10759 & n10760 ) ;
  assign n10762 = ( n10404 & n10759 ) | ( n10404 & n10760 ) | ( n10759 & n10760 ) ;
  assign n10763 = ( n10404 & n10761 ) | ( n10404 & ~n10762 ) | ( n10761 & ~n10762 ) ;
  assign n10764 = ( x70 & n10758 ) | ( x70 & ~n10763 ) | ( n10758 & ~n10763 ) ;
  assign n10765 = ( x70 & n10405 ) | ( x70 & ~n10724 ) | ( n10405 & ~n10724 ) ;
  assign n10766 = x70 & n10405 ;
  assign n10767 = ( ~n10410 & n10765 ) | ( ~n10410 & n10766 ) | ( n10765 & n10766 ) ;
  assign n10768 = ( n10410 & n10765 ) | ( n10410 & n10766 ) | ( n10765 & n10766 ) ;
  assign n10769 = ( n10410 & n10767 ) | ( n10410 & ~n10768 ) | ( n10767 & ~n10768 ) ;
  assign n10770 = ( x71 & n10764 ) | ( x71 & ~n10769 ) | ( n10764 & ~n10769 ) ;
  assign n10771 = ( x71 & n10411 ) | ( x71 & ~n10724 ) | ( n10411 & ~n10724 ) ;
  assign n10772 = x71 & n10411 ;
  assign n10773 = ( ~n10416 & n10771 ) | ( ~n10416 & n10772 ) | ( n10771 & n10772 ) ;
  assign n10774 = ( n10416 & n10771 ) | ( n10416 & n10772 ) | ( n10771 & n10772 ) ;
  assign n10775 = ( n10416 & n10773 ) | ( n10416 & ~n10774 ) | ( n10773 & ~n10774 ) ;
  assign n10776 = ( x72 & n10770 ) | ( x72 & ~n10775 ) | ( n10770 & ~n10775 ) ;
  assign n10777 = ( x72 & n10417 ) | ( x72 & ~n10724 ) | ( n10417 & ~n10724 ) ;
  assign n10778 = x72 & n10417 ;
  assign n10779 = ( ~n10422 & n10777 ) | ( ~n10422 & n10778 ) | ( n10777 & n10778 ) ;
  assign n10780 = ( n10422 & n10777 ) | ( n10422 & n10778 ) | ( n10777 & n10778 ) ;
  assign n10781 = ( n10422 & n10779 ) | ( n10422 & ~n10780 ) | ( n10779 & ~n10780 ) ;
  assign n10782 = ( x73 & n10776 ) | ( x73 & ~n10781 ) | ( n10776 & ~n10781 ) ;
  assign n10783 = ( x73 & n10423 ) | ( x73 & ~n10724 ) | ( n10423 & ~n10724 ) ;
  assign n10784 = x73 & n10423 ;
  assign n10785 = ( ~n10428 & n10783 ) | ( ~n10428 & n10784 ) | ( n10783 & n10784 ) ;
  assign n10786 = ( n10428 & n10783 ) | ( n10428 & n10784 ) | ( n10783 & n10784 ) ;
  assign n10787 = ( n10428 & n10785 ) | ( n10428 & ~n10786 ) | ( n10785 & ~n10786 ) ;
  assign n10788 = ( x74 & n10782 ) | ( x74 & ~n10787 ) | ( n10782 & ~n10787 ) ;
  assign n10789 = ( x74 & n10429 ) | ( x74 & ~n10724 ) | ( n10429 & ~n10724 ) ;
  assign n10790 = x74 & n10429 ;
  assign n10791 = ( ~n10434 & n10789 ) | ( ~n10434 & n10790 ) | ( n10789 & n10790 ) ;
  assign n10792 = ( n10434 & n10789 ) | ( n10434 & n10790 ) | ( n10789 & n10790 ) ;
  assign n10793 = ( n10434 & n10791 ) | ( n10434 & ~n10792 ) | ( n10791 & ~n10792 ) ;
  assign n10794 = ( x75 & n10788 ) | ( x75 & ~n10793 ) | ( n10788 & ~n10793 ) ;
  assign n10795 = ( x75 & n10435 ) | ( x75 & ~n10724 ) | ( n10435 & ~n10724 ) ;
  assign n10796 = x75 & n10435 ;
  assign n10797 = ( ~n10440 & n10795 ) | ( ~n10440 & n10796 ) | ( n10795 & n10796 ) ;
  assign n10798 = ( n10440 & n10795 ) | ( n10440 & n10796 ) | ( n10795 & n10796 ) ;
  assign n10799 = ( n10440 & n10797 ) | ( n10440 & ~n10798 ) | ( n10797 & ~n10798 ) ;
  assign n10800 = ( x76 & n10794 ) | ( x76 & ~n10799 ) | ( n10794 & ~n10799 ) ;
  assign n10801 = ( x76 & n10441 ) | ( x76 & ~n10724 ) | ( n10441 & ~n10724 ) ;
  assign n10802 = x76 & n10441 ;
  assign n10803 = ( ~n10446 & n10801 ) | ( ~n10446 & n10802 ) | ( n10801 & n10802 ) ;
  assign n10804 = ( n10446 & n10801 ) | ( n10446 & n10802 ) | ( n10801 & n10802 ) ;
  assign n10805 = ( n10446 & n10803 ) | ( n10446 & ~n10804 ) | ( n10803 & ~n10804 ) ;
  assign n10806 = ( x77 & n10800 ) | ( x77 & ~n10805 ) | ( n10800 & ~n10805 ) ;
  assign n10807 = ( x77 & n10447 ) | ( x77 & ~n10724 ) | ( n10447 & ~n10724 ) ;
  assign n10808 = x77 & n10447 ;
  assign n10809 = ( ~n10452 & n10807 ) | ( ~n10452 & n10808 ) | ( n10807 & n10808 ) ;
  assign n10810 = ( n10452 & n10807 ) | ( n10452 & n10808 ) | ( n10807 & n10808 ) ;
  assign n10811 = ( n10452 & n10809 ) | ( n10452 & ~n10810 ) | ( n10809 & ~n10810 ) ;
  assign n10812 = ( x78 & n10806 ) | ( x78 & ~n10811 ) | ( n10806 & ~n10811 ) ;
  assign n10813 = ( x78 & n10453 ) | ( x78 & ~n10724 ) | ( n10453 & ~n10724 ) ;
  assign n10814 = x78 & n10453 ;
  assign n10815 = ( ~n10458 & n10813 ) | ( ~n10458 & n10814 ) | ( n10813 & n10814 ) ;
  assign n10816 = ( n10458 & n10813 ) | ( n10458 & n10814 ) | ( n10813 & n10814 ) ;
  assign n10817 = ( n10458 & n10815 ) | ( n10458 & ~n10816 ) | ( n10815 & ~n10816 ) ;
  assign n10818 = ( x79 & n10812 ) | ( x79 & ~n10817 ) | ( n10812 & ~n10817 ) ;
  assign n10819 = ( x79 & n10459 ) | ( x79 & ~n10724 ) | ( n10459 & ~n10724 ) ;
  assign n10820 = x79 & n10459 ;
  assign n10821 = ( ~n10464 & n10819 ) | ( ~n10464 & n10820 ) | ( n10819 & n10820 ) ;
  assign n10822 = ( n10464 & n10819 ) | ( n10464 & n10820 ) | ( n10819 & n10820 ) ;
  assign n10823 = ( n10464 & n10821 ) | ( n10464 & ~n10822 ) | ( n10821 & ~n10822 ) ;
  assign n10824 = ( x80 & n10818 ) | ( x80 & ~n10823 ) | ( n10818 & ~n10823 ) ;
  assign n10825 = ( x80 & n10465 ) | ( x80 & ~n10724 ) | ( n10465 & ~n10724 ) ;
  assign n10826 = x80 & n10465 ;
  assign n10827 = ( ~n10470 & n10825 ) | ( ~n10470 & n10826 ) | ( n10825 & n10826 ) ;
  assign n10828 = ( n10470 & n10825 ) | ( n10470 & n10826 ) | ( n10825 & n10826 ) ;
  assign n10829 = ( n10470 & n10827 ) | ( n10470 & ~n10828 ) | ( n10827 & ~n10828 ) ;
  assign n10830 = ( x81 & n10824 ) | ( x81 & ~n10829 ) | ( n10824 & ~n10829 ) ;
  assign n10831 = ( x81 & n10471 ) | ( x81 & ~n10724 ) | ( n10471 & ~n10724 ) ;
  assign n10832 = x81 & n10471 ;
  assign n10833 = ( ~n10476 & n10831 ) | ( ~n10476 & n10832 ) | ( n10831 & n10832 ) ;
  assign n10834 = ( n10476 & n10831 ) | ( n10476 & n10832 ) | ( n10831 & n10832 ) ;
  assign n10835 = ( n10476 & n10833 ) | ( n10476 & ~n10834 ) | ( n10833 & ~n10834 ) ;
  assign n10836 = ( x82 & n10830 ) | ( x82 & ~n10835 ) | ( n10830 & ~n10835 ) ;
  assign n10837 = ( x82 & n10477 ) | ( x82 & ~n10724 ) | ( n10477 & ~n10724 ) ;
  assign n10838 = x82 & n10477 ;
  assign n10839 = ( ~n10482 & n10837 ) | ( ~n10482 & n10838 ) | ( n10837 & n10838 ) ;
  assign n10840 = ( n10482 & n10837 ) | ( n10482 & n10838 ) | ( n10837 & n10838 ) ;
  assign n10841 = ( n10482 & n10839 ) | ( n10482 & ~n10840 ) | ( n10839 & ~n10840 ) ;
  assign n10842 = ( x83 & n10836 ) | ( x83 & ~n10841 ) | ( n10836 & ~n10841 ) ;
  assign n10843 = ( x83 & n10483 ) | ( x83 & ~n10724 ) | ( n10483 & ~n10724 ) ;
  assign n10844 = x83 & n10483 ;
  assign n10845 = ( ~n10488 & n10843 ) | ( ~n10488 & n10844 ) | ( n10843 & n10844 ) ;
  assign n10846 = ( n10488 & n10843 ) | ( n10488 & n10844 ) | ( n10843 & n10844 ) ;
  assign n10847 = ( n10488 & n10845 ) | ( n10488 & ~n10846 ) | ( n10845 & ~n10846 ) ;
  assign n10848 = ( x84 & n10842 ) | ( x84 & ~n10847 ) | ( n10842 & ~n10847 ) ;
  assign n10849 = ( x84 & n10489 ) | ( x84 & ~n10724 ) | ( n10489 & ~n10724 ) ;
  assign n10850 = x84 & n10489 ;
  assign n10851 = ( ~n10494 & n10849 ) | ( ~n10494 & n10850 ) | ( n10849 & n10850 ) ;
  assign n10852 = ( n10494 & n10849 ) | ( n10494 & n10850 ) | ( n10849 & n10850 ) ;
  assign n10853 = ( n10494 & n10851 ) | ( n10494 & ~n10852 ) | ( n10851 & ~n10852 ) ;
  assign n10854 = ( x85 & n10848 ) | ( x85 & ~n10853 ) | ( n10848 & ~n10853 ) ;
  assign n10855 = ( x85 & n10495 ) | ( x85 & ~n10724 ) | ( n10495 & ~n10724 ) ;
  assign n10856 = x85 & n10495 ;
  assign n10857 = ( ~n10500 & n10855 ) | ( ~n10500 & n10856 ) | ( n10855 & n10856 ) ;
  assign n10858 = ( n10500 & n10855 ) | ( n10500 & n10856 ) | ( n10855 & n10856 ) ;
  assign n10859 = ( n10500 & n10857 ) | ( n10500 & ~n10858 ) | ( n10857 & ~n10858 ) ;
  assign n10860 = ( x86 & n10854 ) | ( x86 & ~n10859 ) | ( n10854 & ~n10859 ) ;
  assign n10861 = ( x86 & n10501 ) | ( x86 & ~n10724 ) | ( n10501 & ~n10724 ) ;
  assign n10862 = x86 & n10501 ;
  assign n10863 = ( ~n10506 & n10861 ) | ( ~n10506 & n10862 ) | ( n10861 & n10862 ) ;
  assign n10864 = ( n10506 & n10861 ) | ( n10506 & n10862 ) | ( n10861 & n10862 ) ;
  assign n10865 = ( n10506 & n10863 ) | ( n10506 & ~n10864 ) | ( n10863 & ~n10864 ) ;
  assign n10866 = ( x87 & n10860 ) | ( x87 & ~n10865 ) | ( n10860 & ~n10865 ) ;
  assign n10867 = ( x87 & n10507 ) | ( x87 & ~n10724 ) | ( n10507 & ~n10724 ) ;
  assign n10868 = x87 & n10507 ;
  assign n10869 = ( ~n10512 & n10867 ) | ( ~n10512 & n10868 ) | ( n10867 & n10868 ) ;
  assign n10870 = ( n10512 & n10867 ) | ( n10512 & n10868 ) | ( n10867 & n10868 ) ;
  assign n10871 = ( n10512 & n10869 ) | ( n10512 & ~n10870 ) | ( n10869 & ~n10870 ) ;
  assign n10872 = ( x88 & n10866 ) | ( x88 & ~n10871 ) | ( n10866 & ~n10871 ) ;
  assign n10873 = ( x88 & n10513 ) | ( x88 & ~n10724 ) | ( n10513 & ~n10724 ) ;
  assign n10874 = x88 & n10513 ;
  assign n10875 = ( ~n10518 & n10873 ) | ( ~n10518 & n10874 ) | ( n10873 & n10874 ) ;
  assign n10876 = ( n10518 & n10873 ) | ( n10518 & n10874 ) | ( n10873 & n10874 ) ;
  assign n10877 = ( n10518 & n10875 ) | ( n10518 & ~n10876 ) | ( n10875 & ~n10876 ) ;
  assign n10878 = ( x89 & n10872 ) | ( x89 & ~n10877 ) | ( n10872 & ~n10877 ) ;
  assign n10879 = ( x89 & n10519 ) | ( x89 & ~n10724 ) | ( n10519 & ~n10724 ) ;
  assign n10880 = x89 & n10519 ;
  assign n10881 = ( ~n10524 & n10879 ) | ( ~n10524 & n10880 ) | ( n10879 & n10880 ) ;
  assign n10882 = ( n10524 & n10879 ) | ( n10524 & n10880 ) | ( n10879 & n10880 ) ;
  assign n10883 = ( n10524 & n10881 ) | ( n10524 & ~n10882 ) | ( n10881 & ~n10882 ) ;
  assign n10884 = ( x90 & n10878 ) | ( x90 & ~n10883 ) | ( n10878 & ~n10883 ) ;
  assign n10885 = ( x90 & n10525 ) | ( x90 & ~n10724 ) | ( n10525 & ~n10724 ) ;
  assign n10886 = x90 & n10525 ;
  assign n10887 = ( ~n10530 & n10885 ) | ( ~n10530 & n10886 ) | ( n10885 & n10886 ) ;
  assign n10888 = ( n10530 & n10885 ) | ( n10530 & n10886 ) | ( n10885 & n10886 ) ;
  assign n10889 = ( n10530 & n10887 ) | ( n10530 & ~n10888 ) | ( n10887 & ~n10888 ) ;
  assign n10890 = ( x91 & n10884 ) | ( x91 & ~n10889 ) | ( n10884 & ~n10889 ) ;
  assign n10891 = ( x91 & n10531 ) | ( x91 & ~n10724 ) | ( n10531 & ~n10724 ) ;
  assign n10892 = x91 & n10531 ;
  assign n10893 = ( ~n10536 & n10891 ) | ( ~n10536 & n10892 ) | ( n10891 & n10892 ) ;
  assign n10894 = ( n10536 & n10891 ) | ( n10536 & n10892 ) | ( n10891 & n10892 ) ;
  assign n10895 = ( n10536 & n10893 ) | ( n10536 & ~n10894 ) | ( n10893 & ~n10894 ) ;
  assign n10896 = ( x92 & n10890 ) | ( x92 & ~n10895 ) | ( n10890 & ~n10895 ) ;
  assign n10897 = ( x92 & n10537 ) | ( x92 & ~n10724 ) | ( n10537 & ~n10724 ) ;
  assign n10898 = x92 & n10537 ;
  assign n10899 = ( ~n10542 & n10897 ) | ( ~n10542 & n10898 ) | ( n10897 & n10898 ) ;
  assign n10900 = ( n10542 & n10897 ) | ( n10542 & n10898 ) | ( n10897 & n10898 ) ;
  assign n10901 = ( n10542 & n10899 ) | ( n10542 & ~n10900 ) | ( n10899 & ~n10900 ) ;
  assign n10902 = ( x93 & n10896 ) | ( x93 & ~n10901 ) | ( n10896 & ~n10901 ) ;
  assign n10903 = ( x93 & n10543 ) | ( x93 & ~n10724 ) | ( n10543 & ~n10724 ) ;
  assign n10904 = x93 & n10543 ;
  assign n10905 = ( ~n10548 & n10903 ) | ( ~n10548 & n10904 ) | ( n10903 & n10904 ) ;
  assign n10906 = ( n10548 & n10903 ) | ( n10548 & n10904 ) | ( n10903 & n10904 ) ;
  assign n10907 = ( n10548 & n10905 ) | ( n10548 & ~n10906 ) | ( n10905 & ~n10906 ) ;
  assign n10908 = ( x94 & n10902 ) | ( x94 & ~n10907 ) | ( n10902 & ~n10907 ) ;
  assign n10909 = ( x94 & n10549 ) | ( x94 & ~n10724 ) | ( n10549 & ~n10724 ) ;
  assign n10910 = x94 & n10549 ;
  assign n10911 = ( ~n10554 & n10909 ) | ( ~n10554 & n10910 ) | ( n10909 & n10910 ) ;
  assign n10912 = ( n10554 & n10909 ) | ( n10554 & n10910 ) | ( n10909 & n10910 ) ;
  assign n10913 = ( n10554 & n10911 ) | ( n10554 & ~n10912 ) | ( n10911 & ~n10912 ) ;
  assign n10914 = ( x95 & n10908 ) | ( x95 & ~n10913 ) | ( n10908 & ~n10913 ) ;
  assign n10915 = ( x95 & n10555 ) | ( x95 & ~n10724 ) | ( n10555 & ~n10724 ) ;
  assign n10916 = x95 & n10555 ;
  assign n10917 = ( ~n10560 & n10915 ) | ( ~n10560 & n10916 ) | ( n10915 & n10916 ) ;
  assign n10918 = ( n10560 & n10915 ) | ( n10560 & n10916 ) | ( n10915 & n10916 ) ;
  assign n10919 = ( n10560 & n10917 ) | ( n10560 & ~n10918 ) | ( n10917 & ~n10918 ) ;
  assign n10920 = ( x96 & n10914 ) | ( x96 & ~n10919 ) | ( n10914 & ~n10919 ) ;
  assign n10921 = ( x96 & n10561 ) | ( x96 & ~n10724 ) | ( n10561 & ~n10724 ) ;
  assign n10922 = x96 & n10561 ;
  assign n10923 = ( ~n10566 & n10921 ) | ( ~n10566 & n10922 ) | ( n10921 & n10922 ) ;
  assign n10924 = ( n10566 & n10921 ) | ( n10566 & n10922 ) | ( n10921 & n10922 ) ;
  assign n10925 = ( n10566 & n10923 ) | ( n10566 & ~n10924 ) | ( n10923 & ~n10924 ) ;
  assign n10926 = ( x97 & n10920 ) | ( x97 & ~n10925 ) | ( n10920 & ~n10925 ) ;
  assign n10927 = ( x97 & n10567 ) | ( x97 & ~n10724 ) | ( n10567 & ~n10724 ) ;
  assign n10928 = x97 & n10567 ;
  assign n10929 = ( ~n10572 & n10927 ) | ( ~n10572 & n10928 ) | ( n10927 & n10928 ) ;
  assign n10930 = ( n10572 & n10927 ) | ( n10572 & n10928 ) | ( n10927 & n10928 ) ;
  assign n10931 = ( n10572 & n10929 ) | ( n10572 & ~n10930 ) | ( n10929 & ~n10930 ) ;
  assign n10932 = ( x98 & n10926 ) | ( x98 & ~n10931 ) | ( n10926 & ~n10931 ) ;
  assign n10933 = ( x98 & n10573 ) | ( x98 & ~n10724 ) | ( n10573 & ~n10724 ) ;
  assign n10934 = x98 & n10573 ;
  assign n10935 = ( ~n10578 & n10933 ) | ( ~n10578 & n10934 ) | ( n10933 & n10934 ) ;
  assign n10936 = ( n10578 & n10933 ) | ( n10578 & n10934 ) | ( n10933 & n10934 ) ;
  assign n10937 = ( n10578 & n10935 ) | ( n10578 & ~n10936 ) | ( n10935 & ~n10936 ) ;
  assign n10938 = ( x99 & n10932 ) | ( x99 & ~n10937 ) | ( n10932 & ~n10937 ) ;
  assign n10939 = ( x99 & n10579 ) | ( x99 & ~n10724 ) | ( n10579 & ~n10724 ) ;
  assign n10940 = x99 & n10579 ;
  assign n10941 = ( ~n10584 & n10939 ) | ( ~n10584 & n10940 ) | ( n10939 & n10940 ) ;
  assign n10942 = ( n10584 & n10939 ) | ( n10584 & n10940 ) | ( n10939 & n10940 ) ;
  assign n10943 = ( n10584 & n10941 ) | ( n10584 & ~n10942 ) | ( n10941 & ~n10942 ) ;
  assign n10944 = ( x100 & n10938 ) | ( x100 & ~n10943 ) | ( n10938 & ~n10943 ) ;
  assign n10945 = ( x100 & n10585 ) | ( x100 & ~n10724 ) | ( n10585 & ~n10724 ) ;
  assign n10946 = x100 & n10585 ;
  assign n10947 = ( ~n10590 & n10945 ) | ( ~n10590 & n10946 ) | ( n10945 & n10946 ) ;
  assign n10948 = ( n10590 & n10945 ) | ( n10590 & n10946 ) | ( n10945 & n10946 ) ;
  assign n10949 = ( n10590 & n10947 ) | ( n10590 & ~n10948 ) | ( n10947 & ~n10948 ) ;
  assign n10950 = ( x101 & n10944 ) | ( x101 & ~n10949 ) | ( n10944 & ~n10949 ) ;
  assign n10951 = ( x101 & n10591 ) | ( x101 & ~n10724 ) | ( n10591 & ~n10724 ) ;
  assign n10952 = x101 & n10591 ;
  assign n10953 = ( ~n10596 & n10951 ) | ( ~n10596 & n10952 ) | ( n10951 & n10952 ) ;
  assign n10954 = ( n10596 & n10951 ) | ( n10596 & n10952 ) | ( n10951 & n10952 ) ;
  assign n10955 = ( n10596 & n10953 ) | ( n10596 & ~n10954 ) | ( n10953 & ~n10954 ) ;
  assign n10956 = ( x102 & n10950 ) | ( x102 & ~n10955 ) | ( n10950 & ~n10955 ) ;
  assign n10957 = ( x102 & n10597 ) | ( x102 & ~n10724 ) | ( n10597 & ~n10724 ) ;
  assign n10958 = x102 & n10597 ;
  assign n10959 = ( ~n10602 & n10957 ) | ( ~n10602 & n10958 ) | ( n10957 & n10958 ) ;
  assign n10960 = ( n10602 & n10957 ) | ( n10602 & n10958 ) | ( n10957 & n10958 ) ;
  assign n10961 = ( n10602 & n10959 ) | ( n10602 & ~n10960 ) | ( n10959 & ~n10960 ) ;
  assign n10962 = ( x103 & n10956 ) | ( x103 & ~n10961 ) | ( n10956 & ~n10961 ) ;
  assign n10963 = ( x103 & n10603 ) | ( x103 & ~n10724 ) | ( n10603 & ~n10724 ) ;
  assign n10964 = x103 & n10603 ;
  assign n10965 = ( ~n10608 & n10963 ) | ( ~n10608 & n10964 ) | ( n10963 & n10964 ) ;
  assign n10966 = ( n10608 & n10963 ) | ( n10608 & n10964 ) | ( n10963 & n10964 ) ;
  assign n10967 = ( n10608 & n10965 ) | ( n10608 & ~n10966 ) | ( n10965 & ~n10966 ) ;
  assign n10968 = ( x104 & n10962 ) | ( x104 & ~n10967 ) | ( n10962 & ~n10967 ) ;
  assign n10969 = ( x104 & n10609 ) | ( x104 & ~n10724 ) | ( n10609 & ~n10724 ) ;
  assign n10970 = x104 & n10609 ;
  assign n10971 = ( ~n10614 & n10969 ) | ( ~n10614 & n10970 ) | ( n10969 & n10970 ) ;
  assign n10972 = ( n10614 & n10969 ) | ( n10614 & n10970 ) | ( n10969 & n10970 ) ;
  assign n10973 = ( n10614 & n10971 ) | ( n10614 & ~n10972 ) | ( n10971 & ~n10972 ) ;
  assign n10974 = ( x105 & n10968 ) | ( x105 & ~n10973 ) | ( n10968 & ~n10973 ) ;
  assign n10975 = ( x105 & n10615 ) | ( x105 & ~n10724 ) | ( n10615 & ~n10724 ) ;
  assign n10976 = x105 & n10615 ;
  assign n10977 = ( ~n10620 & n10975 ) | ( ~n10620 & n10976 ) | ( n10975 & n10976 ) ;
  assign n10978 = ( n10620 & n10975 ) | ( n10620 & n10976 ) | ( n10975 & n10976 ) ;
  assign n10979 = ( n10620 & n10977 ) | ( n10620 & ~n10978 ) | ( n10977 & ~n10978 ) ;
  assign n10980 = ( x106 & n10974 ) | ( x106 & ~n10979 ) | ( n10974 & ~n10979 ) ;
  assign n10981 = ( x106 & n10621 ) | ( x106 & ~n10724 ) | ( n10621 & ~n10724 ) ;
  assign n10982 = x106 & n10621 ;
  assign n10983 = ( ~n10626 & n10981 ) | ( ~n10626 & n10982 ) | ( n10981 & n10982 ) ;
  assign n10984 = ( n10626 & n10981 ) | ( n10626 & n10982 ) | ( n10981 & n10982 ) ;
  assign n10985 = ( n10626 & n10983 ) | ( n10626 & ~n10984 ) | ( n10983 & ~n10984 ) ;
  assign n10986 = ( x107 & n10980 ) | ( x107 & ~n10985 ) | ( n10980 & ~n10985 ) ;
  assign n10987 = ( x107 & n10627 ) | ( x107 & ~n10724 ) | ( n10627 & ~n10724 ) ;
  assign n10988 = x107 & n10627 ;
  assign n10989 = ( ~n10632 & n10987 ) | ( ~n10632 & n10988 ) | ( n10987 & n10988 ) ;
  assign n10990 = ( n10632 & n10987 ) | ( n10632 & n10988 ) | ( n10987 & n10988 ) ;
  assign n10991 = ( n10632 & n10989 ) | ( n10632 & ~n10990 ) | ( n10989 & ~n10990 ) ;
  assign n10992 = ( x108 & n10986 ) | ( x108 & ~n10991 ) | ( n10986 & ~n10991 ) ;
  assign n10993 = ( x108 & n10633 ) | ( x108 & ~n10724 ) | ( n10633 & ~n10724 ) ;
  assign n10994 = x108 & n10633 ;
  assign n10995 = ( ~n10638 & n10993 ) | ( ~n10638 & n10994 ) | ( n10993 & n10994 ) ;
  assign n10996 = ( n10638 & n10993 ) | ( n10638 & n10994 ) | ( n10993 & n10994 ) ;
  assign n10997 = ( n10638 & n10995 ) | ( n10638 & ~n10996 ) | ( n10995 & ~n10996 ) ;
  assign n10998 = ( x109 & n10992 ) | ( x109 & ~n10997 ) | ( n10992 & ~n10997 ) ;
  assign n10999 = ( x109 & n10639 ) | ( x109 & ~n10724 ) | ( n10639 & ~n10724 ) ;
  assign n11000 = x109 & n10639 ;
  assign n11001 = ( ~n10644 & n10999 ) | ( ~n10644 & n11000 ) | ( n10999 & n11000 ) ;
  assign n11002 = ( n10644 & n10999 ) | ( n10644 & n11000 ) | ( n10999 & n11000 ) ;
  assign n11003 = ( n10644 & n11001 ) | ( n10644 & ~n11002 ) | ( n11001 & ~n11002 ) ;
  assign n11004 = ( x110 & n10998 ) | ( x110 & ~n11003 ) | ( n10998 & ~n11003 ) ;
  assign n11005 = ( x110 & n10645 ) | ( x110 & ~n10724 ) | ( n10645 & ~n10724 ) ;
  assign n11006 = x110 & n10645 ;
  assign n11007 = ( ~n10650 & n11005 ) | ( ~n10650 & n11006 ) | ( n11005 & n11006 ) ;
  assign n11008 = ( n10650 & n11005 ) | ( n10650 & n11006 ) | ( n11005 & n11006 ) ;
  assign n11009 = ( n10650 & n11007 ) | ( n10650 & ~n11008 ) | ( n11007 & ~n11008 ) ;
  assign n11010 = ( x111 & n11004 ) | ( x111 & ~n11009 ) | ( n11004 & ~n11009 ) ;
  assign n11011 = ( x111 & n10651 ) | ( x111 & ~n10724 ) | ( n10651 & ~n10724 ) ;
  assign n11012 = x111 & n10651 ;
  assign n11013 = ( ~n10656 & n11011 ) | ( ~n10656 & n11012 ) | ( n11011 & n11012 ) ;
  assign n11014 = ( n10656 & n11011 ) | ( n10656 & n11012 ) | ( n11011 & n11012 ) ;
  assign n11015 = ( n10656 & n11013 ) | ( n10656 & ~n11014 ) | ( n11013 & ~n11014 ) ;
  assign n11016 = ( x112 & n11010 ) | ( x112 & ~n11015 ) | ( n11010 & ~n11015 ) ;
  assign n11017 = ( x112 & n10657 ) | ( x112 & ~n10724 ) | ( n10657 & ~n10724 ) ;
  assign n11018 = x112 & n10657 ;
  assign n11019 = ( ~n10662 & n11017 ) | ( ~n10662 & n11018 ) | ( n11017 & n11018 ) ;
  assign n11020 = ( n10662 & n11017 ) | ( n10662 & n11018 ) | ( n11017 & n11018 ) ;
  assign n11021 = ( n10662 & n11019 ) | ( n10662 & ~n11020 ) | ( n11019 & ~n11020 ) ;
  assign n11022 = ( x113 & n11016 ) | ( x113 & ~n11021 ) | ( n11016 & ~n11021 ) ;
  assign n11023 = ( x113 & n10663 ) | ( x113 & ~n10724 ) | ( n10663 & ~n10724 ) ;
  assign n11024 = x113 & n10663 ;
  assign n11025 = ( ~n10668 & n11023 ) | ( ~n10668 & n11024 ) | ( n11023 & n11024 ) ;
  assign n11026 = ( n10668 & n11023 ) | ( n10668 & n11024 ) | ( n11023 & n11024 ) ;
  assign n11027 = ( n10668 & n11025 ) | ( n10668 & ~n11026 ) | ( n11025 & ~n11026 ) ;
  assign n11028 = ( x114 & n11022 ) | ( x114 & ~n11027 ) | ( n11022 & ~n11027 ) ;
  assign n11029 = ( x114 & n10669 ) | ( x114 & ~n10724 ) | ( n10669 & ~n10724 ) ;
  assign n11030 = x114 & n10669 ;
  assign n11031 = ( ~n10674 & n11029 ) | ( ~n10674 & n11030 ) | ( n11029 & n11030 ) ;
  assign n11032 = ( n10674 & n11029 ) | ( n10674 & n11030 ) | ( n11029 & n11030 ) ;
  assign n11033 = ( n10674 & n11031 ) | ( n10674 & ~n11032 ) | ( n11031 & ~n11032 ) ;
  assign n11034 = ( x115 & n11028 ) | ( x115 & ~n11033 ) | ( n11028 & ~n11033 ) ;
  assign n11035 = ( x115 & n10675 ) | ( x115 & ~n10724 ) | ( n10675 & ~n10724 ) ;
  assign n11036 = x115 & n10675 ;
  assign n11037 = ( ~n10680 & n11035 ) | ( ~n10680 & n11036 ) | ( n11035 & n11036 ) ;
  assign n11038 = ( n10680 & n11035 ) | ( n10680 & n11036 ) | ( n11035 & n11036 ) ;
  assign n11039 = ( n10680 & n11037 ) | ( n10680 & ~n11038 ) | ( n11037 & ~n11038 ) ;
  assign n11040 = ( x116 & n11034 ) | ( x116 & ~n11039 ) | ( n11034 & ~n11039 ) ;
  assign n11041 = ( x116 & n10681 ) | ( x116 & ~n10724 ) | ( n10681 & ~n10724 ) ;
  assign n11042 = x116 & n10681 ;
  assign n11043 = ( ~n10686 & n11041 ) | ( ~n10686 & n11042 ) | ( n11041 & n11042 ) ;
  assign n11044 = ( n10686 & n11041 ) | ( n10686 & n11042 ) | ( n11041 & n11042 ) ;
  assign n11045 = ( n10686 & n11043 ) | ( n10686 & ~n11044 ) | ( n11043 & ~n11044 ) ;
  assign n11046 = ( x117 & n11040 ) | ( x117 & ~n11045 ) | ( n11040 & ~n11045 ) ;
  assign n11047 = ( x117 & n10687 ) | ( x117 & ~n10724 ) | ( n10687 & ~n10724 ) ;
  assign n11048 = x117 & n10687 ;
  assign n11049 = ( ~n10692 & n11047 ) | ( ~n10692 & n11048 ) | ( n11047 & n11048 ) ;
  assign n11050 = ( n10692 & n11047 ) | ( n10692 & n11048 ) | ( n11047 & n11048 ) ;
  assign n11051 = ( n10692 & n11049 ) | ( n10692 & ~n11050 ) | ( n11049 & ~n11050 ) ;
  assign n11052 = ( x118 & n11046 ) | ( x118 & ~n11051 ) | ( n11046 & ~n11051 ) ;
  assign n11053 = ( x118 & n10693 ) | ( x118 & ~n10724 ) | ( n10693 & ~n10724 ) ;
  assign n11054 = x118 & n10693 ;
  assign n11055 = ( ~n10698 & n11053 ) | ( ~n10698 & n11054 ) | ( n11053 & n11054 ) ;
  assign n11056 = ( n10698 & n11053 ) | ( n10698 & n11054 ) | ( n11053 & n11054 ) ;
  assign n11057 = ( n10698 & n11055 ) | ( n10698 & ~n11056 ) | ( n11055 & ~n11056 ) ;
  assign n11058 = ( x119 & n11052 ) | ( x119 & ~n11057 ) | ( n11052 & ~n11057 ) ;
  assign n11059 = ( x119 & n10699 ) | ( x119 & ~n10724 ) | ( n10699 & ~n10724 ) ;
  assign n11060 = x119 & n10699 ;
  assign n11061 = ( ~n10704 & n11059 ) | ( ~n10704 & n11060 ) | ( n11059 & n11060 ) ;
  assign n11062 = ( n10704 & n11059 ) | ( n10704 & n11060 ) | ( n11059 & n11060 ) ;
  assign n11063 = ( n10704 & n11061 ) | ( n10704 & ~n11062 ) | ( n11061 & ~n11062 ) ;
  assign n11064 = ( x120 & n11058 ) | ( x120 & ~n11063 ) | ( n11058 & ~n11063 ) ;
  assign n11065 = ( x120 & n10705 ) | ( x120 & ~n10724 ) | ( n10705 & ~n10724 ) ;
  assign n11066 = x120 & n10705 ;
  assign n11067 = ( ~n10710 & n11065 ) | ( ~n10710 & n11066 ) | ( n11065 & n11066 ) ;
  assign n11068 = ( n10710 & n11065 ) | ( n10710 & n11066 ) | ( n11065 & n11066 ) ;
  assign n11069 = ( n10710 & n11067 ) | ( n10710 & ~n11068 ) | ( n11067 & ~n11068 ) ;
  assign n11070 = ( x121 & n11064 ) | ( x121 & ~n11069 ) | ( n11064 & ~n11069 ) ;
  assign n11071 = ( x121 & n10711 ) | ( x121 & ~n10724 ) | ( n10711 & ~n10724 ) ;
  assign n11072 = x121 & n10711 ;
  assign n11073 = ( ~n10716 & n11071 ) | ( ~n10716 & n11072 ) | ( n11071 & n11072 ) ;
  assign n11074 = ( n10716 & n11071 ) | ( n10716 & n11072 ) | ( n11071 & n11072 ) ;
  assign n11075 = ( n10716 & n11073 ) | ( n10716 & ~n11074 ) | ( n11073 & ~n11074 ) ;
  assign n11076 = ( x122 & n11070 ) | ( x122 & ~n11075 ) | ( n11070 & ~n11075 ) ;
  assign n11077 = ( x123 & ~n10729 ) | ( x123 & n11076 ) | ( ~n10729 & n11076 ) ;
  assign n11078 = n132 | n11077 ;
  assign n11079 = ( ~x123 & n133 ) | ( ~x123 & n10722 ) | ( n133 & n10722 ) ;
  assign n11080 = ( ~x123 & n10721 ) | ( ~x123 & n10722 ) | ( n10721 & n10722 ) ;
  assign n11081 = ~n11079 & n11080 ;
  assign n11082 = x124 & ~n10721 ;
  assign n11083 = ( n11078 & ~n11081 ) | ( n11078 & n11082 ) | ( ~n11081 & n11082 ) ;
  assign n11084 = x3 & n11083 ;
  assign n11085 = ( x3 & x64 ) | ( x3 & ~n11083 ) | ( x64 & ~n11083 ) ;
  assign n11086 = x3 & x64 ;
  assign n11087 = ( n11084 & n11085 ) | ( n11084 & ~n11086 ) | ( n11085 & ~n11086 ) ;
  assign n11088 = ( x65 & n391 ) | ( x65 & ~n11087 ) | ( n391 & ~n11087 ) ;
  assign n11089 = ( x65 & n10730 ) | ( x65 & n11083 ) | ( n10730 & n11083 ) ;
  assign n11090 = x65 | n10730 ;
  assign n11091 = ( ~n10733 & n11089 ) | ( ~n10733 & n11090 ) | ( n11089 & n11090 ) ;
  assign n11092 = ( n10733 & n11089 ) | ( n10733 & n11090 ) | ( n11089 & n11090 ) ;
  assign n11093 = ( n10733 & n11091 ) | ( n10733 & ~n11092 ) | ( n11091 & ~n11092 ) ;
  assign n11094 = ( x66 & n11088 ) | ( x66 & ~n11093 ) | ( n11088 & ~n11093 ) ;
  assign n11095 = ( x66 & n10734 ) | ( x66 & n11083 ) | ( n10734 & n11083 ) ;
  assign n11096 = x66 | n10734 ;
  assign n11097 = ( ~n10739 & n11095 ) | ( ~n10739 & n11096 ) | ( n11095 & n11096 ) ;
  assign n11098 = ( n10739 & n11095 ) | ( n10739 & n11096 ) | ( n11095 & n11096 ) ;
  assign n11099 = ( n10739 & n11097 ) | ( n10739 & ~n11098 ) | ( n11097 & ~n11098 ) ;
  assign n11100 = ( x67 & n11094 ) | ( x67 & ~n11099 ) | ( n11094 & ~n11099 ) ;
  assign n11101 = ( x67 & n10740 ) | ( x67 & ~n11083 ) | ( n10740 & ~n11083 ) ;
  assign n11102 = x67 & n10740 ;
  assign n11103 = ( ~n10745 & n11101 ) | ( ~n10745 & n11102 ) | ( n11101 & n11102 ) ;
  assign n11104 = ( n10745 & n11101 ) | ( n10745 & n11102 ) | ( n11101 & n11102 ) ;
  assign n11105 = ( n10745 & n11103 ) | ( n10745 & ~n11104 ) | ( n11103 & ~n11104 ) ;
  assign n11106 = ( x68 & n11100 ) | ( x68 & ~n11105 ) | ( n11100 & ~n11105 ) ;
  assign n11107 = ( x68 & n10746 ) | ( x68 & ~n11083 ) | ( n10746 & ~n11083 ) ;
  assign n11108 = x68 & n10746 ;
  assign n11109 = ( ~n10751 & n11107 ) | ( ~n10751 & n11108 ) | ( n11107 & n11108 ) ;
  assign n11110 = ( n10751 & n11107 ) | ( n10751 & n11108 ) | ( n11107 & n11108 ) ;
  assign n11111 = ( n10751 & n11109 ) | ( n10751 & ~n11110 ) | ( n11109 & ~n11110 ) ;
  assign n11112 = ( x69 & n11106 ) | ( x69 & ~n11111 ) | ( n11106 & ~n11111 ) ;
  assign n11113 = ( x69 & n10752 ) | ( x69 & ~n11083 ) | ( n10752 & ~n11083 ) ;
  assign n11114 = x69 & n10752 ;
  assign n11115 = ( ~n10757 & n11113 ) | ( ~n10757 & n11114 ) | ( n11113 & n11114 ) ;
  assign n11116 = ( n10757 & n11113 ) | ( n10757 & n11114 ) | ( n11113 & n11114 ) ;
  assign n11117 = ( n10757 & n11115 ) | ( n10757 & ~n11116 ) | ( n11115 & ~n11116 ) ;
  assign n11118 = ( x70 & n11112 ) | ( x70 & ~n11117 ) | ( n11112 & ~n11117 ) ;
  assign n11119 = ( x70 & n10758 ) | ( x70 & ~n11083 ) | ( n10758 & ~n11083 ) ;
  assign n11120 = x70 & n10758 ;
  assign n11121 = ( ~n10763 & n11119 ) | ( ~n10763 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11122 = ( n10763 & n11119 ) | ( n10763 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11123 = ( n10763 & n11121 ) | ( n10763 & ~n11122 ) | ( n11121 & ~n11122 ) ;
  assign n11124 = ( x71 & n11118 ) | ( x71 & ~n11123 ) | ( n11118 & ~n11123 ) ;
  assign n11125 = ( x71 & n10764 ) | ( x71 & ~n11083 ) | ( n10764 & ~n11083 ) ;
  assign n11126 = x71 & n10764 ;
  assign n11127 = ( ~n10769 & n11125 ) | ( ~n10769 & n11126 ) | ( n11125 & n11126 ) ;
  assign n11128 = ( n10769 & n11125 ) | ( n10769 & n11126 ) | ( n11125 & n11126 ) ;
  assign n11129 = ( n10769 & n11127 ) | ( n10769 & ~n11128 ) | ( n11127 & ~n11128 ) ;
  assign n11130 = ( x72 & n11124 ) | ( x72 & ~n11129 ) | ( n11124 & ~n11129 ) ;
  assign n11131 = ( x72 & n10770 ) | ( x72 & ~n11083 ) | ( n10770 & ~n11083 ) ;
  assign n11132 = x72 & n10770 ;
  assign n11133 = ( ~n10775 & n11131 ) | ( ~n10775 & n11132 ) | ( n11131 & n11132 ) ;
  assign n11134 = ( n10775 & n11131 ) | ( n10775 & n11132 ) | ( n11131 & n11132 ) ;
  assign n11135 = ( n10775 & n11133 ) | ( n10775 & ~n11134 ) | ( n11133 & ~n11134 ) ;
  assign n11136 = ( x73 & n11130 ) | ( x73 & ~n11135 ) | ( n11130 & ~n11135 ) ;
  assign n11137 = ( x73 & n10776 ) | ( x73 & ~n11083 ) | ( n10776 & ~n11083 ) ;
  assign n11138 = x73 & n10776 ;
  assign n11139 = ( ~n10781 & n11137 ) | ( ~n10781 & n11138 ) | ( n11137 & n11138 ) ;
  assign n11140 = ( n10781 & n11137 ) | ( n10781 & n11138 ) | ( n11137 & n11138 ) ;
  assign n11141 = ( n10781 & n11139 ) | ( n10781 & ~n11140 ) | ( n11139 & ~n11140 ) ;
  assign n11142 = ( x74 & n11136 ) | ( x74 & ~n11141 ) | ( n11136 & ~n11141 ) ;
  assign n11143 = ( x74 & n10782 ) | ( x74 & ~n11083 ) | ( n10782 & ~n11083 ) ;
  assign n11144 = x74 & n10782 ;
  assign n11145 = ( ~n10787 & n11143 ) | ( ~n10787 & n11144 ) | ( n11143 & n11144 ) ;
  assign n11146 = ( n10787 & n11143 ) | ( n10787 & n11144 ) | ( n11143 & n11144 ) ;
  assign n11147 = ( n10787 & n11145 ) | ( n10787 & ~n11146 ) | ( n11145 & ~n11146 ) ;
  assign n11148 = ( x75 & n11142 ) | ( x75 & ~n11147 ) | ( n11142 & ~n11147 ) ;
  assign n11149 = ( x75 & n10788 ) | ( x75 & ~n11083 ) | ( n10788 & ~n11083 ) ;
  assign n11150 = x75 & n10788 ;
  assign n11151 = ( ~n10793 & n11149 ) | ( ~n10793 & n11150 ) | ( n11149 & n11150 ) ;
  assign n11152 = ( n10793 & n11149 ) | ( n10793 & n11150 ) | ( n11149 & n11150 ) ;
  assign n11153 = ( n10793 & n11151 ) | ( n10793 & ~n11152 ) | ( n11151 & ~n11152 ) ;
  assign n11154 = ( x76 & n11148 ) | ( x76 & ~n11153 ) | ( n11148 & ~n11153 ) ;
  assign n11155 = ( x76 & n10794 ) | ( x76 & ~n11083 ) | ( n10794 & ~n11083 ) ;
  assign n11156 = x76 & n10794 ;
  assign n11157 = ( ~n10799 & n11155 ) | ( ~n10799 & n11156 ) | ( n11155 & n11156 ) ;
  assign n11158 = ( n10799 & n11155 ) | ( n10799 & n11156 ) | ( n11155 & n11156 ) ;
  assign n11159 = ( n10799 & n11157 ) | ( n10799 & ~n11158 ) | ( n11157 & ~n11158 ) ;
  assign n11160 = ( x77 & n11154 ) | ( x77 & ~n11159 ) | ( n11154 & ~n11159 ) ;
  assign n11161 = ( x77 & n10800 ) | ( x77 & ~n11083 ) | ( n10800 & ~n11083 ) ;
  assign n11162 = x77 & n10800 ;
  assign n11163 = ( ~n10805 & n11161 ) | ( ~n10805 & n11162 ) | ( n11161 & n11162 ) ;
  assign n11164 = ( n10805 & n11161 ) | ( n10805 & n11162 ) | ( n11161 & n11162 ) ;
  assign n11165 = ( n10805 & n11163 ) | ( n10805 & ~n11164 ) | ( n11163 & ~n11164 ) ;
  assign n11166 = ( x78 & n11160 ) | ( x78 & ~n11165 ) | ( n11160 & ~n11165 ) ;
  assign n11167 = ( x78 & n10806 ) | ( x78 & ~n11083 ) | ( n10806 & ~n11083 ) ;
  assign n11168 = x78 & n10806 ;
  assign n11169 = ( ~n10811 & n11167 ) | ( ~n10811 & n11168 ) | ( n11167 & n11168 ) ;
  assign n11170 = ( n10811 & n11167 ) | ( n10811 & n11168 ) | ( n11167 & n11168 ) ;
  assign n11171 = ( n10811 & n11169 ) | ( n10811 & ~n11170 ) | ( n11169 & ~n11170 ) ;
  assign n11172 = ( x79 & n11166 ) | ( x79 & ~n11171 ) | ( n11166 & ~n11171 ) ;
  assign n11173 = ( x79 & n10812 ) | ( x79 & ~n11083 ) | ( n10812 & ~n11083 ) ;
  assign n11174 = x79 & n10812 ;
  assign n11175 = ( ~n10817 & n11173 ) | ( ~n10817 & n11174 ) | ( n11173 & n11174 ) ;
  assign n11176 = ( n10817 & n11173 ) | ( n10817 & n11174 ) | ( n11173 & n11174 ) ;
  assign n11177 = ( n10817 & n11175 ) | ( n10817 & ~n11176 ) | ( n11175 & ~n11176 ) ;
  assign n11178 = ( x80 & n11172 ) | ( x80 & ~n11177 ) | ( n11172 & ~n11177 ) ;
  assign n11179 = ( x80 & n10818 ) | ( x80 & ~n11083 ) | ( n10818 & ~n11083 ) ;
  assign n11180 = x80 & n10818 ;
  assign n11181 = ( ~n10823 & n11179 ) | ( ~n10823 & n11180 ) | ( n11179 & n11180 ) ;
  assign n11182 = ( n10823 & n11179 ) | ( n10823 & n11180 ) | ( n11179 & n11180 ) ;
  assign n11183 = ( n10823 & n11181 ) | ( n10823 & ~n11182 ) | ( n11181 & ~n11182 ) ;
  assign n11184 = ( x81 & n11178 ) | ( x81 & ~n11183 ) | ( n11178 & ~n11183 ) ;
  assign n11185 = ( x81 & n10824 ) | ( x81 & ~n11083 ) | ( n10824 & ~n11083 ) ;
  assign n11186 = x81 & n10824 ;
  assign n11187 = ( ~n10829 & n11185 ) | ( ~n10829 & n11186 ) | ( n11185 & n11186 ) ;
  assign n11188 = ( n10829 & n11185 ) | ( n10829 & n11186 ) | ( n11185 & n11186 ) ;
  assign n11189 = ( n10829 & n11187 ) | ( n10829 & ~n11188 ) | ( n11187 & ~n11188 ) ;
  assign n11190 = ( x82 & n11184 ) | ( x82 & ~n11189 ) | ( n11184 & ~n11189 ) ;
  assign n11191 = ( x82 & n10830 ) | ( x82 & ~n11083 ) | ( n10830 & ~n11083 ) ;
  assign n11192 = x82 & n10830 ;
  assign n11193 = ( ~n10835 & n11191 ) | ( ~n10835 & n11192 ) | ( n11191 & n11192 ) ;
  assign n11194 = ( n10835 & n11191 ) | ( n10835 & n11192 ) | ( n11191 & n11192 ) ;
  assign n11195 = ( n10835 & n11193 ) | ( n10835 & ~n11194 ) | ( n11193 & ~n11194 ) ;
  assign n11196 = ( x83 & n11190 ) | ( x83 & ~n11195 ) | ( n11190 & ~n11195 ) ;
  assign n11197 = ( x83 & n10836 ) | ( x83 & ~n11083 ) | ( n10836 & ~n11083 ) ;
  assign n11198 = x83 & n10836 ;
  assign n11199 = ( ~n10841 & n11197 ) | ( ~n10841 & n11198 ) | ( n11197 & n11198 ) ;
  assign n11200 = ( n10841 & n11197 ) | ( n10841 & n11198 ) | ( n11197 & n11198 ) ;
  assign n11201 = ( n10841 & n11199 ) | ( n10841 & ~n11200 ) | ( n11199 & ~n11200 ) ;
  assign n11202 = ( x84 & n11196 ) | ( x84 & ~n11201 ) | ( n11196 & ~n11201 ) ;
  assign n11203 = ( x84 & n10842 ) | ( x84 & ~n11083 ) | ( n10842 & ~n11083 ) ;
  assign n11204 = x84 & n10842 ;
  assign n11205 = ( ~n10847 & n11203 ) | ( ~n10847 & n11204 ) | ( n11203 & n11204 ) ;
  assign n11206 = ( n10847 & n11203 ) | ( n10847 & n11204 ) | ( n11203 & n11204 ) ;
  assign n11207 = ( n10847 & n11205 ) | ( n10847 & ~n11206 ) | ( n11205 & ~n11206 ) ;
  assign n11208 = ( x85 & n11202 ) | ( x85 & ~n11207 ) | ( n11202 & ~n11207 ) ;
  assign n11209 = ( x85 & n10848 ) | ( x85 & ~n11083 ) | ( n10848 & ~n11083 ) ;
  assign n11210 = x85 & n10848 ;
  assign n11211 = ( ~n10853 & n11209 ) | ( ~n10853 & n11210 ) | ( n11209 & n11210 ) ;
  assign n11212 = ( n10853 & n11209 ) | ( n10853 & n11210 ) | ( n11209 & n11210 ) ;
  assign n11213 = ( n10853 & n11211 ) | ( n10853 & ~n11212 ) | ( n11211 & ~n11212 ) ;
  assign n11214 = ( x86 & n11208 ) | ( x86 & ~n11213 ) | ( n11208 & ~n11213 ) ;
  assign n11215 = ( x86 & n10854 ) | ( x86 & ~n11083 ) | ( n10854 & ~n11083 ) ;
  assign n11216 = x86 & n10854 ;
  assign n11217 = ( ~n10859 & n11215 ) | ( ~n10859 & n11216 ) | ( n11215 & n11216 ) ;
  assign n11218 = ( n10859 & n11215 ) | ( n10859 & n11216 ) | ( n11215 & n11216 ) ;
  assign n11219 = ( n10859 & n11217 ) | ( n10859 & ~n11218 ) | ( n11217 & ~n11218 ) ;
  assign n11220 = ( x87 & n11214 ) | ( x87 & ~n11219 ) | ( n11214 & ~n11219 ) ;
  assign n11221 = ( x87 & n10860 ) | ( x87 & ~n11083 ) | ( n10860 & ~n11083 ) ;
  assign n11222 = x87 & n10860 ;
  assign n11223 = ( ~n10865 & n11221 ) | ( ~n10865 & n11222 ) | ( n11221 & n11222 ) ;
  assign n11224 = ( n10865 & n11221 ) | ( n10865 & n11222 ) | ( n11221 & n11222 ) ;
  assign n11225 = ( n10865 & n11223 ) | ( n10865 & ~n11224 ) | ( n11223 & ~n11224 ) ;
  assign n11226 = ( x88 & n11220 ) | ( x88 & ~n11225 ) | ( n11220 & ~n11225 ) ;
  assign n11227 = ( x88 & n10866 ) | ( x88 & ~n11083 ) | ( n10866 & ~n11083 ) ;
  assign n11228 = x88 & n10866 ;
  assign n11229 = ( ~n10871 & n11227 ) | ( ~n10871 & n11228 ) | ( n11227 & n11228 ) ;
  assign n11230 = ( n10871 & n11227 ) | ( n10871 & n11228 ) | ( n11227 & n11228 ) ;
  assign n11231 = ( n10871 & n11229 ) | ( n10871 & ~n11230 ) | ( n11229 & ~n11230 ) ;
  assign n11232 = ( x89 & n11226 ) | ( x89 & ~n11231 ) | ( n11226 & ~n11231 ) ;
  assign n11233 = ( x89 & n10872 ) | ( x89 & ~n11083 ) | ( n10872 & ~n11083 ) ;
  assign n11234 = x89 & n10872 ;
  assign n11235 = ( ~n10877 & n11233 ) | ( ~n10877 & n11234 ) | ( n11233 & n11234 ) ;
  assign n11236 = ( n10877 & n11233 ) | ( n10877 & n11234 ) | ( n11233 & n11234 ) ;
  assign n11237 = ( n10877 & n11235 ) | ( n10877 & ~n11236 ) | ( n11235 & ~n11236 ) ;
  assign n11238 = ( x90 & n11232 ) | ( x90 & ~n11237 ) | ( n11232 & ~n11237 ) ;
  assign n11239 = ( x90 & n10878 ) | ( x90 & ~n11083 ) | ( n10878 & ~n11083 ) ;
  assign n11240 = x90 & n10878 ;
  assign n11241 = ( ~n10883 & n11239 ) | ( ~n10883 & n11240 ) | ( n11239 & n11240 ) ;
  assign n11242 = ( n10883 & n11239 ) | ( n10883 & n11240 ) | ( n11239 & n11240 ) ;
  assign n11243 = ( n10883 & n11241 ) | ( n10883 & ~n11242 ) | ( n11241 & ~n11242 ) ;
  assign n11244 = ( x91 & n11238 ) | ( x91 & ~n11243 ) | ( n11238 & ~n11243 ) ;
  assign n11245 = ( x91 & n10884 ) | ( x91 & ~n11083 ) | ( n10884 & ~n11083 ) ;
  assign n11246 = x91 & n10884 ;
  assign n11247 = ( ~n10889 & n11245 ) | ( ~n10889 & n11246 ) | ( n11245 & n11246 ) ;
  assign n11248 = ( n10889 & n11245 ) | ( n10889 & n11246 ) | ( n11245 & n11246 ) ;
  assign n11249 = ( n10889 & n11247 ) | ( n10889 & ~n11248 ) | ( n11247 & ~n11248 ) ;
  assign n11250 = ( x92 & n11244 ) | ( x92 & ~n11249 ) | ( n11244 & ~n11249 ) ;
  assign n11251 = ( x92 & n10890 ) | ( x92 & ~n11083 ) | ( n10890 & ~n11083 ) ;
  assign n11252 = x92 & n10890 ;
  assign n11253 = ( ~n10895 & n11251 ) | ( ~n10895 & n11252 ) | ( n11251 & n11252 ) ;
  assign n11254 = ( n10895 & n11251 ) | ( n10895 & n11252 ) | ( n11251 & n11252 ) ;
  assign n11255 = ( n10895 & n11253 ) | ( n10895 & ~n11254 ) | ( n11253 & ~n11254 ) ;
  assign n11256 = ( x93 & n11250 ) | ( x93 & ~n11255 ) | ( n11250 & ~n11255 ) ;
  assign n11257 = ( x93 & n10896 ) | ( x93 & ~n11083 ) | ( n10896 & ~n11083 ) ;
  assign n11258 = x93 & n10896 ;
  assign n11259 = ( ~n10901 & n11257 ) | ( ~n10901 & n11258 ) | ( n11257 & n11258 ) ;
  assign n11260 = ( n10901 & n11257 ) | ( n10901 & n11258 ) | ( n11257 & n11258 ) ;
  assign n11261 = ( n10901 & n11259 ) | ( n10901 & ~n11260 ) | ( n11259 & ~n11260 ) ;
  assign n11262 = ( x94 & n11256 ) | ( x94 & ~n11261 ) | ( n11256 & ~n11261 ) ;
  assign n11263 = ( x94 & n10902 ) | ( x94 & ~n11083 ) | ( n10902 & ~n11083 ) ;
  assign n11264 = x94 & n10902 ;
  assign n11265 = ( ~n10907 & n11263 ) | ( ~n10907 & n11264 ) | ( n11263 & n11264 ) ;
  assign n11266 = ( n10907 & n11263 ) | ( n10907 & n11264 ) | ( n11263 & n11264 ) ;
  assign n11267 = ( n10907 & n11265 ) | ( n10907 & ~n11266 ) | ( n11265 & ~n11266 ) ;
  assign n11268 = ( x95 & n11262 ) | ( x95 & ~n11267 ) | ( n11262 & ~n11267 ) ;
  assign n11269 = ( x95 & n10908 ) | ( x95 & ~n11083 ) | ( n10908 & ~n11083 ) ;
  assign n11270 = x95 & n10908 ;
  assign n11271 = ( ~n10913 & n11269 ) | ( ~n10913 & n11270 ) | ( n11269 & n11270 ) ;
  assign n11272 = ( n10913 & n11269 ) | ( n10913 & n11270 ) | ( n11269 & n11270 ) ;
  assign n11273 = ( n10913 & n11271 ) | ( n10913 & ~n11272 ) | ( n11271 & ~n11272 ) ;
  assign n11274 = ( x96 & n11268 ) | ( x96 & ~n11273 ) | ( n11268 & ~n11273 ) ;
  assign n11275 = ( x96 & n10914 ) | ( x96 & ~n11083 ) | ( n10914 & ~n11083 ) ;
  assign n11276 = x96 & n10914 ;
  assign n11277 = ( ~n10919 & n11275 ) | ( ~n10919 & n11276 ) | ( n11275 & n11276 ) ;
  assign n11278 = ( n10919 & n11275 ) | ( n10919 & n11276 ) | ( n11275 & n11276 ) ;
  assign n11279 = ( n10919 & n11277 ) | ( n10919 & ~n11278 ) | ( n11277 & ~n11278 ) ;
  assign n11280 = ( x97 & n11274 ) | ( x97 & ~n11279 ) | ( n11274 & ~n11279 ) ;
  assign n11281 = ( x97 & n10920 ) | ( x97 & ~n11083 ) | ( n10920 & ~n11083 ) ;
  assign n11282 = x97 & n10920 ;
  assign n11283 = ( ~n10925 & n11281 ) | ( ~n10925 & n11282 ) | ( n11281 & n11282 ) ;
  assign n11284 = ( n10925 & n11281 ) | ( n10925 & n11282 ) | ( n11281 & n11282 ) ;
  assign n11285 = ( n10925 & n11283 ) | ( n10925 & ~n11284 ) | ( n11283 & ~n11284 ) ;
  assign n11286 = ( x98 & n11280 ) | ( x98 & ~n11285 ) | ( n11280 & ~n11285 ) ;
  assign n11287 = ( x98 & n10926 ) | ( x98 & ~n11083 ) | ( n10926 & ~n11083 ) ;
  assign n11288 = x98 & n10926 ;
  assign n11289 = ( ~n10931 & n11287 ) | ( ~n10931 & n11288 ) | ( n11287 & n11288 ) ;
  assign n11290 = ( n10931 & n11287 ) | ( n10931 & n11288 ) | ( n11287 & n11288 ) ;
  assign n11291 = ( n10931 & n11289 ) | ( n10931 & ~n11290 ) | ( n11289 & ~n11290 ) ;
  assign n11292 = ( x99 & n11286 ) | ( x99 & ~n11291 ) | ( n11286 & ~n11291 ) ;
  assign n11293 = ( x99 & n10932 ) | ( x99 & ~n11083 ) | ( n10932 & ~n11083 ) ;
  assign n11294 = x99 & n10932 ;
  assign n11295 = ( ~n10937 & n11293 ) | ( ~n10937 & n11294 ) | ( n11293 & n11294 ) ;
  assign n11296 = ( n10937 & n11293 ) | ( n10937 & n11294 ) | ( n11293 & n11294 ) ;
  assign n11297 = ( n10937 & n11295 ) | ( n10937 & ~n11296 ) | ( n11295 & ~n11296 ) ;
  assign n11298 = ( x100 & n11292 ) | ( x100 & ~n11297 ) | ( n11292 & ~n11297 ) ;
  assign n11299 = ( x100 & n10938 ) | ( x100 & ~n11083 ) | ( n10938 & ~n11083 ) ;
  assign n11300 = x100 & n10938 ;
  assign n11301 = ( ~n10943 & n11299 ) | ( ~n10943 & n11300 ) | ( n11299 & n11300 ) ;
  assign n11302 = ( n10943 & n11299 ) | ( n10943 & n11300 ) | ( n11299 & n11300 ) ;
  assign n11303 = ( n10943 & n11301 ) | ( n10943 & ~n11302 ) | ( n11301 & ~n11302 ) ;
  assign n11304 = ( x101 & n11298 ) | ( x101 & ~n11303 ) | ( n11298 & ~n11303 ) ;
  assign n11305 = ( x101 & n10944 ) | ( x101 & ~n11083 ) | ( n10944 & ~n11083 ) ;
  assign n11306 = x101 & n10944 ;
  assign n11307 = ( ~n10949 & n11305 ) | ( ~n10949 & n11306 ) | ( n11305 & n11306 ) ;
  assign n11308 = ( n10949 & n11305 ) | ( n10949 & n11306 ) | ( n11305 & n11306 ) ;
  assign n11309 = ( n10949 & n11307 ) | ( n10949 & ~n11308 ) | ( n11307 & ~n11308 ) ;
  assign n11310 = ( x102 & n11304 ) | ( x102 & ~n11309 ) | ( n11304 & ~n11309 ) ;
  assign n11311 = ( x102 & n10950 ) | ( x102 & ~n11083 ) | ( n10950 & ~n11083 ) ;
  assign n11312 = x102 & n10950 ;
  assign n11313 = ( ~n10955 & n11311 ) | ( ~n10955 & n11312 ) | ( n11311 & n11312 ) ;
  assign n11314 = ( n10955 & n11311 ) | ( n10955 & n11312 ) | ( n11311 & n11312 ) ;
  assign n11315 = ( n10955 & n11313 ) | ( n10955 & ~n11314 ) | ( n11313 & ~n11314 ) ;
  assign n11316 = ( x103 & n11310 ) | ( x103 & ~n11315 ) | ( n11310 & ~n11315 ) ;
  assign n11317 = ( x103 & n10956 ) | ( x103 & ~n11083 ) | ( n10956 & ~n11083 ) ;
  assign n11318 = x103 & n10956 ;
  assign n11319 = ( ~n10961 & n11317 ) | ( ~n10961 & n11318 ) | ( n11317 & n11318 ) ;
  assign n11320 = ( n10961 & n11317 ) | ( n10961 & n11318 ) | ( n11317 & n11318 ) ;
  assign n11321 = ( n10961 & n11319 ) | ( n10961 & ~n11320 ) | ( n11319 & ~n11320 ) ;
  assign n11322 = ( x104 & n11316 ) | ( x104 & ~n11321 ) | ( n11316 & ~n11321 ) ;
  assign n11323 = ( x104 & n10962 ) | ( x104 & ~n11083 ) | ( n10962 & ~n11083 ) ;
  assign n11324 = x104 & n10962 ;
  assign n11325 = ( ~n10967 & n11323 ) | ( ~n10967 & n11324 ) | ( n11323 & n11324 ) ;
  assign n11326 = ( n10967 & n11323 ) | ( n10967 & n11324 ) | ( n11323 & n11324 ) ;
  assign n11327 = ( n10967 & n11325 ) | ( n10967 & ~n11326 ) | ( n11325 & ~n11326 ) ;
  assign n11328 = ( x105 & n11322 ) | ( x105 & ~n11327 ) | ( n11322 & ~n11327 ) ;
  assign n11329 = ( x105 & n10968 ) | ( x105 & ~n11083 ) | ( n10968 & ~n11083 ) ;
  assign n11330 = x105 & n10968 ;
  assign n11331 = ( ~n10973 & n11329 ) | ( ~n10973 & n11330 ) | ( n11329 & n11330 ) ;
  assign n11332 = ( n10973 & n11329 ) | ( n10973 & n11330 ) | ( n11329 & n11330 ) ;
  assign n11333 = ( n10973 & n11331 ) | ( n10973 & ~n11332 ) | ( n11331 & ~n11332 ) ;
  assign n11334 = ( x106 & n11328 ) | ( x106 & ~n11333 ) | ( n11328 & ~n11333 ) ;
  assign n11335 = ( x106 & n10974 ) | ( x106 & ~n11083 ) | ( n10974 & ~n11083 ) ;
  assign n11336 = x106 & n10974 ;
  assign n11337 = ( ~n10979 & n11335 ) | ( ~n10979 & n11336 ) | ( n11335 & n11336 ) ;
  assign n11338 = ( n10979 & n11335 ) | ( n10979 & n11336 ) | ( n11335 & n11336 ) ;
  assign n11339 = ( n10979 & n11337 ) | ( n10979 & ~n11338 ) | ( n11337 & ~n11338 ) ;
  assign n11340 = ( x107 & n11334 ) | ( x107 & ~n11339 ) | ( n11334 & ~n11339 ) ;
  assign n11341 = ( x107 & n10980 ) | ( x107 & ~n11083 ) | ( n10980 & ~n11083 ) ;
  assign n11342 = x107 & n10980 ;
  assign n11343 = ( ~n10985 & n11341 ) | ( ~n10985 & n11342 ) | ( n11341 & n11342 ) ;
  assign n11344 = ( n10985 & n11341 ) | ( n10985 & n11342 ) | ( n11341 & n11342 ) ;
  assign n11345 = ( n10985 & n11343 ) | ( n10985 & ~n11344 ) | ( n11343 & ~n11344 ) ;
  assign n11346 = ( x108 & n11340 ) | ( x108 & ~n11345 ) | ( n11340 & ~n11345 ) ;
  assign n11347 = ( x108 & n10986 ) | ( x108 & ~n11083 ) | ( n10986 & ~n11083 ) ;
  assign n11348 = x108 & n10986 ;
  assign n11349 = ( ~n10991 & n11347 ) | ( ~n10991 & n11348 ) | ( n11347 & n11348 ) ;
  assign n11350 = ( n10991 & n11347 ) | ( n10991 & n11348 ) | ( n11347 & n11348 ) ;
  assign n11351 = ( n10991 & n11349 ) | ( n10991 & ~n11350 ) | ( n11349 & ~n11350 ) ;
  assign n11352 = ( x109 & n11346 ) | ( x109 & ~n11351 ) | ( n11346 & ~n11351 ) ;
  assign n11353 = ( x109 & n10992 ) | ( x109 & ~n11083 ) | ( n10992 & ~n11083 ) ;
  assign n11354 = x109 & n10992 ;
  assign n11355 = ( ~n10997 & n11353 ) | ( ~n10997 & n11354 ) | ( n11353 & n11354 ) ;
  assign n11356 = ( n10997 & n11353 ) | ( n10997 & n11354 ) | ( n11353 & n11354 ) ;
  assign n11357 = ( n10997 & n11355 ) | ( n10997 & ~n11356 ) | ( n11355 & ~n11356 ) ;
  assign n11358 = ( x110 & n11352 ) | ( x110 & ~n11357 ) | ( n11352 & ~n11357 ) ;
  assign n11359 = ( x110 & n10998 ) | ( x110 & ~n11083 ) | ( n10998 & ~n11083 ) ;
  assign n11360 = x110 & n10998 ;
  assign n11361 = ( ~n11003 & n11359 ) | ( ~n11003 & n11360 ) | ( n11359 & n11360 ) ;
  assign n11362 = ( n11003 & n11359 ) | ( n11003 & n11360 ) | ( n11359 & n11360 ) ;
  assign n11363 = ( n11003 & n11361 ) | ( n11003 & ~n11362 ) | ( n11361 & ~n11362 ) ;
  assign n11364 = ( x111 & n11358 ) | ( x111 & ~n11363 ) | ( n11358 & ~n11363 ) ;
  assign n11365 = ( x111 & n11004 ) | ( x111 & ~n11083 ) | ( n11004 & ~n11083 ) ;
  assign n11366 = x111 & n11004 ;
  assign n11367 = ( ~n11009 & n11365 ) | ( ~n11009 & n11366 ) | ( n11365 & n11366 ) ;
  assign n11368 = ( n11009 & n11365 ) | ( n11009 & n11366 ) | ( n11365 & n11366 ) ;
  assign n11369 = ( n11009 & n11367 ) | ( n11009 & ~n11368 ) | ( n11367 & ~n11368 ) ;
  assign n11370 = ( x112 & n11364 ) | ( x112 & ~n11369 ) | ( n11364 & ~n11369 ) ;
  assign n11371 = ( x112 & n11010 ) | ( x112 & ~n11083 ) | ( n11010 & ~n11083 ) ;
  assign n11372 = x112 & n11010 ;
  assign n11373 = ( ~n11015 & n11371 ) | ( ~n11015 & n11372 ) | ( n11371 & n11372 ) ;
  assign n11374 = ( n11015 & n11371 ) | ( n11015 & n11372 ) | ( n11371 & n11372 ) ;
  assign n11375 = ( n11015 & n11373 ) | ( n11015 & ~n11374 ) | ( n11373 & ~n11374 ) ;
  assign n11376 = ( x113 & n11370 ) | ( x113 & ~n11375 ) | ( n11370 & ~n11375 ) ;
  assign n11377 = ( x113 & n11016 ) | ( x113 & ~n11083 ) | ( n11016 & ~n11083 ) ;
  assign n11378 = x113 & n11016 ;
  assign n11379 = ( ~n11021 & n11377 ) | ( ~n11021 & n11378 ) | ( n11377 & n11378 ) ;
  assign n11380 = ( n11021 & n11377 ) | ( n11021 & n11378 ) | ( n11377 & n11378 ) ;
  assign n11381 = ( n11021 & n11379 ) | ( n11021 & ~n11380 ) | ( n11379 & ~n11380 ) ;
  assign n11382 = ( x114 & n11376 ) | ( x114 & ~n11381 ) | ( n11376 & ~n11381 ) ;
  assign n11383 = ( x114 & n11022 ) | ( x114 & ~n11083 ) | ( n11022 & ~n11083 ) ;
  assign n11384 = x114 & n11022 ;
  assign n11385 = ( ~n11027 & n11383 ) | ( ~n11027 & n11384 ) | ( n11383 & n11384 ) ;
  assign n11386 = ( n11027 & n11383 ) | ( n11027 & n11384 ) | ( n11383 & n11384 ) ;
  assign n11387 = ( n11027 & n11385 ) | ( n11027 & ~n11386 ) | ( n11385 & ~n11386 ) ;
  assign n11388 = ( x115 & n11382 ) | ( x115 & ~n11387 ) | ( n11382 & ~n11387 ) ;
  assign n11389 = ( x115 & n11028 ) | ( x115 & ~n11083 ) | ( n11028 & ~n11083 ) ;
  assign n11390 = x115 & n11028 ;
  assign n11391 = ( ~n11033 & n11389 ) | ( ~n11033 & n11390 ) | ( n11389 & n11390 ) ;
  assign n11392 = ( n11033 & n11389 ) | ( n11033 & n11390 ) | ( n11389 & n11390 ) ;
  assign n11393 = ( n11033 & n11391 ) | ( n11033 & ~n11392 ) | ( n11391 & ~n11392 ) ;
  assign n11394 = ( x116 & n11388 ) | ( x116 & ~n11393 ) | ( n11388 & ~n11393 ) ;
  assign n11395 = ( x116 & n11034 ) | ( x116 & ~n11083 ) | ( n11034 & ~n11083 ) ;
  assign n11396 = x116 & n11034 ;
  assign n11397 = ( ~n11039 & n11395 ) | ( ~n11039 & n11396 ) | ( n11395 & n11396 ) ;
  assign n11398 = ( n11039 & n11395 ) | ( n11039 & n11396 ) | ( n11395 & n11396 ) ;
  assign n11399 = ( n11039 & n11397 ) | ( n11039 & ~n11398 ) | ( n11397 & ~n11398 ) ;
  assign n11400 = ( x117 & n11394 ) | ( x117 & ~n11399 ) | ( n11394 & ~n11399 ) ;
  assign n11401 = ( x117 & n11040 ) | ( x117 & ~n11083 ) | ( n11040 & ~n11083 ) ;
  assign n11402 = x117 & n11040 ;
  assign n11403 = ( ~n11045 & n11401 ) | ( ~n11045 & n11402 ) | ( n11401 & n11402 ) ;
  assign n11404 = ( n11045 & n11401 ) | ( n11045 & n11402 ) | ( n11401 & n11402 ) ;
  assign n11405 = ( n11045 & n11403 ) | ( n11045 & ~n11404 ) | ( n11403 & ~n11404 ) ;
  assign n11406 = ( x118 & n11400 ) | ( x118 & ~n11405 ) | ( n11400 & ~n11405 ) ;
  assign n11407 = ( x118 & n11046 ) | ( x118 & ~n11083 ) | ( n11046 & ~n11083 ) ;
  assign n11408 = x118 & n11046 ;
  assign n11409 = ( ~n11051 & n11407 ) | ( ~n11051 & n11408 ) | ( n11407 & n11408 ) ;
  assign n11410 = ( n11051 & n11407 ) | ( n11051 & n11408 ) | ( n11407 & n11408 ) ;
  assign n11411 = ( n11051 & n11409 ) | ( n11051 & ~n11410 ) | ( n11409 & ~n11410 ) ;
  assign n11412 = ( x119 & n11406 ) | ( x119 & ~n11411 ) | ( n11406 & ~n11411 ) ;
  assign n11413 = ( x119 & n11052 ) | ( x119 & ~n11083 ) | ( n11052 & ~n11083 ) ;
  assign n11414 = x119 & n11052 ;
  assign n11415 = ( ~n11057 & n11413 ) | ( ~n11057 & n11414 ) | ( n11413 & n11414 ) ;
  assign n11416 = ( n11057 & n11413 ) | ( n11057 & n11414 ) | ( n11413 & n11414 ) ;
  assign n11417 = ( n11057 & n11415 ) | ( n11057 & ~n11416 ) | ( n11415 & ~n11416 ) ;
  assign n11418 = ( x120 & n11412 ) | ( x120 & ~n11417 ) | ( n11412 & ~n11417 ) ;
  assign n11419 = ( x120 & n11058 ) | ( x120 & ~n11083 ) | ( n11058 & ~n11083 ) ;
  assign n11420 = x120 & n11058 ;
  assign n11421 = ( ~n11063 & n11419 ) | ( ~n11063 & n11420 ) | ( n11419 & n11420 ) ;
  assign n11422 = ( n11063 & n11419 ) | ( n11063 & n11420 ) | ( n11419 & n11420 ) ;
  assign n11423 = ( n11063 & n11421 ) | ( n11063 & ~n11422 ) | ( n11421 & ~n11422 ) ;
  assign n11424 = ( x121 & n11418 ) | ( x121 & ~n11423 ) | ( n11418 & ~n11423 ) ;
  assign n11425 = ( x121 & n11064 ) | ( x121 & ~n11083 ) | ( n11064 & ~n11083 ) ;
  assign n11426 = x121 & n11064 ;
  assign n11427 = ( ~n11069 & n11425 ) | ( ~n11069 & n11426 ) | ( n11425 & n11426 ) ;
  assign n11428 = ( n11069 & n11425 ) | ( n11069 & n11426 ) | ( n11425 & n11426 ) ;
  assign n11429 = ( n11069 & n11427 ) | ( n11069 & ~n11428 ) | ( n11427 & ~n11428 ) ;
  assign n11430 = ( x122 & n11424 ) | ( x122 & ~n11429 ) | ( n11424 & ~n11429 ) ;
  assign n11431 = ( x122 & n11070 ) | ( x122 & ~n11083 ) | ( n11070 & ~n11083 ) ;
  assign n11432 = x122 & n11070 ;
  assign n11433 = ( ~n11075 & n11431 ) | ( ~n11075 & n11432 ) | ( n11431 & n11432 ) ;
  assign n11434 = ( n11075 & n11431 ) | ( n11075 & n11432 ) | ( n11431 & n11432 ) ;
  assign n11435 = ( n11075 & n11433 ) | ( n11075 & ~n11434 ) | ( n11433 & ~n11434 ) ;
  assign n11436 = ( x123 & n11430 ) | ( x123 & ~n11435 ) | ( n11430 & ~n11435 ) ;
  assign n11437 = ( x123 & n11076 ) | ( x123 & ~n11083 ) | ( n11076 & ~n11083 ) ;
  assign n11438 = x123 & n11076 ;
  assign n11439 = ( ~n10729 & n11437 ) | ( ~n10729 & n11438 ) | ( n11437 & n11438 ) ;
  assign n11440 = ( n10729 & n11437 ) | ( n10729 & n11438 ) | ( n11437 & n11438 ) ;
  assign n11441 = ( n10729 & n11439 ) | ( n10729 & ~n11440 ) | ( n11439 & ~n11440 ) ;
  assign n11442 = ( x124 & n11436 ) | ( x124 & ~n11441 ) | ( n11436 & ~n11441 ) ;
  assign n11443 = n133 & n10019 ;
  assign n11444 = n11078 & n11443 ;
  assign n11445 = n389 | n11444 ;
  assign n11446 = ~x127 & n11445 ;
  assign n11447 = ~x126 & n11446 ;
  assign n11448 = n132 & ~n11447 ;
  assign n11449 = ~x125 & n11447 ;
  assign n11450 = ( n11442 & n11448 ) | ( n11442 & ~n11449 ) | ( n11448 & ~n11449 ) ;
  assign n11451 = ~x2 & n11450 ;
  assign n11452 = ( x2 & ~x64 ) | ( x2 & n11450 ) | ( ~x64 & n11450 ) ;
  assign n11453 = ( n391 & ~n11451 ) | ( n391 & n11452 ) | ( ~n11451 & n11452 ) ;
  assign n11454 = ( x65 & n390 ) | ( x65 & ~n11453 ) | ( n390 & ~n11453 ) ;
  assign n11455 = ( x65 & n391 ) | ( x65 & n11450 ) | ( n391 & n11450 ) ;
  assign n11456 = x65 | n391 ;
  assign n11457 = ( ~n11087 & n11455 ) | ( ~n11087 & n11456 ) | ( n11455 & n11456 ) ;
  assign n11458 = ( n11087 & n11455 ) | ( n11087 & n11456 ) | ( n11455 & n11456 ) ;
  assign n11459 = ( n11087 & n11457 ) | ( n11087 & ~n11458 ) | ( n11457 & ~n11458 ) ;
  assign n11460 = ( x66 & n11454 ) | ( x66 & ~n11459 ) | ( n11454 & ~n11459 ) ;
  assign n11461 = ( x66 & n11088 ) | ( x66 & n11450 ) | ( n11088 & n11450 ) ;
  assign n11462 = x66 | n11088 ;
  assign n11463 = ( ~n11093 & n11461 ) | ( ~n11093 & n11462 ) | ( n11461 & n11462 ) ;
  assign n11464 = ( n11093 & n11461 ) | ( n11093 & n11462 ) | ( n11461 & n11462 ) ;
  assign n11465 = ( n11093 & n11463 ) | ( n11093 & ~n11464 ) | ( n11463 & ~n11464 ) ;
  assign n11466 = ( x67 & n11460 ) | ( x67 & ~n11465 ) | ( n11460 & ~n11465 ) ;
  assign n11467 = ( x67 & n11094 ) | ( x67 & ~n11450 ) | ( n11094 & ~n11450 ) ;
  assign n11468 = x67 & n11094 ;
  assign n11469 = ( ~n11099 & n11467 ) | ( ~n11099 & n11468 ) | ( n11467 & n11468 ) ;
  assign n11470 = ( n11099 & n11467 ) | ( n11099 & n11468 ) | ( n11467 & n11468 ) ;
  assign n11471 = ( n11099 & n11469 ) | ( n11099 & ~n11470 ) | ( n11469 & ~n11470 ) ;
  assign n11472 = ( x68 & n11466 ) | ( x68 & ~n11471 ) | ( n11466 & ~n11471 ) ;
  assign n11473 = ( x68 & n11100 ) | ( x68 & ~n11450 ) | ( n11100 & ~n11450 ) ;
  assign n11474 = x68 & n11100 ;
  assign n11475 = ( ~n11105 & n11473 ) | ( ~n11105 & n11474 ) | ( n11473 & n11474 ) ;
  assign n11476 = ( n11105 & n11473 ) | ( n11105 & n11474 ) | ( n11473 & n11474 ) ;
  assign n11477 = ( n11105 & n11475 ) | ( n11105 & ~n11476 ) | ( n11475 & ~n11476 ) ;
  assign n11478 = ( x69 & n11472 ) | ( x69 & ~n11477 ) | ( n11472 & ~n11477 ) ;
  assign n11479 = ( x69 & n11106 ) | ( x69 & ~n11450 ) | ( n11106 & ~n11450 ) ;
  assign n11480 = x69 & n11106 ;
  assign n11481 = ( ~n11111 & n11479 ) | ( ~n11111 & n11480 ) | ( n11479 & n11480 ) ;
  assign n11482 = ( n11111 & n11479 ) | ( n11111 & n11480 ) | ( n11479 & n11480 ) ;
  assign n11483 = ( n11111 & n11481 ) | ( n11111 & ~n11482 ) | ( n11481 & ~n11482 ) ;
  assign n11484 = ( x70 & n11478 ) | ( x70 & ~n11483 ) | ( n11478 & ~n11483 ) ;
  assign n11485 = ( x70 & n11112 ) | ( x70 & ~n11450 ) | ( n11112 & ~n11450 ) ;
  assign n11486 = x70 & n11112 ;
  assign n11487 = ( ~n11117 & n11485 ) | ( ~n11117 & n11486 ) | ( n11485 & n11486 ) ;
  assign n11488 = ( n11117 & n11485 ) | ( n11117 & n11486 ) | ( n11485 & n11486 ) ;
  assign n11489 = ( n11117 & n11487 ) | ( n11117 & ~n11488 ) | ( n11487 & ~n11488 ) ;
  assign n11490 = ( x71 & n11484 ) | ( x71 & ~n11489 ) | ( n11484 & ~n11489 ) ;
  assign n11491 = ( x71 & n11118 ) | ( x71 & ~n11450 ) | ( n11118 & ~n11450 ) ;
  assign n11492 = x71 & n11118 ;
  assign n11493 = ( ~n11123 & n11491 ) | ( ~n11123 & n11492 ) | ( n11491 & n11492 ) ;
  assign n11494 = ( n11123 & n11491 ) | ( n11123 & n11492 ) | ( n11491 & n11492 ) ;
  assign n11495 = ( n11123 & n11493 ) | ( n11123 & ~n11494 ) | ( n11493 & ~n11494 ) ;
  assign n11496 = ( x72 & n11490 ) | ( x72 & ~n11495 ) | ( n11490 & ~n11495 ) ;
  assign n11497 = ( x72 & n11124 ) | ( x72 & ~n11450 ) | ( n11124 & ~n11450 ) ;
  assign n11498 = x72 & n11124 ;
  assign n11499 = ( ~n11129 & n11497 ) | ( ~n11129 & n11498 ) | ( n11497 & n11498 ) ;
  assign n11500 = ( n11129 & n11497 ) | ( n11129 & n11498 ) | ( n11497 & n11498 ) ;
  assign n11501 = ( n11129 & n11499 ) | ( n11129 & ~n11500 ) | ( n11499 & ~n11500 ) ;
  assign n11502 = ( x73 & n11496 ) | ( x73 & ~n11501 ) | ( n11496 & ~n11501 ) ;
  assign n11503 = ( x73 & n11130 ) | ( x73 & ~n11450 ) | ( n11130 & ~n11450 ) ;
  assign n11504 = x73 & n11130 ;
  assign n11505 = ( ~n11135 & n11503 ) | ( ~n11135 & n11504 ) | ( n11503 & n11504 ) ;
  assign n11506 = ( n11135 & n11503 ) | ( n11135 & n11504 ) | ( n11503 & n11504 ) ;
  assign n11507 = ( n11135 & n11505 ) | ( n11135 & ~n11506 ) | ( n11505 & ~n11506 ) ;
  assign n11508 = ( x74 & n11502 ) | ( x74 & ~n11507 ) | ( n11502 & ~n11507 ) ;
  assign n11509 = ( x74 & n11136 ) | ( x74 & ~n11450 ) | ( n11136 & ~n11450 ) ;
  assign n11510 = x74 & n11136 ;
  assign n11511 = ( ~n11141 & n11509 ) | ( ~n11141 & n11510 ) | ( n11509 & n11510 ) ;
  assign n11512 = ( n11141 & n11509 ) | ( n11141 & n11510 ) | ( n11509 & n11510 ) ;
  assign n11513 = ( n11141 & n11511 ) | ( n11141 & ~n11512 ) | ( n11511 & ~n11512 ) ;
  assign n11514 = ( x75 & n11508 ) | ( x75 & ~n11513 ) | ( n11508 & ~n11513 ) ;
  assign n11515 = ( x75 & n11142 ) | ( x75 & ~n11450 ) | ( n11142 & ~n11450 ) ;
  assign n11516 = x75 & n11142 ;
  assign n11517 = ( ~n11147 & n11515 ) | ( ~n11147 & n11516 ) | ( n11515 & n11516 ) ;
  assign n11518 = ( n11147 & n11515 ) | ( n11147 & n11516 ) | ( n11515 & n11516 ) ;
  assign n11519 = ( n11147 & n11517 ) | ( n11147 & ~n11518 ) | ( n11517 & ~n11518 ) ;
  assign n11520 = ( x76 & n11514 ) | ( x76 & ~n11519 ) | ( n11514 & ~n11519 ) ;
  assign n11521 = ( x76 & n11148 ) | ( x76 & ~n11450 ) | ( n11148 & ~n11450 ) ;
  assign n11522 = x76 & n11148 ;
  assign n11523 = ( ~n11153 & n11521 ) | ( ~n11153 & n11522 ) | ( n11521 & n11522 ) ;
  assign n11524 = ( n11153 & n11521 ) | ( n11153 & n11522 ) | ( n11521 & n11522 ) ;
  assign n11525 = ( n11153 & n11523 ) | ( n11153 & ~n11524 ) | ( n11523 & ~n11524 ) ;
  assign n11526 = ( x77 & n11520 ) | ( x77 & ~n11525 ) | ( n11520 & ~n11525 ) ;
  assign n11527 = ( x77 & n11154 ) | ( x77 & ~n11450 ) | ( n11154 & ~n11450 ) ;
  assign n11528 = x77 & n11154 ;
  assign n11529 = ( ~n11159 & n11527 ) | ( ~n11159 & n11528 ) | ( n11527 & n11528 ) ;
  assign n11530 = ( n11159 & n11527 ) | ( n11159 & n11528 ) | ( n11527 & n11528 ) ;
  assign n11531 = ( n11159 & n11529 ) | ( n11159 & ~n11530 ) | ( n11529 & ~n11530 ) ;
  assign n11532 = ( x78 & n11526 ) | ( x78 & ~n11531 ) | ( n11526 & ~n11531 ) ;
  assign n11533 = ( x78 & n11160 ) | ( x78 & ~n11450 ) | ( n11160 & ~n11450 ) ;
  assign n11534 = x78 & n11160 ;
  assign n11535 = ( ~n11165 & n11533 ) | ( ~n11165 & n11534 ) | ( n11533 & n11534 ) ;
  assign n11536 = ( n11165 & n11533 ) | ( n11165 & n11534 ) | ( n11533 & n11534 ) ;
  assign n11537 = ( n11165 & n11535 ) | ( n11165 & ~n11536 ) | ( n11535 & ~n11536 ) ;
  assign n11538 = ( x79 & n11532 ) | ( x79 & ~n11537 ) | ( n11532 & ~n11537 ) ;
  assign n11539 = ( x79 & n11166 ) | ( x79 & ~n11450 ) | ( n11166 & ~n11450 ) ;
  assign n11540 = x79 & n11166 ;
  assign n11541 = ( ~n11171 & n11539 ) | ( ~n11171 & n11540 ) | ( n11539 & n11540 ) ;
  assign n11542 = ( n11171 & n11539 ) | ( n11171 & n11540 ) | ( n11539 & n11540 ) ;
  assign n11543 = ( n11171 & n11541 ) | ( n11171 & ~n11542 ) | ( n11541 & ~n11542 ) ;
  assign n11544 = ( x80 & n11538 ) | ( x80 & ~n11543 ) | ( n11538 & ~n11543 ) ;
  assign n11545 = ( x80 & n11172 ) | ( x80 & ~n11450 ) | ( n11172 & ~n11450 ) ;
  assign n11546 = x80 & n11172 ;
  assign n11547 = ( ~n11177 & n11545 ) | ( ~n11177 & n11546 ) | ( n11545 & n11546 ) ;
  assign n11548 = ( n11177 & n11545 ) | ( n11177 & n11546 ) | ( n11545 & n11546 ) ;
  assign n11549 = ( n11177 & n11547 ) | ( n11177 & ~n11548 ) | ( n11547 & ~n11548 ) ;
  assign n11550 = ( x81 & n11544 ) | ( x81 & ~n11549 ) | ( n11544 & ~n11549 ) ;
  assign n11551 = ( x81 & n11178 ) | ( x81 & ~n11450 ) | ( n11178 & ~n11450 ) ;
  assign n11552 = x81 & n11178 ;
  assign n11553 = ( ~n11183 & n11551 ) | ( ~n11183 & n11552 ) | ( n11551 & n11552 ) ;
  assign n11554 = ( n11183 & n11551 ) | ( n11183 & n11552 ) | ( n11551 & n11552 ) ;
  assign n11555 = ( n11183 & n11553 ) | ( n11183 & ~n11554 ) | ( n11553 & ~n11554 ) ;
  assign n11556 = ( x82 & n11550 ) | ( x82 & ~n11555 ) | ( n11550 & ~n11555 ) ;
  assign n11557 = ( x82 & n11184 ) | ( x82 & ~n11450 ) | ( n11184 & ~n11450 ) ;
  assign n11558 = x82 & n11184 ;
  assign n11559 = ( ~n11189 & n11557 ) | ( ~n11189 & n11558 ) | ( n11557 & n11558 ) ;
  assign n11560 = ( n11189 & n11557 ) | ( n11189 & n11558 ) | ( n11557 & n11558 ) ;
  assign n11561 = ( n11189 & n11559 ) | ( n11189 & ~n11560 ) | ( n11559 & ~n11560 ) ;
  assign n11562 = ( x83 & n11556 ) | ( x83 & ~n11561 ) | ( n11556 & ~n11561 ) ;
  assign n11563 = ( x83 & n11190 ) | ( x83 & ~n11450 ) | ( n11190 & ~n11450 ) ;
  assign n11564 = x83 & n11190 ;
  assign n11565 = ( ~n11195 & n11563 ) | ( ~n11195 & n11564 ) | ( n11563 & n11564 ) ;
  assign n11566 = ( n11195 & n11563 ) | ( n11195 & n11564 ) | ( n11563 & n11564 ) ;
  assign n11567 = ( n11195 & n11565 ) | ( n11195 & ~n11566 ) | ( n11565 & ~n11566 ) ;
  assign n11568 = ( x84 & n11562 ) | ( x84 & ~n11567 ) | ( n11562 & ~n11567 ) ;
  assign n11569 = ( x84 & n11196 ) | ( x84 & ~n11450 ) | ( n11196 & ~n11450 ) ;
  assign n11570 = x84 & n11196 ;
  assign n11571 = ( ~n11201 & n11569 ) | ( ~n11201 & n11570 ) | ( n11569 & n11570 ) ;
  assign n11572 = ( n11201 & n11569 ) | ( n11201 & n11570 ) | ( n11569 & n11570 ) ;
  assign n11573 = ( n11201 & n11571 ) | ( n11201 & ~n11572 ) | ( n11571 & ~n11572 ) ;
  assign n11574 = ( x85 & n11568 ) | ( x85 & ~n11573 ) | ( n11568 & ~n11573 ) ;
  assign n11575 = ( x85 & n11202 ) | ( x85 & ~n11450 ) | ( n11202 & ~n11450 ) ;
  assign n11576 = x85 & n11202 ;
  assign n11577 = ( ~n11207 & n11575 ) | ( ~n11207 & n11576 ) | ( n11575 & n11576 ) ;
  assign n11578 = ( n11207 & n11575 ) | ( n11207 & n11576 ) | ( n11575 & n11576 ) ;
  assign n11579 = ( n11207 & n11577 ) | ( n11207 & ~n11578 ) | ( n11577 & ~n11578 ) ;
  assign n11580 = ( x86 & n11574 ) | ( x86 & ~n11579 ) | ( n11574 & ~n11579 ) ;
  assign n11581 = ( x86 & n11208 ) | ( x86 & ~n11450 ) | ( n11208 & ~n11450 ) ;
  assign n11582 = x86 & n11208 ;
  assign n11583 = ( ~n11213 & n11581 ) | ( ~n11213 & n11582 ) | ( n11581 & n11582 ) ;
  assign n11584 = ( n11213 & n11581 ) | ( n11213 & n11582 ) | ( n11581 & n11582 ) ;
  assign n11585 = ( n11213 & n11583 ) | ( n11213 & ~n11584 ) | ( n11583 & ~n11584 ) ;
  assign n11586 = ( x87 & n11580 ) | ( x87 & ~n11585 ) | ( n11580 & ~n11585 ) ;
  assign n11587 = ( x87 & n11214 ) | ( x87 & ~n11450 ) | ( n11214 & ~n11450 ) ;
  assign n11588 = x87 & n11214 ;
  assign n11589 = ( ~n11219 & n11587 ) | ( ~n11219 & n11588 ) | ( n11587 & n11588 ) ;
  assign n11590 = ( n11219 & n11587 ) | ( n11219 & n11588 ) | ( n11587 & n11588 ) ;
  assign n11591 = ( n11219 & n11589 ) | ( n11219 & ~n11590 ) | ( n11589 & ~n11590 ) ;
  assign n11592 = ( x88 & n11586 ) | ( x88 & ~n11591 ) | ( n11586 & ~n11591 ) ;
  assign n11593 = ( x88 & n11220 ) | ( x88 & ~n11450 ) | ( n11220 & ~n11450 ) ;
  assign n11594 = x88 & n11220 ;
  assign n11595 = ( ~n11225 & n11593 ) | ( ~n11225 & n11594 ) | ( n11593 & n11594 ) ;
  assign n11596 = ( n11225 & n11593 ) | ( n11225 & n11594 ) | ( n11593 & n11594 ) ;
  assign n11597 = ( n11225 & n11595 ) | ( n11225 & ~n11596 ) | ( n11595 & ~n11596 ) ;
  assign n11598 = ( x89 & n11592 ) | ( x89 & ~n11597 ) | ( n11592 & ~n11597 ) ;
  assign n11599 = ( x89 & n11226 ) | ( x89 & ~n11450 ) | ( n11226 & ~n11450 ) ;
  assign n11600 = x89 & n11226 ;
  assign n11601 = ( ~n11231 & n11599 ) | ( ~n11231 & n11600 ) | ( n11599 & n11600 ) ;
  assign n11602 = ( n11231 & n11599 ) | ( n11231 & n11600 ) | ( n11599 & n11600 ) ;
  assign n11603 = ( n11231 & n11601 ) | ( n11231 & ~n11602 ) | ( n11601 & ~n11602 ) ;
  assign n11604 = ( x90 & n11598 ) | ( x90 & ~n11603 ) | ( n11598 & ~n11603 ) ;
  assign n11605 = ( x90 & n11232 ) | ( x90 & ~n11450 ) | ( n11232 & ~n11450 ) ;
  assign n11606 = x90 & n11232 ;
  assign n11607 = ( ~n11237 & n11605 ) | ( ~n11237 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11608 = ( n11237 & n11605 ) | ( n11237 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11609 = ( n11237 & n11607 ) | ( n11237 & ~n11608 ) | ( n11607 & ~n11608 ) ;
  assign n11610 = ( x91 & n11604 ) | ( x91 & ~n11609 ) | ( n11604 & ~n11609 ) ;
  assign n11611 = ( x91 & n11238 ) | ( x91 & ~n11450 ) | ( n11238 & ~n11450 ) ;
  assign n11612 = x91 & n11238 ;
  assign n11613 = ( ~n11243 & n11611 ) | ( ~n11243 & n11612 ) | ( n11611 & n11612 ) ;
  assign n11614 = ( n11243 & n11611 ) | ( n11243 & n11612 ) | ( n11611 & n11612 ) ;
  assign n11615 = ( n11243 & n11613 ) | ( n11243 & ~n11614 ) | ( n11613 & ~n11614 ) ;
  assign n11616 = ( x92 & n11610 ) | ( x92 & ~n11615 ) | ( n11610 & ~n11615 ) ;
  assign n11617 = ( x92 & n11244 ) | ( x92 & ~n11450 ) | ( n11244 & ~n11450 ) ;
  assign n11618 = x92 & n11244 ;
  assign n11619 = ( ~n11249 & n11617 ) | ( ~n11249 & n11618 ) | ( n11617 & n11618 ) ;
  assign n11620 = ( n11249 & n11617 ) | ( n11249 & n11618 ) | ( n11617 & n11618 ) ;
  assign n11621 = ( n11249 & n11619 ) | ( n11249 & ~n11620 ) | ( n11619 & ~n11620 ) ;
  assign n11622 = ( x93 & n11616 ) | ( x93 & ~n11621 ) | ( n11616 & ~n11621 ) ;
  assign n11623 = ( x93 & n11250 ) | ( x93 & ~n11450 ) | ( n11250 & ~n11450 ) ;
  assign n11624 = x93 & n11250 ;
  assign n11625 = ( ~n11255 & n11623 ) | ( ~n11255 & n11624 ) | ( n11623 & n11624 ) ;
  assign n11626 = ( n11255 & n11623 ) | ( n11255 & n11624 ) | ( n11623 & n11624 ) ;
  assign n11627 = ( n11255 & n11625 ) | ( n11255 & ~n11626 ) | ( n11625 & ~n11626 ) ;
  assign n11628 = ( x94 & n11622 ) | ( x94 & ~n11627 ) | ( n11622 & ~n11627 ) ;
  assign n11629 = ( x94 & n11256 ) | ( x94 & ~n11450 ) | ( n11256 & ~n11450 ) ;
  assign n11630 = x94 & n11256 ;
  assign n11631 = ( ~n11261 & n11629 ) | ( ~n11261 & n11630 ) | ( n11629 & n11630 ) ;
  assign n11632 = ( n11261 & n11629 ) | ( n11261 & n11630 ) | ( n11629 & n11630 ) ;
  assign n11633 = ( n11261 & n11631 ) | ( n11261 & ~n11632 ) | ( n11631 & ~n11632 ) ;
  assign n11634 = ( x95 & n11628 ) | ( x95 & ~n11633 ) | ( n11628 & ~n11633 ) ;
  assign n11635 = ( x95 & n11262 ) | ( x95 & ~n11450 ) | ( n11262 & ~n11450 ) ;
  assign n11636 = x95 & n11262 ;
  assign n11637 = ( ~n11267 & n11635 ) | ( ~n11267 & n11636 ) | ( n11635 & n11636 ) ;
  assign n11638 = ( n11267 & n11635 ) | ( n11267 & n11636 ) | ( n11635 & n11636 ) ;
  assign n11639 = ( n11267 & n11637 ) | ( n11267 & ~n11638 ) | ( n11637 & ~n11638 ) ;
  assign n11640 = ( x96 & n11634 ) | ( x96 & ~n11639 ) | ( n11634 & ~n11639 ) ;
  assign n11641 = ( x96 & n11268 ) | ( x96 & ~n11450 ) | ( n11268 & ~n11450 ) ;
  assign n11642 = x96 & n11268 ;
  assign n11643 = ( ~n11273 & n11641 ) | ( ~n11273 & n11642 ) | ( n11641 & n11642 ) ;
  assign n11644 = ( n11273 & n11641 ) | ( n11273 & n11642 ) | ( n11641 & n11642 ) ;
  assign n11645 = ( n11273 & n11643 ) | ( n11273 & ~n11644 ) | ( n11643 & ~n11644 ) ;
  assign n11646 = ( x97 & n11640 ) | ( x97 & ~n11645 ) | ( n11640 & ~n11645 ) ;
  assign n11647 = ( x97 & n11274 ) | ( x97 & ~n11450 ) | ( n11274 & ~n11450 ) ;
  assign n11648 = x97 & n11274 ;
  assign n11649 = ( ~n11279 & n11647 ) | ( ~n11279 & n11648 ) | ( n11647 & n11648 ) ;
  assign n11650 = ( n11279 & n11647 ) | ( n11279 & n11648 ) | ( n11647 & n11648 ) ;
  assign n11651 = ( n11279 & n11649 ) | ( n11279 & ~n11650 ) | ( n11649 & ~n11650 ) ;
  assign n11652 = ( x98 & n11646 ) | ( x98 & ~n11651 ) | ( n11646 & ~n11651 ) ;
  assign n11653 = ( x98 & n11280 ) | ( x98 & ~n11450 ) | ( n11280 & ~n11450 ) ;
  assign n11654 = x98 & n11280 ;
  assign n11655 = ( ~n11285 & n11653 ) | ( ~n11285 & n11654 ) | ( n11653 & n11654 ) ;
  assign n11656 = ( n11285 & n11653 ) | ( n11285 & n11654 ) | ( n11653 & n11654 ) ;
  assign n11657 = ( n11285 & n11655 ) | ( n11285 & ~n11656 ) | ( n11655 & ~n11656 ) ;
  assign n11658 = ( x99 & n11652 ) | ( x99 & ~n11657 ) | ( n11652 & ~n11657 ) ;
  assign n11659 = ( x99 & n11286 ) | ( x99 & ~n11450 ) | ( n11286 & ~n11450 ) ;
  assign n11660 = x99 & n11286 ;
  assign n11661 = ( ~n11291 & n11659 ) | ( ~n11291 & n11660 ) | ( n11659 & n11660 ) ;
  assign n11662 = ( n11291 & n11659 ) | ( n11291 & n11660 ) | ( n11659 & n11660 ) ;
  assign n11663 = ( n11291 & n11661 ) | ( n11291 & ~n11662 ) | ( n11661 & ~n11662 ) ;
  assign n11664 = ( x100 & n11658 ) | ( x100 & ~n11663 ) | ( n11658 & ~n11663 ) ;
  assign n11665 = ( x100 & n11292 ) | ( x100 & ~n11450 ) | ( n11292 & ~n11450 ) ;
  assign n11666 = x100 & n11292 ;
  assign n11667 = ( ~n11297 & n11665 ) | ( ~n11297 & n11666 ) | ( n11665 & n11666 ) ;
  assign n11668 = ( n11297 & n11665 ) | ( n11297 & n11666 ) | ( n11665 & n11666 ) ;
  assign n11669 = ( n11297 & n11667 ) | ( n11297 & ~n11668 ) | ( n11667 & ~n11668 ) ;
  assign n11670 = ( x101 & n11664 ) | ( x101 & ~n11669 ) | ( n11664 & ~n11669 ) ;
  assign n11671 = ( x101 & n11298 ) | ( x101 & ~n11450 ) | ( n11298 & ~n11450 ) ;
  assign n11672 = x101 & n11298 ;
  assign n11673 = ( ~n11303 & n11671 ) | ( ~n11303 & n11672 ) | ( n11671 & n11672 ) ;
  assign n11674 = ( n11303 & n11671 ) | ( n11303 & n11672 ) | ( n11671 & n11672 ) ;
  assign n11675 = ( n11303 & n11673 ) | ( n11303 & ~n11674 ) | ( n11673 & ~n11674 ) ;
  assign n11676 = ( x102 & n11670 ) | ( x102 & ~n11675 ) | ( n11670 & ~n11675 ) ;
  assign n11677 = ( x102 & n11304 ) | ( x102 & ~n11450 ) | ( n11304 & ~n11450 ) ;
  assign n11678 = x102 & n11304 ;
  assign n11679 = ( ~n11309 & n11677 ) | ( ~n11309 & n11678 ) | ( n11677 & n11678 ) ;
  assign n11680 = ( n11309 & n11677 ) | ( n11309 & n11678 ) | ( n11677 & n11678 ) ;
  assign n11681 = ( n11309 & n11679 ) | ( n11309 & ~n11680 ) | ( n11679 & ~n11680 ) ;
  assign n11682 = ( x103 & n11676 ) | ( x103 & ~n11681 ) | ( n11676 & ~n11681 ) ;
  assign n11683 = ( x103 & n11310 ) | ( x103 & ~n11450 ) | ( n11310 & ~n11450 ) ;
  assign n11684 = x103 & n11310 ;
  assign n11685 = ( ~n11315 & n11683 ) | ( ~n11315 & n11684 ) | ( n11683 & n11684 ) ;
  assign n11686 = ( n11315 & n11683 ) | ( n11315 & n11684 ) | ( n11683 & n11684 ) ;
  assign n11687 = ( n11315 & n11685 ) | ( n11315 & ~n11686 ) | ( n11685 & ~n11686 ) ;
  assign n11688 = ( x104 & n11682 ) | ( x104 & ~n11687 ) | ( n11682 & ~n11687 ) ;
  assign n11689 = ( x104 & n11316 ) | ( x104 & ~n11450 ) | ( n11316 & ~n11450 ) ;
  assign n11690 = x104 & n11316 ;
  assign n11691 = ( ~n11321 & n11689 ) | ( ~n11321 & n11690 ) | ( n11689 & n11690 ) ;
  assign n11692 = ( n11321 & n11689 ) | ( n11321 & n11690 ) | ( n11689 & n11690 ) ;
  assign n11693 = ( n11321 & n11691 ) | ( n11321 & ~n11692 ) | ( n11691 & ~n11692 ) ;
  assign n11694 = ( x105 & n11688 ) | ( x105 & ~n11693 ) | ( n11688 & ~n11693 ) ;
  assign n11695 = ( x105 & n11322 ) | ( x105 & ~n11450 ) | ( n11322 & ~n11450 ) ;
  assign n11696 = x105 & n11322 ;
  assign n11697 = ( ~n11327 & n11695 ) | ( ~n11327 & n11696 ) | ( n11695 & n11696 ) ;
  assign n11698 = ( n11327 & n11695 ) | ( n11327 & n11696 ) | ( n11695 & n11696 ) ;
  assign n11699 = ( n11327 & n11697 ) | ( n11327 & ~n11698 ) | ( n11697 & ~n11698 ) ;
  assign n11700 = ( x106 & n11694 ) | ( x106 & ~n11699 ) | ( n11694 & ~n11699 ) ;
  assign n11701 = ( x106 & n11328 ) | ( x106 & ~n11450 ) | ( n11328 & ~n11450 ) ;
  assign n11702 = x106 & n11328 ;
  assign n11703 = ( ~n11333 & n11701 ) | ( ~n11333 & n11702 ) | ( n11701 & n11702 ) ;
  assign n11704 = ( n11333 & n11701 ) | ( n11333 & n11702 ) | ( n11701 & n11702 ) ;
  assign n11705 = ( n11333 & n11703 ) | ( n11333 & ~n11704 ) | ( n11703 & ~n11704 ) ;
  assign n11706 = ( x107 & n11700 ) | ( x107 & ~n11705 ) | ( n11700 & ~n11705 ) ;
  assign n11707 = ( x107 & n11334 ) | ( x107 & ~n11450 ) | ( n11334 & ~n11450 ) ;
  assign n11708 = x107 & n11334 ;
  assign n11709 = ( ~n11339 & n11707 ) | ( ~n11339 & n11708 ) | ( n11707 & n11708 ) ;
  assign n11710 = ( n11339 & n11707 ) | ( n11339 & n11708 ) | ( n11707 & n11708 ) ;
  assign n11711 = ( n11339 & n11709 ) | ( n11339 & ~n11710 ) | ( n11709 & ~n11710 ) ;
  assign n11712 = ( x108 & n11706 ) | ( x108 & ~n11711 ) | ( n11706 & ~n11711 ) ;
  assign n11713 = ( x108 & n11340 ) | ( x108 & ~n11450 ) | ( n11340 & ~n11450 ) ;
  assign n11714 = x108 & n11340 ;
  assign n11715 = ( ~n11345 & n11713 ) | ( ~n11345 & n11714 ) | ( n11713 & n11714 ) ;
  assign n11716 = ( n11345 & n11713 ) | ( n11345 & n11714 ) | ( n11713 & n11714 ) ;
  assign n11717 = ( n11345 & n11715 ) | ( n11345 & ~n11716 ) | ( n11715 & ~n11716 ) ;
  assign n11718 = ( x109 & n11712 ) | ( x109 & ~n11717 ) | ( n11712 & ~n11717 ) ;
  assign n11719 = ( x109 & n11346 ) | ( x109 & ~n11450 ) | ( n11346 & ~n11450 ) ;
  assign n11720 = x109 & n11346 ;
  assign n11721 = ( ~n11351 & n11719 ) | ( ~n11351 & n11720 ) | ( n11719 & n11720 ) ;
  assign n11722 = ( n11351 & n11719 ) | ( n11351 & n11720 ) | ( n11719 & n11720 ) ;
  assign n11723 = ( n11351 & n11721 ) | ( n11351 & ~n11722 ) | ( n11721 & ~n11722 ) ;
  assign n11724 = ( x110 & n11718 ) | ( x110 & ~n11723 ) | ( n11718 & ~n11723 ) ;
  assign n11725 = ( x110 & n11352 ) | ( x110 & ~n11450 ) | ( n11352 & ~n11450 ) ;
  assign n11726 = x110 & n11352 ;
  assign n11727 = ( ~n11357 & n11725 ) | ( ~n11357 & n11726 ) | ( n11725 & n11726 ) ;
  assign n11728 = ( n11357 & n11725 ) | ( n11357 & n11726 ) | ( n11725 & n11726 ) ;
  assign n11729 = ( n11357 & n11727 ) | ( n11357 & ~n11728 ) | ( n11727 & ~n11728 ) ;
  assign n11730 = ( x111 & n11724 ) | ( x111 & ~n11729 ) | ( n11724 & ~n11729 ) ;
  assign n11731 = ( x111 & n11358 ) | ( x111 & ~n11450 ) | ( n11358 & ~n11450 ) ;
  assign n11732 = x111 & n11358 ;
  assign n11733 = ( ~n11363 & n11731 ) | ( ~n11363 & n11732 ) | ( n11731 & n11732 ) ;
  assign n11734 = ( n11363 & n11731 ) | ( n11363 & n11732 ) | ( n11731 & n11732 ) ;
  assign n11735 = ( n11363 & n11733 ) | ( n11363 & ~n11734 ) | ( n11733 & ~n11734 ) ;
  assign n11736 = ( x112 & n11730 ) | ( x112 & ~n11735 ) | ( n11730 & ~n11735 ) ;
  assign n11737 = ( x112 & n11364 ) | ( x112 & ~n11450 ) | ( n11364 & ~n11450 ) ;
  assign n11738 = x112 & n11364 ;
  assign n11739 = ( ~n11369 & n11737 ) | ( ~n11369 & n11738 ) | ( n11737 & n11738 ) ;
  assign n11740 = ( n11369 & n11737 ) | ( n11369 & n11738 ) | ( n11737 & n11738 ) ;
  assign n11741 = ( n11369 & n11739 ) | ( n11369 & ~n11740 ) | ( n11739 & ~n11740 ) ;
  assign n11742 = ( x113 & n11736 ) | ( x113 & ~n11741 ) | ( n11736 & ~n11741 ) ;
  assign n11743 = ( x113 & n11370 ) | ( x113 & ~n11450 ) | ( n11370 & ~n11450 ) ;
  assign n11744 = x113 & n11370 ;
  assign n11745 = ( ~n11375 & n11743 ) | ( ~n11375 & n11744 ) | ( n11743 & n11744 ) ;
  assign n11746 = ( n11375 & n11743 ) | ( n11375 & n11744 ) | ( n11743 & n11744 ) ;
  assign n11747 = ( n11375 & n11745 ) | ( n11375 & ~n11746 ) | ( n11745 & ~n11746 ) ;
  assign n11748 = ( x114 & n11742 ) | ( x114 & ~n11747 ) | ( n11742 & ~n11747 ) ;
  assign n11749 = ( x114 & n11376 ) | ( x114 & ~n11450 ) | ( n11376 & ~n11450 ) ;
  assign n11750 = x114 & n11376 ;
  assign n11751 = ( ~n11381 & n11749 ) | ( ~n11381 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11752 = ( n11381 & n11749 ) | ( n11381 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11753 = ( n11381 & n11751 ) | ( n11381 & ~n11752 ) | ( n11751 & ~n11752 ) ;
  assign n11754 = ( x115 & n11748 ) | ( x115 & ~n11753 ) | ( n11748 & ~n11753 ) ;
  assign n11755 = ( x115 & n11382 ) | ( x115 & ~n11450 ) | ( n11382 & ~n11450 ) ;
  assign n11756 = x115 & n11382 ;
  assign n11757 = ( ~n11387 & n11755 ) | ( ~n11387 & n11756 ) | ( n11755 & n11756 ) ;
  assign n11758 = ( n11387 & n11755 ) | ( n11387 & n11756 ) | ( n11755 & n11756 ) ;
  assign n11759 = ( n11387 & n11757 ) | ( n11387 & ~n11758 ) | ( n11757 & ~n11758 ) ;
  assign n11760 = ( x116 & n11754 ) | ( x116 & ~n11759 ) | ( n11754 & ~n11759 ) ;
  assign n11761 = ( x116 & n11388 ) | ( x116 & ~n11450 ) | ( n11388 & ~n11450 ) ;
  assign n11762 = x116 & n11388 ;
  assign n11763 = ( ~n11393 & n11761 ) | ( ~n11393 & n11762 ) | ( n11761 & n11762 ) ;
  assign n11764 = ( n11393 & n11761 ) | ( n11393 & n11762 ) | ( n11761 & n11762 ) ;
  assign n11765 = ( n11393 & n11763 ) | ( n11393 & ~n11764 ) | ( n11763 & ~n11764 ) ;
  assign n11766 = ( x117 & n11760 ) | ( x117 & ~n11765 ) | ( n11760 & ~n11765 ) ;
  assign n11767 = ( x117 & n11394 ) | ( x117 & ~n11450 ) | ( n11394 & ~n11450 ) ;
  assign n11768 = x117 & n11394 ;
  assign n11769 = ( ~n11399 & n11767 ) | ( ~n11399 & n11768 ) | ( n11767 & n11768 ) ;
  assign n11770 = ( n11399 & n11767 ) | ( n11399 & n11768 ) | ( n11767 & n11768 ) ;
  assign n11771 = ( n11399 & n11769 ) | ( n11399 & ~n11770 ) | ( n11769 & ~n11770 ) ;
  assign n11772 = ( x118 & n11766 ) | ( x118 & ~n11771 ) | ( n11766 & ~n11771 ) ;
  assign n11773 = ( x118 & n11400 ) | ( x118 & ~n11450 ) | ( n11400 & ~n11450 ) ;
  assign n11774 = x118 & n11400 ;
  assign n11775 = ( ~n11405 & n11773 ) | ( ~n11405 & n11774 ) | ( n11773 & n11774 ) ;
  assign n11776 = ( n11405 & n11773 ) | ( n11405 & n11774 ) | ( n11773 & n11774 ) ;
  assign n11777 = ( n11405 & n11775 ) | ( n11405 & ~n11776 ) | ( n11775 & ~n11776 ) ;
  assign n11778 = ( x119 & n11772 ) | ( x119 & ~n11777 ) | ( n11772 & ~n11777 ) ;
  assign n11779 = ( x119 & n11406 ) | ( x119 & ~n11450 ) | ( n11406 & ~n11450 ) ;
  assign n11780 = x119 & n11406 ;
  assign n11781 = ( ~n11411 & n11779 ) | ( ~n11411 & n11780 ) | ( n11779 & n11780 ) ;
  assign n11782 = ( n11411 & n11779 ) | ( n11411 & n11780 ) | ( n11779 & n11780 ) ;
  assign n11783 = ( n11411 & n11781 ) | ( n11411 & ~n11782 ) | ( n11781 & ~n11782 ) ;
  assign n11784 = ( x120 & n11778 ) | ( x120 & ~n11783 ) | ( n11778 & ~n11783 ) ;
  assign n11785 = ( x120 & n11412 ) | ( x120 & ~n11450 ) | ( n11412 & ~n11450 ) ;
  assign n11786 = x120 & n11412 ;
  assign n11787 = ( ~n11417 & n11785 ) | ( ~n11417 & n11786 ) | ( n11785 & n11786 ) ;
  assign n11788 = ( n11417 & n11785 ) | ( n11417 & n11786 ) | ( n11785 & n11786 ) ;
  assign n11789 = ( n11417 & n11787 ) | ( n11417 & ~n11788 ) | ( n11787 & ~n11788 ) ;
  assign n11790 = ( x121 & n11784 ) | ( x121 & ~n11789 ) | ( n11784 & ~n11789 ) ;
  assign n11791 = ( x121 & n11418 ) | ( x121 & ~n11450 ) | ( n11418 & ~n11450 ) ;
  assign n11792 = x121 & n11418 ;
  assign n11793 = ( ~n11423 & n11791 ) | ( ~n11423 & n11792 ) | ( n11791 & n11792 ) ;
  assign n11794 = ( n11423 & n11791 ) | ( n11423 & n11792 ) | ( n11791 & n11792 ) ;
  assign n11795 = ( n11423 & n11793 ) | ( n11423 & ~n11794 ) | ( n11793 & ~n11794 ) ;
  assign n11796 = ( x122 & n11790 ) | ( x122 & ~n11795 ) | ( n11790 & ~n11795 ) ;
  assign n11797 = ( x122 & n11424 ) | ( x122 & ~n11450 ) | ( n11424 & ~n11450 ) ;
  assign n11798 = x122 & n11424 ;
  assign n11799 = ( ~n11429 & n11797 ) | ( ~n11429 & n11798 ) | ( n11797 & n11798 ) ;
  assign n11800 = ( n11429 & n11797 ) | ( n11429 & n11798 ) | ( n11797 & n11798 ) ;
  assign n11801 = ( n11429 & n11799 ) | ( n11429 & ~n11800 ) | ( n11799 & ~n11800 ) ;
  assign n11802 = ( x123 & n11796 ) | ( x123 & ~n11801 ) | ( n11796 & ~n11801 ) ;
  assign n11803 = ( x123 & n11430 ) | ( x123 & ~n11450 ) | ( n11430 & ~n11450 ) ;
  assign n11804 = x123 & n11430 ;
  assign n11805 = ( ~n11435 & n11803 ) | ( ~n11435 & n11804 ) | ( n11803 & n11804 ) ;
  assign n11806 = ( n11435 & n11803 ) | ( n11435 & n11804 ) | ( n11803 & n11804 ) ;
  assign n11807 = ( n11435 & n11805 ) | ( n11435 & ~n11806 ) | ( n11805 & ~n11806 ) ;
  assign n11808 = ( x124 & n11802 ) | ( x124 & ~n11807 ) | ( n11802 & ~n11807 ) ;
  assign n11809 = ( x124 & n11436 ) | ( x124 & ~n11450 ) | ( n11436 & ~n11450 ) ;
  assign n11810 = x124 & n11436 ;
  assign n11811 = ( ~n11441 & n11809 ) | ( ~n11441 & n11810 ) | ( n11809 & n11810 ) ;
  assign n11812 = ( n11441 & n11809 ) | ( n11441 & n11810 ) | ( n11809 & n11810 ) ;
  assign n11813 = ( n11441 & n11811 ) | ( n11441 & ~n11812 ) | ( n11811 & ~n11812 ) ;
  assign n11814 = ( x125 & n11808 ) | ( x125 & ~n11813 ) | ( n11808 & ~n11813 ) ;
  assign n11815 = x126 & n11446 ;
  assign n11816 = n389 | n11815 ;
  assign n11817 = ( n389 & n11814 ) | ( n389 & n11816 ) | ( n11814 & n11816 ) ;
  assign n11818 = ~x0 & x64 ;
  assign n11819 = ( x125 & ~n11442 ) | ( x125 & n11447 ) | ( ~n11442 & n11447 ) ;
  assign n11820 = x125 & ~n11442 ;
  assign n11821 = ( n11814 & ~n11819 ) | ( n11814 & n11820 ) | ( ~n11819 & n11820 ) ;
  assign n11822 = n131 & ~n11446 ;
  assign n11823 = n11821 | n11822 ;
  assign n11824 = ~x1 & n11823 ;
  assign n11825 = ( x1 & ~x64 ) | ( x1 & n11823 ) | ( ~x64 & n11823 ) ;
  assign n11826 = ( n390 & ~n11824 ) | ( n390 & n11825 ) | ( ~n11824 & n11825 ) ;
  assign n11827 = ( x65 & n11818 ) | ( x65 & ~n11826 ) | ( n11818 & ~n11826 ) ;
  assign n11828 = ( x65 & n390 ) | ( x65 & n11823 ) | ( n390 & n11823 ) ;
  assign n11829 = x65 | n390 ;
  assign n11830 = ( ~n11453 & n11828 ) | ( ~n11453 & n11829 ) | ( n11828 & n11829 ) ;
  assign n11831 = ( n11453 & n11828 ) | ( n11453 & n11829 ) | ( n11828 & n11829 ) ;
  assign n11832 = ( n11453 & n11830 ) | ( n11453 & ~n11831 ) | ( n11830 & ~n11831 ) ;
  assign n11833 = ( x66 & n11827 ) | ( x66 & ~n11832 ) | ( n11827 & ~n11832 ) ;
  assign n11834 = ( x66 & n11454 ) | ( x66 & n11823 ) | ( n11454 & n11823 ) ;
  assign n11835 = x66 | n11454 ;
  assign n11836 = ( ~n11459 & n11834 ) | ( ~n11459 & n11835 ) | ( n11834 & n11835 ) ;
  assign n11837 = ( n11459 & n11834 ) | ( n11459 & n11835 ) | ( n11834 & n11835 ) ;
  assign n11838 = ( n11459 & n11836 ) | ( n11459 & ~n11837 ) | ( n11836 & ~n11837 ) ;
  assign n11839 = ( x67 & n11833 ) | ( x67 & ~n11838 ) | ( n11833 & ~n11838 ) ;
  assign n11840 = ( x67 & n11460 ) | ( x67 & ~n11823 ) | ( n11460 & ~n11823 ) ;
  assign n11841 = x67 & n11460 ;
  assign n11842 = ( ~n11465 & n11840 ) | ( ~n11465 & n11841 ) | ( n11840 & n11841 ) ;
  assign n11843 = ( n11465 & n11840 ) | ( n11465 & n11841 ) | ( n11840 & n11841 ) ;
  assign n11844 = ( n11465 & n11842 ) | ( n11465 & ~n11843 ) | ( n11842 & ~n11843 ) ;
  assign n11845 = ( x68 & n11839 ) | ( x68 & ~n11844 ) | ( n11839 & ~n11844 ) ;
  assign n11846 = ( x68 & n11466 ) | ( x68 & ~n11823 ) | ( n11466 & ~n11823 ) ;
  assign n11847 = x68 & n11466 ;
  assign n11848 = ( ~n11471 & n11846 ) | ( ~n11471 & n11847 ) | ( n11846 & n11847 ) ;
  assign n11849 = ( n11471 & n11846 ) | ( n11471 & n11847 ) | ( n11846 & n11847 ) ;
  assign n11850 = ( n11471 & n11848 ) | ( n11471 & ~n11849 ) | ( n11848 & ~n11849 ) ;
  assign n11851 = ( x69 & n11845 ) | ( x69 & ~n11850 ) | ( n11845 & ~n11850 ) ;
  assign n11852 = ( x69 & n11472 ) | ( x69 & ~n11823 ) | ( n11472 & ~n11823 ) ;
  assign n11853 = x69 & n11472 ;
  assign n11854 = ( ~n11477 & n11852 ) | ( ~n11477 & n11853 ) | ( n11852 & n11853 ) ;
  assign n11855 = ( n11477 & n11852 ) | ( n11477 & n11853 ) | ( n11852 & n11853 ) ;
  assign n11856 = ( n11477 & n11854 ) | ( n11477 & ~n11855 ) | ( n11854 & ~n11855 ) ;
  assign n11857 = ( x70 & n11851 ) | ( x70 & ~n11856 ) | ( n11851 & ~n11856 ) ;
  assign n11858 = ( x70 & n11478 ) | ( x70 & ~n11823 ) | ( n11478 & ~n11823 ) ;
  assign n11859 = x70 & n11478 ;
  assign n11860 = ( ~n11483 & n11858 ) | ( ~n11483 & n11859 ) | ( n11858 & n11859 ) ;
  assign n11861 = ( n11483 & n11858 ) | ( n11483 & n11859 ) | ( n11858 & n11859 ) ;
  assign n11862 = ( n11483 & n11860 ) | ( n11483 & ~n11861 ) | ( n11860 & ~n11861 ) ;
  assign n11863 = ( x71 & n11857 ) | ( x71 & ~n11862 ) | ( n11857 & ~n11862 ) ;
  assign n11864 = ( x71 & n11484 ) | ( x71 & ~n11823 ) | ( n11484 & ~n11823 ) ;
  assign n11865 = x71 & n11484 ;
  assign n11866 = ( ~n11489 & n11864 ) | ( ~n11489 & n11865 ) | ( n11864 & n11865 ) ;
  assign n11867 = ( n11489 & n11864 ) | ( n11489 & n11865 ) | ( n11864 & n11865 ) ;
  assign n11868 = ( n11489 & n11866 ) | ( n11489 & ~n11867 ) | ( n11866 & ~n11867 ) ;
  assign n11869 = ( x72 & n11863 ) | ( x72 & ~n11868 ) | ( n11863 & ~n11868 ) ;
  assign n11870 = ( x72 & n11490 ) | ( x72 & ~n11823 ) | ( n11490 & ~n11823 ) ;
  assign n11871 = x72 & n11490 ;
  assign n11872 = ( ~n11495 & n11870 ) | ( ~n11495 & n11871 ) | ( n11870 & n11871 ) ;
  assign n11873 = ( n11495 & n11870 ) | ( n11495 & n11871 ) | ( n11870 & n11871 ) ;
  assign n11874 = ( n11495 & n11872 ) | ( n11495 & ~n11873 ) | ( n11872 & ~n11873 ) ;
  assign n11875 = ( x73 & n11869 ) | ( x73 & ~n11874 ) | ( n11869 & ~n11874 ) ;
  assign n11876 = ( x73 & n11496 ) | ( x73 & ~n11823 ) | ( n11496 & ~n11823 ) ;
  assign n11877 = x73 & n11496 ;
  assign n11878 = ( ~n11501 & n11876 ) | ( ~n11501 & n11877 ) | ( n11876 & n11877 ) ;
  assign n11879 = ( n11501 & n11876 ) | ( n11501 & n11877 ) | ( n11876 & n11877 ) ;
  assign n11880 = ( n11501 & n11878 ) | ( n11501 & ~n11879 ) | ( n11878 & ~n11879 ) ;
  assign n11881 = ( x74 & n11875 ) | ( x74 & ~n11880 ) | ( n11875 & ~n11880 ) ;
  assign n11882 = ( x74 & n11502 ) | ( x74 & ~n11823 ) | ( n11502 & ~n11823 ) ;
  assign n11883 = x74 & n11502 ;
  assign n11884 = ( ~n11507 & n11882 ) | ( ~n11507 & n11883 ) | ( n11882 & n11883 ) ;
  assign n11885 = ( n11507 & n11882 ) | ( n11507 & n11883 ) | ( n11882 & n11883 ) ;
  assign n11886 = ( n11507 & n11884 ) | ( n11507 & ~n11885 ) | ( n11884 & ~n11885 ) ;
  assign n11887 = ( x75 & n11881 ) | ( x75 & ~n11886 ) | ( n11881 & ~n11886 ) ;
  assign n11888 = ( x75 & n11508 ) | ( x75 & ~n11823 ) | ( n11508 & ~n11823 ) ;
  assign n11889 = x75 & n11508 ;
  assign n11890 = ( ~n11513 & n11888 ) | ( ~n11513 & n11889 ) | ( n11888 & n11889 ) ;
  assign n11891 = ( n11513 & n11888 ) | ( n11513 & n11889 ) | ( n11888 & n11889 ) ;
  assign n11892 = ( n11513 & n11890 ) | ( n11513 & ~n11891 ) | ( n11890 & ~n11891 ) ;
  assign n11893 = ( x76 & n11887 ) | ( x76 & ~n11892 ) | ( n11887 & ~n11892 ) ;
  assign n11894 = ( x76 & n11514 ) | ( x76 & ~n11823 ) | ( n11514 & ~n11823 ) ;
  assign n11895 = x76 & n11514 ;
  assign n11896 = ( ~n11519 & n11894 ) | ( ~n11519 & n11895 ) | ( n11894 & n11895 ) ;
  assign n11897 = ( n11519 & n11894 ) | ( n11519 & n11895 ) | ( n11894 & n11895 ) ;
  assign n11898 = ( n11519 & n11896 ) | ( n11519 & ~n11897 ) | ( n11896 & ~n11897 ) ;
  assign n11899 = ( x77 & n11893 ) | ( x77 & ~n11898 ) | ( n11893 & ~n11898 ) ;
  assign n11900 = ( x77 & n11520 ) | ( x77 & ~n11823 ) | ( n11520 & ~n11823 ) ;
  assign n11901 = x77 & n11520 ;
  assign n11902 = ( ~n11525 & n11900 ) | ( ~n11525 & n11901 ) | ( n11900 & n11901 ) ;
  assign n11903 = ( n11525 & n11900 ) | ( n11525 & n11901 ) | ( n11900 & n11901 ) ;
  assign n11904 = ( n11525 & n11902 ) | ( n11525 & ~n11903 ) | ( n11902 & ~n11903 ) ;
  assign n11905 = ( x78 & n11899 ) | ( x78 & ~n11904 ) | ( n11899 & ~n11904 ) ;
  assign n11906 = ( x78 & n11526 ) | ( x78 & ~n11823 ) | ( n11526 & ~n11823 ) ;
  assign n11907 = x78 & n11526 ;
  assign n11908 = ( ~n11531 & n11906 ) | ( ~n11531 & n11907 ) | ( n11906 & n11907 ) ;
  assign n11909 = ( n11531 & n11906 ) | ( n11531 & n11907 ) | ( n11906 & n11907 ) ;
  assign n11910 = ( n11531 & n11908 ) | ( n11531 & ~n11909 ) | ( n11908 & ~n11909 ) ;
  assign n11911 = ( x79 & n11905 ) | ( x79 & ~n11910 ) | ( n11905 & ~n11910 ) ;
  assign n11912 = ( x79 & n11532 ) | ( x79 & ~n11823 ) | ( n11532 & ~n11823 ) ;
  assign n11913 = x79 & n11532 ;
  assign n11914 = ( ~n11537 & n11912 ) | ( ~n11537 & n11913 ) | ( n11912 & n11913 ) ;
  assign n11915 = ( n11537 & n11912 ) | ( n11537 & n11913 ) | ( n11912 & n11913 ) ;
  assign n11916 = ( n11537 & n11914 ) | ( n11537 & ~n11915 ) | ( n11914 & ~n11915 ) ;
  assign n11917 = ( x80 & n11911 ) | ( x80 & ~n11916 ) | ( n11911 & ~n11916 ) ;
  assign n11918 = ( x80 & n11538 ) | ( x80 & ~n11823 ) | ( n11538 & ~n11823 ) ;
  assign n11919 = x80 & n11538 ;
  assign n11920 = ( ~n11543 & n11918 ) | ( ~n11543 & n11919 ) | ( n11918 & n11919 ) ;
  assign n11921 = ( n11543 & n11918 ) | ( n11543 & n11919 ) | ( n11918 & n11919 ) ;
  assign n11922 = ( n11543 & n11920 ) | ( n11543 & ~n11921 ) | ( n11920 & ~n11921 ) ;
  assign n11923 = ( x81 & n11917 ) | ( x81 & ~n11922 ) | ( n11917 & ~n11922 ) ;
  assign n11924 = ( x81 & n11544 ) | ( x81 & ~n11823 ) | ( n11544 & ~n11823 ) ;
  assign n11925 = x81 & n11544 ;
  assign n11926 = ( ~n11549 & n11924 ) | ( ~n11549 & n11925 ) | ( n11924 & n11925 ) ;
  assign n11927 = ( n11549 & n11924 ) | ( n11549 & n11925 ) | ( n11924 & n11925 ) ;
  assign n11928 = ( n11549 & n11926 ) | ( n11549 & ~n11927 ) | ( n11926 & ~n11927 ) ;
  assign n11929 = ( x82 & n11923 ) | ( x82 & ~n11928 ) | ( n11923 & ~n11928 ) ;
  assign n11930 = ( x82 & n11550 ) | ( x82 & ~n11823 ) | ( n11550 & ~n11823 ) ;
  assign n11931 = x82 & n11550 ;
  assign n11932 = ( ~n11555 & n11930 ) | ( ~n11555 & n11931 ) | ( n11930 & n11931 ) ;
  assign n11933 = ( n11555 & n11930 ) | ( n11555 & n11931 ) | ( n11930 & n11931 ) ;
  assign n11934 = ( n11555 & n11932 ) | ( n11555 & ~n11933 ) | ( n11932 & ~n11933 ) ;
  assign n11935 = ( x83 & n11929 ) | ( x83 & ~n11934 ) | ( n11929 & ~n11934 ) ;
  assign n11936 = ( x83 & n11556 ) | ( x83 & ~n11823 ) | ( n11556 & ~n11823 ) ;
  assign n11937 = x83 & n11556 ;
  assign n11938 = ( ~n11561 & n11936 ) | ( ~n11561 & n11937 ) | ( n11936 & n11937 ) ;
  assign n11939 = ( n11561 & n11936 ) | ( n11561 & n11937 ) | ( n11936 & n11937 ) ;
  assign n11940 = ( n11561 & n11938 ) | ( n11561 & ~n11939 ) | ( n11938 & ~n11939 ) ;
  assign n11941 = ( x84 & n11935 ) | ( x84 & ~n11940 ) | ( n11935 & ~n11940 ) ;
  assign n11942 = ( x84 & n11562 ) | ( x84 & ~n11823 ) | ( n11562 & ~n11823 ) ;
  assign n11943 = x84 & n11562 ;
  assign n11944 = ( ~n11567 & n11942 ) | ( ~n11567 & n11943 ) | ( n11942 & n11943 ) ;
  assign n11945 = ( n11567 & n11942 ) | ( n11567 & n11943 ) | ( n11942 & n11943 ) ;
  assign n11946 = ( n11567 & n11944 ) | ( n11567 & ~n11945 ) | ( n11944 & ~n11945 ) ;
  assign n11947 = ( x85 & n11941 ) | ( x85 & ~n11946 ) | ( n11941 & ~n11946 ) ;
  assign n11948 = ( x85 & n11568 ) | ( x85 & ~n11823 ) | ( n11568 & ~n11823 ) ;
  assign n11949 = x85 & n11568 ;
  assign n11950 = ( ~n11573 & n11948 ) | ( ~n11573 & n11949 ) | ( n11948 & n11949 ) ;
  assign n11951 = ( n11573 & n11948 ) | ( n11573 & n11949 ) | ( n11948 & n11949 ) ;
  assign n11952 = ( n11573 & n11950 ) | ( n11573 & ~n11951 ) | ( n11950 & ~n11951 ) ;
  assign n11953 = ( x86 & n11947 ) | ( x86 & ~n11952 ) | ( n11947 & ~n11952 ) ;
  assign n11954 = ( x86 & n11574 ) | ( x86 & ~n11823 ) | ( n11574 & ~n11823 ) ;
  assign n11955 = x86 & n11574 ;
  assign n11956 = ( ~n11579 & n11954 ) | ( ~n11579 & n11955 ) | ( n11954 & n11955 ) ;
  assign n11957 = ( n11579 & n11954 ) | ( n11579 & n11955 ) | ( n11954 & n11955 ) ;
  assign n11958 = ( n11579 & n11956 ) | ( n11579 & ~n11957 ) | ( n11956 & ~n11957 ) ;
  assign n11959 = ( x87 & n11953 ) | ( x87 & ~n11958 ) | ( n11953 & ~n11958 ) ;
  assign n11960 = ( x87 & n11580 ) | ( x87 & ~n11823 ) | ( n11580 & ~n11823 ) ;
  assign n11961 = x87 & n11580 ;
  assign n11962 = ( ~n11585 & n11960 ) | ( ~n11585 & n11961 ) | ( n11960 & n11961 ) ;
  assign n11963 = ( n11585 & n11960 ) | ( n11585 & n11961 ) | ( n11960 & n11961 ) ;
  assign n11964 = ( n11585 & n11962 ) | ( n11585 & ~n11963 ) | ( n11962 & ~n11963 ) ;
  assign n11965 = ( x88 & n11959 ) | ( x88 & ~n11964 ) | ( n11959 & ~n11964 ) ;
  assign n11966 = ( x88 & n11586 ) | ( x88 & ~n11823 ) | ( n11586 & ~n11823 ) ;
  assign n11967 = x88 & n11586 ;
  assign n11968 = ( ~n11591 & n11966 ) | ( ~n11591 & n11967 ) | ( n11966 & n11967 ) ;
  assign n11969 = ( n11591 & n11966 ) | ( n11591 & n11967 ) | ( n11966 & n11967 ) ;
  assign n11970 = ( n11591 & n11968 ) | ( n11591 & ~n11969 ) | ( n11968 & ~n11969 ) ;
  assign n11971 = ( x89 & n11965 ) | ( x89 & ~n11970 ) | ( n11965 & ~n11970 ) ;
  assign n11972 = ( x89 & n11592 ) | ( x89 & ~n11823 ) | ( n11592 & ~n11823 ) ;
  assign n11973 = x89 & n11592 ;
  assign n11974 = ( ~n11597 & n11972 ) | ( ~n11597 & n11973 ) | ( n11972 & n11973 ) ;
  assign n11975 = ( n11597 & n11972 ) | ( n11597 & n11973 ) | ( n11972 & n11973 ) ;
  assign n11976 = ( n11597 & n11974 ) | ( n11597 & ~n11975 ) | ( n11974 & ~n11975 ) ;
  assign n11977 = ( x90 & n11971 ) | ( x90 & ~n11976 ) | ( n11971 & ~n11976 ) ;
  assign n11978 = ( x90 & n11598 ) | ( x90 & ~n11823 ) | ( n11598 & ~n11823 ) ;
  assign n11979 = x90 & n11598 ;
  assign n11980 = ( ~n11603 & n11978 ) | ( ~n11603 & n11979 ) | ( n11978 & n11979 ) ;
  assign n11981 = ( n11603 & n11978 ) | ( n11603 & n11979 ) | ( n11978 & n11979 ) ;
  assign n11982 = ( n11603 & n11980 ) | ( n11603 & ~n11981 ) | ( n11980 & ~n11981 ) ;
  assign n11983 = ( x91 & n11977 ) | ( x91 & ~n11982 ) | ( n11977 & ~n11982 ) ;
  assign n11984 = ( x91 & n11604 ) | ( x91 & ~n11823 ) | ( n11604 & ~n11823 ) ;
  assign n11985 = x91 & n11604 ;
  assign n11986 = ( ~n11609 & n11984 ) | ( ~n11609 & n11985 ) | ( n11984 & n11985 ) ;
  assign n11987 = ( n11609 & n11984 ) | ( n11609 & n11985 ) | ( n11984 & n11985 ) ;
  assign n11988 = ( n11609 & n11986 ) | ( n11609 & ~n11987 ) | ( n11986 & ~n11987 ) ;
  assign n11989 = ( x92 & n11983 ) | ( x92 & ~n11988 ) | ( n11983 & ~n11988 ) ;
  assign n11990 = ( x92 & n11610 ) | ( x92 & ~n11823 ) | ( n11610 & ~n11823 ) ;
  assign n11991 = x92 & n11610 ;
  assign n11992 = ( ~n11615 & n11990 ) | ( ~n11615 & n11991 ) | ( n11990 & n11991 ) ;
  assign n11993 = ( n11615 & n11990 ) | ( n11615 & n11991 ) | ( n11990 & n11991 ) ;
  assign n11994 = ( n11615 & n11992 ) | ( n11615 & ~n11993 ) | ( n11992 & ~n11993 ) ;
  assign n11995 = ( x93 & n11989 ) | ( x93 & ~n11994 ) | ( n11989 & ~n11994 ) ;
  assign n11996 = ( x93 & n11616 ) | ( x93 & ~n11823 ) | ( n11616 & ~n11823 ) ;
  assign n11997 = x93 & n11616 ;
  assign n11998 = ( ~n11621 & n11996 ) | ( ~n11621 & n11997 ) | ( n11996 & n11997 ) ;
  assign n11999 = ( n11621 & n11996 ) | ( n11621 & n11997 ) | ( n11996 & n11997 ) ;
  assign n12000 = ( n11621 & n11998 ) | ( n11621 & ~n11999 ) | ( n11998 & ~n11999 ) ;
  assign n12001 = ( x94 & n11995 ) | ( x94 & ~n12000 ) | ( n11995 & ~n12000 ) ;
  assign n12002 = ( x94 & n11622 ) | ( x94 & ~n11823 ) | ( n11622 & ~n11823 ) ;
  assign n12003 = x94 & n11622 ;
  assign n12004 = ( ~n11627 & n12002 ) | ( ~n11627 & n12003 ) | ( n12002 & n12003 ) ;
  assign n12005 = ( n11627 & n12002 ) | ( n11627 & n12003 ) | ( n12002 & n12003 ) ;
  assign n12006 = ( n11627 & n12004 ) | ( n11627 & ~n12005 ) | ( n12004 & ~n12005 ) ;
  assign n12007 = ( x95 & n12001 ) | ( x95 & ~n12006 ) | ( n12001 & ~n12006 ) ;
  assign n12008 = ( x95 & n11628 ) | ( x95 & ~n11823 ) | ( n11628 & ~n11823 ) ;
  assign n12009 = x95 & n11628 ;
  assign n12010 = ( ~n11633 & n12008 ) | ( ~n11633 & n12009 ) | ( n12008 & n12009 ) ;
  assign n12011 = ( n11633 & n12008 ) | ( n11633 & n12009 ) | ( n12008 & n12009 ) ;
  assign n12012 = ( n11633 & n12010 ) | ( n11633 & ~n12011 ) | ( n12010 & ~n12011 ) ;
  assign n12013 = ( x96 & n12007 ) | ( x96 & ~n12012 ) | ( n12007 & ~n12012 ) ;
  assign n12014 = ( x96 & n11634 ) | ( x96 & ~n11823 ) | ( n11634 & ~n11823 ) ;
  assign n12015 = x96 & n11634 ;
  assign n12016 = ( ~n11639 & n12014 ) | ( ~n11639 & n12015 ) | ( n12014 & n12015 ) ;
  assign n12017 = ( n11639 & n12014 ) | ( n11639 & n12015 ) | ( n12014 & n12015 ) ;
  assign n12018 = ( n11639 & n12016 ) | ( n11639 & ~n12017 ) | ( n12016 & ~n12017 ) ;
  assign n12019 = ( x97 & n12013 ) | ( x97 & ~n12018 ) | ( n12013 & ~n12018 ) ;
  assign n12020 = ( x97 & n11640 ) | ( x97 & ~n11823 ) | ( n11640 & ~n11823 ) ;
  assign n12021 = x97 & n11640 ;
  assign n12022 = ( ~n11645 & n12020 ) | ( ~n11645 & n12021 ) | ( n12020 & n12021 ) ;
  assign n12023 = ( n11645 & n12020 ) | ( n11645 & n12021 ) | ( n12020 & n12021 ) ;
  assign n12024 = ( n11645 & n12022 ) | ( n11645 & ~n12023 ) | ( n12022 & ~n12023 ) ;
  assign n12025 = ( x98 & n12019 ) | ( x98 & ~n12024 ) | ( n12019 & ~n12024 ) ;
  assign n12026 = ( x98 & n11646 ) | ( x98 & ~n11823 ) | ( n11646 & ~n11823 ) ;
  assign n12027 = x98 & n11646 ;
  assign n12028 = ( ~n11651 & n12026 ) | ( ~n11651 & n12027 ) | ( n12026 & n12027 ) ;
  assign n12029 = ( n11651 & n12026 ) | ( n11651 & n12027 ) | ( n12026 & n12027 ) ;
  assign n12030 = ( n11651 & n12028 ) | ( n11651 & ~n12029 ) | ( n12028 & ~n12029 ) ;
  assign n12031 = ( x99 & n12025 ) | ( x99 & ~n12030 ) | ( n12025 & ~n12030 ) ;
  assign n12032 = ( x99 & n11652 ) | ( x99 & ~n11823 ) | ( n11652 & ~n11823 ) ;
  assign n12033 = x99 & n11652 ;
  assign n12034 = ( ~n11657 & n12032 ) | ( ~n11657 & n12033 ) | ( n12032 & n12033 ) ;
  assign n12035 = ( n11657 & n12032 ) | ( n11657 & n12033 ) | ( n12032 & n12033 ) ;
  assign n12036 = ( n11657 & n12034 ) | ( n11657 & ~n12035 ) | ( n12034 & ~n12035 ) ;
  assign n12037 = ( x100 & n12031 ) | ( x100 & ~n12036 ) | ( n12031 & ~n12036 ) ;
  assign n12038 = ( x100 & n11658 ) | ( x100 & ~n11823 ) | ( n11658 & ~n11823 ) ;
  assign n12039 = x100 & n11658 ;
  assign n12040 = ( ~n11663 & n12038 ) | ( ~n11663 & n12039 ) | ( n12038 & n12039 ) ;
  assign n12041 = ( n11663 & n12038 ) | ( n11663 & n12039 ) | ( n12038 & n12039 ) ;
  assign n12042 = ( n11663 & n12040 ) | ( n11663 & ~n12041 ) | ( n12040 & ~n12041 ) ;
  assign n12043 = ( x101 & n12037 ) | ( x101 & ~n12042 ) | ( n12037 & ~n12042 ) ;
  assign n12044 = ( x101 & n11664 ) | ( x101 & ~n11823 ) | ( n11664 & ~n11823 ) ;
  assign n12045 = x101 & n11664 ;
  assign n12046 = ( ~n11669 & n12044 ) | ( ~n11669 & n12045 ) | ( n12044 & n12045 ) ;
  assign n12047 = ( n11669 & n12044 ) | ( n11669 & n12045 ) | ( n12044 & n12045 ) ;
  assign n12048 = ( n11669 & n12046 ) | ( n11669 & ~n12047 ) | ( n12046 & ~n12047 ) ;
  assign n12049 = ( x102 & n12043 ) | ( x102 & ~n12048 ) | ( n12043 & ~n12048 ) ;
  assign n12050 = ( x102 & n11670 ) | ( x102 & ~n11823 ) | ( n11670 & ~n11823 ) ;
  assign n12051 = x102 & n11670 ;
  assign n12052 = ( ~n11675 & n12050 ) | ( ~n11675 & n12051 ) | ( n12050 & n12051 ) ;
  assign n12053 = ( n11675 & n12050 ) | ( n11675 & n12051 ) | ( n12050 & n12051 ) ;
  assign n12054 = ( n11675 & n12052 ) | ( n11675 & ~n12053 ) | ( n12052 & ~n12053 ) ;
  assign n12055 = ( x103 & n12049 ) | ( x103 & ~n12054 ) | ( n12049 & ~n12054 ) ;
  assign n12056 = ( x103 & n11676 ) | ( x103 & ~n11823 ) | ( n11676 & ~n11823 ) ;
  assign n12057 = x103 & n11676 ;
  assign n12058 = ( ~n11681 & n12056 ) | ( ~n11681 & n12057 ) | ( n12056 & n12057 ) ;
  assign n12059 = ( n11681 & n12056 ) | ( n11681 & n12057 ) | ( n12056 & n12057 ) ;
  assign n12060 = ( n11681 & n12058 ) | ( n11681 & ~n12059 ) | ( n12058 & ~n12059 ) ;
  assign n12061 = ( x104 & n12055 ) | ( x104 & ~n12060 ) | ( n12055 & ~n12060 ) ;
  assign n12062 = ( x104 & n11682 ) | ( x104 & ~n11823 ) | ( n11682 & ~n11823 ) ;
  assign n12063 = x104 & n11682 ;
  assign n12064 = ( ~n11687 & n12062 ) | ( ~n11687 & n12063 ) | ( n12062 & n12063 ) ;
  assign n12065 = ( n11687 & n12062 ) | ( n11687 & n12063 ) | ( n12062 & n12063 ) ;
  assign n12066 = ( n11687 & n12064 ) | ( n11687 & ~n12065 ) | ( n12064 & ~n12065 ) ;
  assign n12067 = ( x105 & n12061 ) | ( x105 & ~n12066 ) | ( n12061 & ~n12066 ) ;
  assign n12068 = ( x105 & n11688 ) | ( x105 & ~n11823 ) | ( n11688 & ~n11823 ) ;
  assign n12069 = x105 & n11688 ;
  assign n12070 = ( ~n11693 & n12068 ) | ( ~n11693 & n12069 ) | ( n12068 & n12069 ) ;
  assign n12071 = ( n11693 & n12068 ) | ( n11693 & n12069 ) | ( n12068 & n12069 ) ;
  assign n12072 = ( n11693 & n12070 ) | ( n11693 & ~n12071 ) | ( n12070 & ~n12071 ) ;
  assign n12073 = ( x106 & n12067 ) | ( x106 & ~n12072 ) | ( n12067 & ~n12072 ) ;
  assign n12074 = ( x106 & n11694 ) | ( x106 & ~n11823 ) | ( n11694 & ~n11823 ) ;
  assign n12075 = x106 & n11694 ;
  assign n12076 = ( ~n11699 & n12074 ) | ( ~n11699 & n12075 ) | ( n12074 & n12075 ) ;
  assign n12077 = ( n11699 & n12074 ) | ( n11699 & n12075 ) | ( n12074 & n12075 ) ;
  assign n12078 = ( n11699 & n12076 ) | ( n11699 & ~n12077 ) | ( n12076 & ~n12077 ) ;
  assign n12079 = ( x107 & n12073 ) | ( x107 & ~n12078 ) | ( n12073 & ~n12078 ) ;
  assign n12080 = ( x107 & n11700 ) | ( x107 & ~n11823 ) | ( n11700 & ~n11823 ) ;
  assign n12081 = x107 & n11700 ;
  assign n12082 = ( ~n11705 & n12080 ) | ( ~n11705 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12083 = ( n11705 & n12080 ) | ( n11705 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12084 = ( n11705 & n12082 ) | ( n11705 & ~n12083 ) | ( n12082 & ~n12083 ) ;
  assign n12085 = ( x108 & n12079 ) | ( x108 & ~n12084 ) | ( n12079 & ~n12084 ) ;
  assign n12086 = ( x108 & n11706 ) | ( x108 & ~n11823 ) | ( n11706 & ~n11823 ) ;
  assign n12087 = x108 & n11706 ;
  assign n12088 = ( ~n11711 & n12086 ) | ( ~n11711 & n12087 ) | ( n12086 & n12087 ) ;
  assign n12089 = ( n11711 & n12086 ) | ( n11711 & n12087 ) | ( n12086 & n12087 ) ;
  assign n12090 = ( n11711 & n12088 ) | ( n11711 & ~n12089 ) | ( n12088 & ~n12089 ) ;
  assign n12091 = ( x109 & n12085 ) | ( x109 & ~n12090 ) | ( n12085 & ~n12090 ) ;
  assign n12092 = ( x109 & n11712 ) | ( x109 & ~n11823 ) | ( n11712 & ~n11823 ) ;
  assign n12093 = x109 & n11712 ;
  assign n12094 = ( ~n11717 & n12092 ) | ( ~n11717 & n12093 ) | ( n12092 & n12093 ) ;
  assign n12095 = ( n11717 & n12092 ) | ( n11717 & n12093 ) | ( n12092 & n12093 ) ;
  assign n12096 = ( n11717 & n12094 ) | ( n11717 & ~n12095 ) | ( n12094 & ~n12095 ) ;
  assign n12097 = ( x110 & n12091 ) | ( x110 & ~n12096 ) | ( n12091 & ~n12096 ) ;
  assign n12098 = ( x110 & n11718 ) | ( x110 & ~n11823 ) | ( n11718 & ~n11823 ) ;
  assign n12099 = x110 & n11718 ;
  assign n12100 = ( ~n11723 & n12098 ) | ( ~n11723 & n12099 ) | ( n12098 & n12099 ) ;
  assign n12101 = ( n11723 & n12098 ) | ( n11723 & n12099 ) | ( n12098 & n12099 ) ;
  assign n12102 = ( n11723 & n12100 ) | ( n11723 & ~n12101 ) | ( n12100 & ~n12101 ) ;
  assign n12103 = ( x111 & n12097 ) | ( x111 & ~n12102 ) | ( n12097 & ~n12102 ) ;
  assign n12104 = ( x111 & n11724 ) | ( x111 & ~n11823 ) | ( n11724 & ~n11823 ) ;
  assign n12105 = x111 & n11724 ;
  assign n12106 = ( ~n11729 & n12104 ) | ( ~n11729 & n12105 ) | ( n12104 & n12105 ) ;
  assign n12107 = ( n11729 & n12104 ) | ( n11729 & n12105 ) | ( n12104 & n12105 ) ;
  assign n12108 = ( n11729 & n12106 ) | ( n11729 & ~n12107 ) | ( n12106 & ~n12107 ) ;
  assign n12109 = ( x112 & n12103 ) | ( x112 & ~n12108 ) | ( n12103 & ~n12108 ) ;
  assign n12110 = ( x112 & n11730 ) | ( x112 & ~n11823 ) | ( n11730 & ~n11823 ) ;
  assign n12111 = x112 & n11730 ;
  assign n12112 = ( ~n11735 & n12110 ) | ( ~n11735 & n12111 ) | ( n12110 & n12111 ) ;
  assign n12113 = ( n11735 & n12110 ) | ( n11735 & n12111 ) | ( n12110 & n12111 ) ;
  assign n12114 = ( n11735 & n12112 ) | ( n11735 & ~n12113 ) | ( n12112 & ~n12113 ) ;
  assign n12115 = ( x113 & n12109 ) | ( x113 & ~n12114 ) | ( n12109 & ~n12114 ) ;
  assign n12116 = ( x113 & n11736 ) | ( x113 & ~n11823 ) | ( n11736 & ~n11823 ) ;
  assign n12117 = x113 & n11736 ;
  assign n12118 = ( ~n11741 & n12116 ) | ( ~n11741 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12119 = ( n11741 & n12116 ) | ( n11741 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12120 = ( n11741 & n12118 ) | ( n11741 & ~n12119 ) | ( n12118 & ~n12119 ) ;
  assign n12121 = ( x114 & n12115 ) | ( x114 & ~n12120 ) | ( n12115 & ~n12120 ) ;
  assign n12122 = ( x114 & n11742 ) | ( x114 & ~n11823 ) | ( n11742 & ~n11823 ) ;
  assign n12123 = x114 & n11742 ;
  assign n12124 = ( ~n11747 & n12122 ) | ( ~n11747 & n12123 ) | ( n12122 & n12123 ) ;
  assign n12125 = ( n11747 & n12122 ) | ( n11747 & n12123 ) | ( n12122 & n12123 ) ;
  assign n12126 = ( n11747 & n12124 ) | ( n11747 & ~n12125 ) | ( n12124 & ~n12125 ) ;
  assign n12127 = ( x115 & n12121 ) | ( x115 & ~n12126 ) | ( n12121 & ~n12126 ) ;
  assign n12128 = ( x115 & n11748 ) | ( x115 & ~n11823 ) | ( n11748 & ~n11823 ) ;
  assign n12129 = x115 & n11748 ;
  assign n12130 = ( ~n11753 & n12128 ) | ( ~n11753 & n12129 ) | ( n12128 & n12129 ) ;
  assign n12131 = ( n11753 & n12128 ) | ( n11753 & n12129 ) | ( n12128 & n12129 ) ;
  assign n12132 = ( n11753 & n12130 ) | ( n11753 & ~n12131 ) | ( n12130 & ~n12131 ) ;
  assign n12133 = ( x116 & n12127 ) | ( x116 & ~n12132 ) | ( n12127 & ~n12132 ) ;
  assign n12134 = ( x116 & n11754 ) | ( x116 & ~n11823 ) | ( n11754 & ~n11823 ) ;
  assign n12135 = x116 & n11754 ;
  assign n12136 = ( ~n11759 & n12134 ) | ( ~n11759 & n12135 ) | ( n12134 & n12135 ) ;
  assign n12137 = ( n11759 & n12134 ) | ( n11759 & n12135 ) | ( n12134 & n12135 ) ;
  assign n12138 = ( n11759 & n12136 ) | ( n11759 & ~n12137 ) | ( n12136 & ~n12137 ) ;
  assign n12139 = ( x117 & n12133 ) | ( x117 & ~n12138 ) | ( n12133 & ~n12138 ) ;
  assign n12140 = ( x117 & n11760 ) | ( x117 & ~n11823 ) | ( n11760 & ~n11823 ) ;
  assign n12141 = x117 & n11760 ;
  assign n12142 = ( ~n11765 & n12140 ) | ( ~n11765 & n12141 ) | ( n12140 & n12141 ) ;
  assign n12143 = ( n11765 & n12140 ) | ( n11765 & n12141 ) | ( n12140 & n12141 ) ;
  assign n12144 = ( n11765 & n12142 ) | ( n11765 & ~n12143 ) | ( n12142 & ~n12143 ) ;
  assign n12145 = ( x118 & n12139 ) | ( x118 & ~n12144 ) | ( n12139 & ~n12144 ) ;
  assign n12146 = ( x118 & n11766 ) | ( x118 & ~n11823 ) | ( n11766 & ~n11823 ) ;
  assign n12147 = x118 & n11766 ;
  assign n12148 = ( ~n11771 & n12146 ) | ( ~n11771 & n12147 ) | ( n12146 & n12147 ) ;
  assign n12149 = ( n11771 & n12146 ) | ( n11771 & n12147 ) | ( n12146 & n12147 ) ;
  assign n12150 = ( n11771 & n12148 ) | ( n11771 & ~n12149 ) | ( n12148 & ~n12149 ) ;
  assign n12151 = ( x119 & n12145 ) | ( x119 & ~n12150 ) | ( n12145 & ~n12150 ) ;
  assign n12152 = ( x119 & n11772 ) | ( x119 & ~n11823 ) | ( n11772 & ~n11823 ) ;
  assign n12153 = x119 & n11772 ;
  assign n12154 = ( ~n11777 & n12152 ) | ( ~n11777 & n12153 ) | ( n12152 & n12153 ) ;
  assign n12155 = ( n11777 & n12152 ) | ( n11777 & n12153 ) | ( n12152 & n12153 ) ;
  assign n12156 = ( n11777 & n12154 ) | ( n11777 & ~n12155 ) | ( n12154 & ~n12155 ) ;
  assign n12157 = ( x120 & n12151 ) | ( x120 & ~n12156 ) | ( n12151 & ~n12156 ) ;
  assign n12158 = ( x120 & n11778 ) | ( x120 & ~n11823 ) | ( n11778 & ~n11823 ) ;
  assign n12159 = x120 & n11778 ;
  assign n12160 = ( ~n11783 & n12158 ) | ( ~n11783 & n12159 ) | ( n12158 & n12159 ) ;
  assign n12161 = ( n11783 & n12158 ) | ( n11783 & n12159 ) | ( n12158 & n12159 ) ;
  assign n12162 = ( n11783 & n12160 ) | ( n11783 & ~n12161 ) | ( n12160 & ~n12161 ) ;
  assign n12163 = ( x121 & n12157 ) | ( x121 & ~n12162 ) | ( n12157 & ~n12162 ) ;
  assign n12164 = ( x121 & n11784 ) | ( x121 & ~n11823 ) | ( n11784 & ~n11823 ) ;
  assign n12165 = x121 & n11784 ;
  assign n12166 = ( ~n11789 & n12164 ) | ( ~n11789 & n12165 ) | ( n12164 & n12165 ) ;
  assign n12167 = ( n11789 & n12164 ) | ( n11789 & n12165 ) | ( n12164 & n12165 ) ;
  assign n12168 = ( n11789 & n12166 ) | ( n11789 & ~n12167 ) | ( n12166 & ~n12167 ) ;
  assign n12169 = ( x122 & n12163 ) | ( x122 & ~n12168 ) | ( n12163 & ~n12168 ) ;
  assign n12170 = ( x122 & n11790 ) | ( x122 & ~n11823 ) | ( n11790 & ~n11823 ) ;
  assign n12171 = x122 & n11790 ;
  assign n12172 = ( ~n11795 & n12170 ) | ( ~n11795 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12173 = ( n11795 & n12170 ) | ( n11795 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12174 = ( n11795 & n12172 ) | ( n11795 & ~n12173 ) | ( n12172 & ~n12173 ) ;
  assign n12175 = ( x123 & n12169 ) | ( x123 & ~n12174 ) | ( n12169 & ~n12174 ) ;
  assign n12176 = ( x123 & n11796 ) | ( x123 & ~n11823 ) | ( n11796 & ~n11823 ) ;
  assign n12177 = x123 & n11796 ;
  assign n12178 = ( ~n11801 & n12176 ) | ( ~n11801 & n12177 ) | ( n12176 & n12177 ) ;
  assign n12179 = ( n11801 & n12176 ) | ( n11801 & n12177 ) | ( n12176 & n12177 ) ;
  assign n12180 = ( n11801 & n12178 ) | ( n11801 & ~n12179 ) | ( n12178 & ~n12179 ) ;
  assign n12181 = ( x124 & n12175 ) | ( x124 & ~n12180 ) | ( n12175 & ~n12180 ) ;
  assign n12182 = ( x124 & n11802 ) | ( x124 & ~n11823 ) | ( n11802 & ~n11823 ) ;
  assign n12183 = x124 & n11802 ;
  assign n12184 = ( ~n11807 & n12182 ) | ( ~n11807 & n12183 ) | ( n12182 & n12183 ) ;
  assign n12185 = ( n11807 & n12182 ) | ( n11807 & n12183 ) | ( n12182 & n12183 ) ;
  assign n12186 = ( n11807 & n12184 ) | ( n11807 & ~n12185 ) | ( n12184 & ~n12185 ) ;
  assign n12187 = ( x125 & n12181 ) | ( x125 & ~n12186 ) | ( n12181 & ~n12186 ) ;
  assign n12188 = ( x125 & n11808 ) | ( x125 & ~n11823 ) | ( n11808 & ~n11823 ) ;
  assign n12189 = x125 & n11808 ;
  assign n12190 = ( ~n11813 & n12188 ) | ( ~n11813 & n12189 ) | ( n12188 & n12189 ) ;
  assign n12191 = ( n11813 & n12188 ) | ( n11813 & n12189 ) | ( n12188 & n12189 ) ;
  assign n12192 = ( n11813 & n12190 ) | ( n11813 & ~n12191 ) | ( n12190 & ~n12191 ) ;
  assign n12193 = ( x126 & n12187 ) | ( x126 & ~n12192 ) | ( n12187 & ~n12192 ) ;
  assign n12194 = x127 & ~n11445 ;
  assign n12195 = ~n11817 & n12194 ;
  assign n12196 = ( ~n11817 & n12193 ) | ( ~n11817 & n12195 ) | ( n12193 & n12195 ) ;
  assign n12197 = n192 | n199 ;
  assign n12198 = ~x63 & x64 ;
  assign n12199 = n197 | n12198 ;
  assign n12200 = n190 | n12199 ;
  assign n12201 = x0 & n12196 ;
  assign n12202 = ( x0 & x64 ) | ( x0 & ~n12196 ) | ( x64 & ~n12196 ) ;
  assign n12203 = x0 & x64 ;
  assign n12204 = ( n12201 & n12202 ) | ( n12201 & ~n12203 ) | ( n12202 & ~n12203 ) ;
  assign n12205 = ( x65 & n11818 ) | ( x65 & n12196 ) | ( n11818 & n12196 ) ;
  assign n12206 = x65 | n11818 ;
  assign n12207 = ( ~n11826 & n12205 ) | ( ~n11826 & n12206 ) | ( n12205 & n12206 ) ;
  assign n12208 = ( n11826 & n12205 ) | ( n11826 & n12206 ) | ( n12205 & n12206 ) ;
  assign n12209 = ( n11826 & n12207 ) | ( n11826 & ~n12208 ) | ( n12207 & ~n12208 ) ;
  assign n12210 = ( x66 & n11827 ) | ( x66 & n12196 ) | ( n11827 & n12196 ) ;
  assign n12211 = x66 | n11827 ;
  assign n12212 = ( ~n11832 & n12210 ) | ( ~n11832 & n12211 ) | ( n12210 & n12211 ) ;
  assign n12213 = ( n11832 & n12210 ) | ( n11832 & n12211 ) | ( n12210 & n12211 ) ;
  assign n12214 = ( n11832 & n12212 ) | ( n11832 & ~n12213 ) | ( n12212 & ~n12213 ) ;
  assign n12215 = ( x67 & n11833 ) | ( x67 & ~n12196 ) | ( n11833 & ~n12196 ) ;
  assign n12216 = x67 & n11833 ;
  assign n12217 = ( ~n11838 & n12215 ) | ( ~n11838 & n12216 ) | ( n12215 & n12216 ) ;
  assign n12218 = ( n11838 & n12215 ) | ( n11838 & n12216 ) | ( n12215 & n12216 ) ;
  assign n12219 = ( n11838 & n12217 ) | ( n11838 & ~n12218 ) | ( n12217 & ~n12218 ) ;
  assign n12220 = ( x68 & n11839 ) | ( x68 & ~n12196 ) | ( n11839 & ~n12196 ) ;
  assign n12221 = x68 & n11839 ;
  assign n12222 = ( ~n11844 & n12220 ) | ( ~n11844 & n12221 ) | ( n12220 & n12221 ) ;
  assign n12223 = ( n11844 & n12220 ) | ( n11844 & n12221 ) | ( n12220 & n12221 ) ;
  assign n12224 = ( n11844 & n12222 ) | ( n11844 & ~n12223 ) | ( n12222 & ~n12223 ) ;
  assign n12225 = ( x69 & n11845 ) | ( x69 & ~n12196 ) | ( n11845 & ~n12196 ) ;
  assign n12226 = x69 & n11845 ;
  assign n12227 = ( ~n11850 & n12225 ) | ( ~n11850 & n12226 ) | ( n12225 & n12226 ) ;
  assign n12228 = ( n11850 & n12225 ) | ( n11850 & n12226 ) | ( n12225 & n12226 ) ;
  assign n12229 = ( n11850 & n12227 ) | ( n11850 & ~n12228 ) | ( n12227 & ~n12228 ) ;
  assign n12230 = ( x70 & n11851 ) | ( x70 & ~n12196 ) | ( n11851 & ~n12196 ) ;
  assign n12231 = x70 & n11851 ;
  assign n12232 = ( ~n11856 & n12230 ) | ( ~n11856 & n12231 ) | ( n12230 & n12231 ) ;
  assign n12233 = ( n11856 & n12230 ) | ( n11856 & n12231 ) | ( n12230 & n12231 ) ;
  assign n12234 = ( n11856 & n12232 ) | ( n11856 & ~n12233 ) | ( n12232 & ~n12233 ) ;
  assign n12235 = ( x71 & n11857 ) | ( x71 & ~n12196 ) | ( n11857 & ~n12196 ) ;
  assign n12236 = x71 & n11857 ;
  assign n12237 = ( ~n11862 & n12235 ) | ( ~n11862 & n12236 ) | ( n12235 & n12236 ) ;
  assign n12238 = ( n11862 & n12235 ) | ( n11862 & n12236 ) | ( n12235 & n12236 ) ;
  assign n12239 = ( n11862 & n12237 ) | ( n11862 & ~n12238 ) | ( n12237 & ~n12238 ) ;
  assign n12240 = ( x72 & n11863 ) | ( x72 & ~n12196 ) | ( n11863 & ~n12196 ) ;
  assign n12241 = x72 & n11863 ;
  assign n12242 = ( ~n11868 & n12240 ) | ( ~n11868 & n12241 ) | ( n12240 & n12241 ) ;
  assign n12243 = ( n11868 & n12240 ) | ( n11868 & n12241 ) | ( n12240 & n12241 ) ;
  assign n12244 = ( n11868 & n12242 ) | ( n11868 & ~n12243 ) | ( n12242 & ~n12243 ) ;
  assign n12245 = ( x73 & n11869 ) | ( x73 & ~n12196 ) | ( n11869 & ~n12196 ) ;
  assign n12246 = x73 & n11869 ;
  assign n12247 = ( ~n11874 & n12245 ) | ( ~n11874 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12248 = ( n11874 & n12245 ) | ( n11874 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12249 = ( n11874 & n12247 ) | ( n11874 & ~n12248 ) | ( n12247 & ~n12248 ) ;
  assign n12250 = ( x74 & n11875 ) | ( x74 & ~n12196 ) | ( n11875 & ~n12196 ) ;
  assign n12251 = x74 & n11875 ;
  assign n12252 = ( ~n11880 & n12250 ) | ( ~n11880 & n12251 ) | ( n12250 & n12251 ) ;
  assign n12253 = ( n11880 & n12250 ) | ( n11880 & n12251 ) | ( n12250 & n12251 ) ;
  assign n12254 = ( n11880 & n12252 ) | ( n11880 & ~n12253 ) | ( n12252 & ~n12253 ) ;
  assign n12255 = ( x75 & n11881 ) | ( x75 & ~n12196 ) | ( n11881 & ~n12196 ) ;
  assign n12256 = x75 & n11881 ;
  assign n12257 = ( ~n11886 & n12255 ) | ( ~n11886 & n12256 ) | ( n12255 & n12256 ) ;
  assign n12258 = ( n11886 & n12255 ) | ( n11886 & n12256 ) | ( n12255 & n12256 ) ;
  assign n12259 = ( n11886 & n12257 ) | ( n11886 & ~n12258 ) | ( n12257 & ~n12258 ) ;
  assign n12260 = ( x76 & n11887 ) | ( x76 & ~n12196 ) | ( n11887 & ~n12196 ) ;
  assign n12261 = x76 & n11887 ;
  assign n12262 = ( ~n11892 & n12260 ) | ( ~n11892 & n12261 ) | ( n12260 & n12261 ) ;
  assign n12263 = ( n11892 & n12260 ) | ( n11892 & n12261 ) | ( n12260 & n12261 ) ;
  assign n12264 = ( n11892 & n12262 ) | ( n11892 & ~n12263 ) | ( n12262 & ~n12263 ) ;
  assign n12265 = ( x77 & n11893 ) | ( x77 & ~n12196 ) | ( n11893 & ~n12196 ) ;
  assign n12266 = x77 & n11893 ;
  assign n12267 = ( ~n11898 & n12265 ) | ( ~n11898 & n12266 ) | ( n12265 & n12266 ) ;
  assign n12268 = ( n11898 & n12265 ) | ( n11898 & n12266 ) | ( n12265 & n12266 ) ;
  assign n12269 = ( n11898 & n12267 ) | ( n11898 & ~n12268 ) | ( n12267 & ~n12268 ) ;
  assign n12270 = ( x78 & n11899 ) | ( x78 & ~n12196 ) | ( n11899 & ~n12196 ) ;
  assign n12271 = x78 & n11899 ;
  assign n12272 = ( ~n11904 & n12270 ) | ( ~n11904 & n12271 ) | ( n12270 & n12271 ) ;
  assign n12273 = ( n11904 & n12270 ) | ( n11904 & n12271 ) | ( n12270 & n12271 ) ;
  assign n12274 = ( n11904 & n12272 ) | ( n11904 & ~n12273 ) | ( n12272 & ~n12273 ) ;
  assign n12275 = ( x79 & n11905 ) | ( x79 & ~n12196 ) | ( n11905 & ~n12196 ) ;
  assign n12276 = x79 & n11905 ;
  assign n12277 = ( ~n11910 & n12275 ) | ( ~n11910 & n12276 ) | ( n12275 & n12276 ) ;
  assign n12278 = ( n11910 & n12275 ) | ( n11910 & n12276 ) | ( n12275 & n12276 ) ;
  assign n12279 = ( n11910 & n12277 ) | ( n11910 & ~n12278 ) | ( n12277 & ~n12278 ) ;
  assign n12280 = ( x80 & n11911 ) | ( x80 & ~n12196 ) | ( n11911 & ~n12196 ) ;
  assign n12281 = x80 & n11911 ;
  assign n12282 = ( ~n11916 & n12280 ) | ( ~n11916 & n12281 ) | ( n12280 & n12281 ) ;
  assign n12283 = ( n11916 & n12280 ) | ( n11916 & n12281 ) | ( n12280 & n12281 ) ;
  assign n12284 = ( n11916 & n12282 ) | ( n11916 & ~n12283 ) | ( n12282 & ~n12283 ) ;
  assign n12285 = ( x81 & n11917 ) | ( x81 & ~n12196 ) | ( n11917 & ~n12196 ) ;
  assign n12286 = x81 & n11917 ;
  assign n12287 = ( ~n11922 & n12285 ) | ( ~n11922 & n12286 ) | ( n12285 & n12286 ) ;
  assign n12288 = ( n11922 & n12285 ) | ( n11922 & n12286 ) | ( n12285 & n12286 ) ;
  assign n12289 = ( n11922 & n12287 ) | ( n11922 & ~n12288 ) | ( n12287 & ~n12288 ) ;
  assign n12290 = ( x82 & n11923 ) | ( x82 & ~n12196 ) | ( n11923 & ~n12196 ) ;
  assign n12291 = x82 & n11923 ;
  assign n12292 = ( ~n11928 & n12290 ) | ( ~n11928 & n12291 ) | ( n12290 & n12291 ) ;
  assign n12293 = ( n11928 & n12290 ) | ( n11928 & n12291 ) | ( n12290 & n12291 ) ;
  assign n12294 = ( n11928 & n12292 ) | ( n11928 & ~n12293 ) | ( n12292 & ~n12293 ) ;
  assign n12295 = ( x83 & n11929 ) | ( x83 & ~n12196 ) | ( n11929 & ~n12196 ) ;
  assign n12296 = x83 & n11929 ;
  assign n12297 = ( ~n11934 & n12295 ) | ( ~n11934 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12298 = ( n11934 & n12295 ) | ( n11934 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12299 = ( n11934 & n12297 ) | ( n11934 & ~n12298 ) | ( n12297 & ~n12298 ) ;
  assign n12300 = ( x84 & n11935 ) | ( x84 & ~n12196 ) | ( n11935 & ~n12196 ) ;
  assign n12301 = x84 & n11935 ;
  assign n12302 = ( ~n11940 & n12300 ) | ( ~n11940 & n12301 ) | ( n12300 & n12301 ) ;
  assign n12303 = ( n11940 & n12300 ) | ( n11940 & n12301 ) | ( n12300 & n12301 ) ;
  assign n12304 = ( n11940 & n12302 ) | ( n11940 & ~n12303 ) | ( n12302 & ~n12303 ) ;
  assign n12305 = ( x85 & n11941 ) | ( x85 & ~n12196 ) | ( n11941 & ~n12196 ) ;
  assign n12306 = x85 & n11941 ;
  assign n12307 = ( ~n11946 & n12305 ) | ( ~n11946 & n12306 ) | ( n12305 & n12306 ) ;
  assign n12308 = ( n11946 & n12305 ) | ( n11946 & n12306 ) | ( n12305 & n12306 ) ;
  assign n12309 = ( n11946 & n12307 ) | ( n11946 & ~n12308 ) | ( n12307 & ~n12308 ) ;
  assign n12310 = ( x86 & n11947 ) | ( x86 & ~n12196 ) | ( n11947 & ~n12196 ) ;
  assign n12311 = x86 & n11947 ;
  assign n12312 = ( ~n11952 & n12310 ) | ( ~n11952 & n12311 ) | ( n12310 & n12311 ) ;
  assign n12313 = ( n11952 & n12310 ) | ( n11952 & n12311 ) | ( n12310 & n12311 ) ;
  assign n12314 = ( n11952 & n12312 ) | ( n11952 & ~n12313 ) | ( n12312 & ~n12313 ) ;
  assign n12315 = ( x87 & n11953 ) | ( x87 & ~n12196 ) | ( n11953 & ~n12196 ) ;
  assign n12316 = x87 & n11953 ;
  assign n12317 = ( ~n11958 & n12315 ) | ( ~n11958 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12318 = ( n11958 & n12315 ) | ( n11958 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12319 = ( n11958 & n12317 ) | ( n11958 & ~n12318 ) | ( n12317 & ~n12318 ) ;
  assign n12320 = ( x88 & n11959 ) | ( x88 & ~n12196 ) | ( n11959 & ~n12196 ) ;
  assign n12321 = x88 & n11959 ;
  assign n12322 = ( ~n11964 & n12320 ) | ( ~n11964 & n12321 ) | ( n12320 & n12321 ) ;
  assign n12323 = ( n11964 & n12320 ) | ( n11964 & n12321 ) | ( n12320 & n12321 ) ;
  assign n12324 = ( n11964 & n12322 ) | ( n11964 & ~n12323 ) | ( n12322 & ~n12323 ) ;
  assign n12325 = ( x89 & n11965 ) | ( x89 & ~n12196 ) | ( n11965 & ~n12196 ) ;
  assign n12326 = x89 & n11965 ;
  assign n12327 = ( ~n11970 & n12325 ) | ( ~n11970 & n12326 ) | ( n12325 & n12326 ) ;
  assign n12328 = ( n11970 & n12325 ) | ( n11970 & n12326 ) | ( n12325 & n12326 ) ;
  assign n12329 = ( n11970 & n12327 ) | ( n11970 & ~n12328 ) | ( n12327 & ~n12328 ) ;
  assign n12330 = ( x90 & n11971 ) | ( x90 & ~n12196 ) | ( n11971 & ~n12196 ) ;
  assign n12331 = x90 & n11971 ;
  assign n12332 = ( ~n11976 & n12330 ) | ( ~n11976 & n12331 ) | ( n12330 & n12331 ) ;
  assign n12333 = ( n11976 & n12330 ) | ( n11976 & n12331 ) | ( n12330 & n12331 ) ;
  assign n12334 = ( n11976 & n12332 ) | ( n11976 & ~n12333 ) | ( n12332 & ~n12333 ) ;
  assign n12335 = ( x91 & n11977 ) | ( x91 & ~n12196 ) | ( n11977 & ~n12196 ) ;
  assign n12336 = x91 & n11977 ;
  assign n12337 = ( ~n11982 & n12335 ) | ( ~n11982 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12338 = ( n11982 & n12335 ) | ( n11982 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12339 = ( n11982 & n12337 ) | ( n11982 & ~n12338 ) | ( n12337 & ~n12338 ) ;
  assign n12340 = ( x92 & n11983 ) | ( x92 & ~n12196 ) | ( n11983 & ~n12196 ) ;
  assign n12341 = x92 & n11983 ;
  assign n12342 = ( ~n11988 & n12340 ) | ( ~n11988 & n12341 ) | ( n12340 & n12341 ) ;
  assign n12343 = ( n11988 & n12340 ) | ( n11988 & n12341 ) | ( n12340 & n12341 ) ;
  assign n12344 = ( n11988 & n12342 ) | ( n11988 & ~n12343 ) | ( n12342 & ~n12343 ) ;
  assign n12345 = ( x93 & n11989 ) | ( x93 & ~n12196 ) | ( n11989 & ~n12196 ) ;
  assign n12346 = x93 & n11989 ;
  assign n12347 = ( ~n11994 & n12345 ) | ( ~n11994 & n12346 ) | ( n12345 & n12346 ) ;
  assign n12348 = ( n11994 & n12345 ) | ( n11994 & n12346 ) | ( n12345 & n12346 ) ;
  assign n12349 = ( n11994 & n12347 ) | ( n11994 & ~n12348 ) | ( n12347 & ~n12348 ) ;
  assign n12350 = ( x94 & n11995 ) | ( x94 & ~n12196 ) | ( n11995 & ~n12196 ) ;
  assign n12351 = x94 & n11995 ;
  assign n12352 = ( ~n12000 & n12350 ) | ( ~n12000 & n12351 ) | ( n12350 & n12351 ) ;
  assign n12353 = ( n12000 & n12350 ) | ( n12000 & n12351 ) | ( n12350 & n12351 ) ;
  assign n12354 = ( n12000 & n12352 ) | ( n12000 & ~n12353 ) | ( n12352 & ~n12353 ) ;
  assign n12355 = ( x95 & n12001 ) | ( x95 & ~n12196 ) | ( n12001 & ~n12196 ) ;
  assign n12356 = x95 & n12001 ;
  assign n12357 = ( ~n12006 & n12355 ) | ( ~n12006 & n12356 ) | ( n12355 & n12356 ) ;
  assign n12358 = ( n12006 & n12355 ) | ( n12006 & n12356 ) | ( n12355 & n12356 ) ;
  assign n12359 = ( n12006 & n12357 ) | ( n12006 & ~n12358 ) | ( n12357 & ~n12358 ) ;
  assign n12360 = ( x96 & n12007 ) | ( x96 & ~n12196 ) | ( n12007 & ~n12196 ) ;
  assign n12361 = x96 & n12007 ;
  assign n12362 = ( ~n12012 & n12360 ) | ( ~n12012 & n12361 ) | ( n12360 & n12361 ) ;
  assign n12363 = ( n12012 & n12360 ) | ( n12012 & n12361 ) | ( n12360 & n12361 ) ;
  assign n12364 = ( n12012 & n12362 ) | ( n12012 & ~n12363 ) | ( n12362 & ~n12363 ) ;
  assign n12365 = ( x97 & n12013 ) | ( x97 & ~n12196 ) | ( n12013 & ~n12196 ) ;
  assign n12366 = x97 & n12013 ;
  assign n12367 = ( ~n12018 & n12365 ) | ( ~n12018 & n12366 ) | ( n12365 & n12366 ) ;
  assign n12368 = ( n12018 & n12365 ) | ( n12018 & n12366 ) | ( n12365 & n12366 ) ;
  assign n12369 = ( n12018 & n12367 ) | ( n12018 & ~n12368 ) | ( n12367 & ~n12368 ) ;
  assign n12370 = ( x98 & n12019 ) | ( x98 & ~n12196 ) | ( n12019 & ~n12196 ) ;
  assign n12371 = x98 & n12019 ;
  assign n12372 = ( ~n12024 & n12370 ) | ( ~n12024 & n12371 ) | ( n12370 & n12371 ) ;
  assign n12373 = ( n12024 & n12370 ) | ( n12024 & n12371 ) | ( n12370 & n12371 ) ;
  assign n12374 = ( n12024 & n12372 ) | ( n12024 & ~n12373 ) | ( n12372 & ~n12373 ) ;
  assign n12375 = ( x99 & n12025 ) | ( x99 & ~n12196 ) | ( n12025 & ~n12196 ) ;
  assign n12376 = x99 & n12025 ;
  assign n12377 = ( ~n12030 & n12375 ) | ( ~n12030 & n12376 ) | ( n12375 & n12376 ) ;
  assign n12378 = ( n12030 & n12375 ) | ( n12030 & n12376 ) | ( n12375 & n12376 ) ;
  assign n12379 = ( n12030 & n12377 ) | ( n12030 & ~n12378 ) | ( n12377 & ~n12378 ) ;
  assign n12380 = ( x100 & n12031 ) | ( x100 & ~n12196 ) | ( n12031 & ~n12196 ) ;
  assign n12381 = x100 & n12031 ;
  assign n12382 = ( ~n12036 & n12380 ) | ( ~n12036 & n12381 ) | ( n12380 & n12381 ) ;
  assign n12383 = ( n12036 & n12380 ) | ( n12036 & n12381 ) | ( n12380 & n12381 ) ;
  assign n12384 = ( n12036 & n12382 ) | ( n12036 & ~n12383 ) | ( n12382 & ~n12383 ) ;
  assign n12385 = ( x101 & n12037 ) | ( x101 & ~n12196 ) | ( n12037 & ~n12196 ) ;
  assign n12386 = x101 & n12037 ;
  assign n12387 = ( ~n12042 & n12385 ) | ( ~n12042 & n12386 ) | ( n12385 & n12386 ) ;
  assign n12388 = ( n12042 & n12385 ) | ( n12042 & n12386 ) | ( n12385 & n12386 ) ;
  assign n12389 = ( n12042 & n12387 ) | ( n12042 & ~n12388 ) | ( n12387 & ~n12388 ) ;
  assign n12390 = ( x102 & n12043 ) | ( x102 & ~n12196 ) | ( n12043 & ~n12196 ) ;
  assign n12391 = x102 & n12043 ;
  assign n12392 = ( ~n12048 & n12390 ) | ( ~n12048 & n12391 ) | ( n12390 & n12391 ) ;
  assign n12393 = ( n12048 & n12390 ) | ( n12048 & n12391 ) | ( n12390 & n12391 ) ;
  assign n12394 = ( n12048 & n12392 ) | ( n12048 & ~n12393 ) | ( n12392 & ~n12393 ) ;
  assign n12395 = ( x103 & n12049 ) | ( x103 & ~n12196 ) | ( n12049 & ~n12196 ) ;
  assign n12396 = x103 & n12049 ;
  assign n12397 = ( ~n12054 & n12395 ) | ( ~n12054 & n12396 ) | ( n12395 & n12396 ) ;
  assign n12398 = ( n12054 & n12395 ) | ( n12054 & n12396 ) | ( n12395 & n12396 ) ;
  assign n12399 = ( n12054 & n12397 ) | ( n12054 & ~n12398 ) | ( n12397 & ~n12398 ) ;
  assign n12400 = ( x104 & n12055 ) | ( x104 & ~n12196 ) | ( n12055 & ~n12196 ) ;
  assign n12401 = x104 & n12055 ;
  assign n12402 = ( ~n12060 & n12400 ) | ( ~n12060 & n12401 ) | ( n12400 & n12401 ) ;
  assign n12403 = ( n12060 & n12400 ) | ( n12060 & n12401 ) | ( n12400 & n12401 ) ;
  assign n12404 = ( n12060 & n12402 ) | ( n12060 & ~n12403 ) | ( n12402 & ~n12403 ) ;
  assign n12405 = ( x105 & n12061 ) | ( x105 & ~n12196 ) | ( n12061 & ~n12196 ) ;
  assign n12406 = x105 & n12061 ;
  assign n12407 = ( ~n12066 & n12405 ) | ( ~n12066 & n12406 ) | ( n12405 & n12406 ) ;
  assign n12408 = ( n12066 & n12405 ) | ( n12066 & n12406 ) | ( n12405 & n12406 ) ;
  assign n12409 = ( n12066 & n12407 ) | ( n12066 & ~n12408 ) | ( n12407 & ~n12408 ) ;
  assign n12410 = ( x106 & n12067 ) | ( x106 & ~n12196 ) | ( n12067 & ~n12196 ) ;
  assign n12411 = x106 & n12067 ;
  assign n12412 = ( ~n12072 & n12410 ) | ( ~n12072 & n12411 ) | ( n12410 & n12411 ) ;
  assign n12413 = ( n12072 & n12410 ) | ( n12072 & n12411 ) | ( n12410 & n12411 ) ;
  assign n12414 = ( n12072 & n12412 ) | ( n12072 & ~n12413 ) | ( n12412 & ~n12413 ) ;
  assign n12415 = ( x107 & n12073 ) | ( x107 & ~n12196 ) | ( n12073 & ~n12196 ) ;
  assign n12416 = x107 & n12073 ;
  assign n12417 = ( ~n12078 & n12415 ) | ( ~n12078 & n12416 ) | ( n12415 & n12416 ) ;
  assign n12418 = ( n12078 & n12415 ) | ( n12078 & n12416 ) | ( n12415 & n12416 ) ;
  assign n12419 = ( n12078 & n12417 ) | ( n12078 & ~n12418 ) | ( n12417 & ~n12418 ) ;
  assign n12420 = ( x108 & n12079 ) | ( x108 & ~n12196 ) | ( n12079 & ~n12196 ) ;
  assign n12421 = x108 & n12079 ;
  assign n12422 = ( ~n12084 & n12420 ) | ( ~n12084 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12423 = ( n12084 & n12420 ) | ( n12084 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12424 = ( n12084 & n12422 ) | ( n12084 & ~n12423 ) | ( n12422 & ~n12423 ) ;
  assign n12425 = ( x109 & n12085 ) | ( x109 & ~n12196 ) | ( n12085 & ~n12196 ) ;
  assign n12426 = x109 & n12085 ;
  assign n12427 = ( ~n12090 & n12425 ) | ( ~n12090 & n12426 ) | ( n12425 & n12426 ) ;
  assign n12428 = ( n12090 & n12425 ) | ( n12090 & n12426 ) | ( n12425 & n12426 ) ;
  assign n12429 = ( n12090 & n12427 ) | ( n12090 & ~n12428 ) | ( n12427 & ~n12428 ) ;
  assign n12430 = ( x110 & n12091 ) | ( x110 & ~n12196 ) | ( n12091 & ~n12196 ) ;
  assign n12431 = x110 & n12091 ;
  assign n12432 = ( ~n12096 & n12430 ) | ( ~n12096 & n12431 ) | ( n12430 & n12431 ) ;
  assign n12433 = ( n12096 & n12430 ) | ( n12096 & n12431 ) | ( n12430 & n12431 ) ;
  assign n12434 = ( n12096 & n12432 ) | ( n12096 & ~n12433 ) | ( n12432 & ~n12433 ) ;
  assign n12435 = ( x111 & n12097 ) | ( x111 & ~n12196 ) | ( n12097 & ~n12196 ) ;
  assign n12436 = x111 & n12097 ;
  assign n12437 = ( ~n12102 & n12435 ) | ( ~n12102 & n12436 ) | ( n12435 & n12436 ) ;
  assign n12438 = ( n12102 & n12435 ) | ( n12102 & n12436 ) | ( n12435 & n12436 ) ;
  assign n12439 = ( n12102 & n12437 ) | ( n12102 & ~n12438 ) | ( n12437 & ~n12438 ) ;
  assign n12440 = ( x112 & n12103 ) | ( x112 & ~n12196 ) | ( n12103 & ~n12196 ) ;
  assign n12441 = x112 & n12103 ;
  assign n12442 = ( ~n12108 & n12440 ) | ( ~n12108 & n12441 ) | ( n12440 & n12441 ) ;
  assign n12443 = ( n12108 & n12440 ) | ( n12108 & n12441 ) | ( n12440 & n12441 ) ;
  assign n12444 = ( n12108 & n12442 ) | ( n12108 & ~n12443 ) | ( n12442 & ~n12443 ) ;
  assign n12445 = ( x113 & n12109 ) | ( x113 & ~n12196 ) | ( n12109 & ~n12196 ) ;
  assign n12446 = x113 & n12109 ;
  assign n12447 = ( ~n12114 & n12445 ) | ( ~n12114 & n12446 ) | ( n12445 & n12446 ) ;
  assign n12448 = ( n12114 & n12445 ) | ( n12114 & n12446 ) | ( n12445 & n12446 ) ;
  assign n12449 = ( n12114 & n12447 ) | ( n12114 & ~n12448 ) | ( n12447 & ~n12448 ) ;
  assign n12450 = ( x114 & n12115 ) | ( x114 & ~n12196 ) | ( n12115 & ~n12196 ) ;
  assign n12451 = x114 & n12115 ;
  assign n12452 = ( ~n12120 & n12450 ) | ( ~n12120 & n12451 ) | ( n12450 & n12451 ) ;
  assign n12453 = ( n12120 & n12450 ) | ( n12120 & n12451 ) | ( n12450 & n12451 ) ;
  assign n12454 = ( n12120 & n12452 ) | ( n12120 & ~n12453 ) | ( n12452 & ~n12453 ) ;
  assign n12455 = ( x115 & n12121 ) | ( x115 & ~n12196 ) | ( n12121 & ~n12196 ) ;
  assign n12456 = x115 & n12121 ;
  assign n12457 = ( ~n12126 & n12455 ) | ( ~n12126 & n12456 ) | ( n12455 & n12456 ) ;
  assign n12458 = ( n12126 & n12455 ) | ( n12126 & n12456 ) | ( n12455 & n12456 ) ;
  assign n12459 = ( n12126 & n12457 ) | ( n12126 & ~n12458 ) | ( n12457 & ~n12458 ) ;
  assign n12460 = ( x116 & n12127 ) | ( x116 & ~n12196 ) | ( n12127 & ~n12196 ) ;
  assign n12461 = x116 & n12127 ;
  assign n12462 = ( ~n12132 & n12460 ) | ( ~n12132 & n12461 ) | ( n12460 & n12461 ) ;
  assign n12463 = ( n12132 & n12460 ) | ( n12132 & n12461 ) | ( n12460 & n12461 ) ;
  assign n12464 = ( n12132 & n12462 ) | ( n12132 & ~n12463 ) | ( n12462 & ~n12463 ) ;
  assign n12465 = ( x117 & n12133 ) | ( x117 & ~n12196 ) | ( n12133 & ~n12196 ) ;
  assign n12466 = x117 & n12133 ;
  assign n12467 = ( ~n12138 & n12465 ) | ( ~n12138 & n12466 ) | ( n12465 & n12466 ) ;
  assign n12468 = ( n12138 & n12465 ) | ( n12138 & n12466 ) | ( n12465 & n12466 ) ;
  assign n12469 = ( n12138 & n12467 ) | ( n12138 & ~n12468 ) | ( n12467 & ~n12468 ) ;
  assign n12470 = ( x118 & n12139 ) | ( x118 & ~n12196 ) | ( n12139 & ~n12196 ) ;
  assign n12471 = x118 & n12139 ;
  assign n12472 = ( ~n12144 & n12470 ) | ( ~n12144 & n12471 ) | ( n12470 & n12471 ) ;
  assign n12473 = ( n12144 & n12470 ) | ( n12144 & n12471 ) | ( n12470 & n12471 ) ;
  assign n12474 = ( n12144 & n12472 ) | ( n12144 & ~n12473 ) | ( n12472 & ~n12473 ) ;
  assign n12475 = ( x119 & n12145 ) | ( x119 & ~n12196 ) | ( n12145 & ~n12196 ) ;
  assign n12476 = x119 & n12145 ;
  assign n12477 = ( ~n12150 & n12475 ) | ( ~n12150 & n12476 ) | ( n12475 & n12476 ) ;
  assign n12478 = ( n12150 & n12475 ) | ( n12150 & n12476 ) | ( n12475 & n12476 ) ;
  assign n12479 = ( n12150 & n12477 ) | ( n12150 & ~n12478 ) | ( n12477 & ~n12478 ) ;
  assign n12480 = ( x120 & n12151 ) | ( x120 & ~n12196 ) | ( n12151 & ~n12196 ) ;
  assign n12481 = x120 & n12151 ;
  assign n12482 = ( ~n12156 & n12480 ) | ( ~n12156 & n12481 ) | ( n12480 & n12481 ) ;
  assign n12483 = ( n12156 & n12480 ) | ( n12156 & n12481 ) | ( n12480 & n12481 ) ;
  assign n12484 = ( n12156 & n12482 ) | ( n12156 & ~n12483 ) | ( n12482 & ~n12483 ) ;
  assign n12485 = ( x121 & n12157 ) | ( x121 & ~n12196 ) | ( n12157 & ~n12196 ) ;
  assign n12486 = x121 & n12157 ;
  assign n12487 = ( ~n12162 & n12485 ) | ( ~n12162 & n12486 ) | ( n12485 & n12486 ) ;
  assign n12488 = ( n12162 & n12485 ) | ( n12162 & n12486 ) | ( n12485 & n12486 ) ;
  assign n12489 = ( n12162 & n12487 ) | ( n12162 & ~n12488 ) | ( n12487 & ~n12488 ) ;
  assign n12490 = ( x122 & n12163 ) | ( x122 & ~n12196 ) | ( n12163 & ~n12196 ) ;
  assign n12491 = x122 & n12163 ;
  assign n12492 = ( ~n12168 & n12490 ) | ( ~n12168 & n12491 ) | ( n12490 & n12491 ) ;
  assign n12493 = ( n12168 & n12490 ) | ( n12168 & n12491 ) | ( n12490 & n12491 ) ;
  assign n12494 = ( n12168 & n12492 ) | ( n12168 & ~n12493 ) | ( n12492 & ~n12493 ) ;
  assign n12495 = ( x123 & n12169 ) | ( x123 & ~n12196 ) | ( n12169 & ~n12196 ) ;
  assign n12496 = x123 & n12169 ;
  assign n12497 = ( ~n12174 & n12495 ) | ( ~n12174 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12498 = ( n12174 & n12495 ) | ( n12174 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12499 = ( n12174 & n12497 ) | ( n12174 & ~n12498 ) | ( n12497 & ~n12498 ) ;
  assign n12500 = ( x124 & n12175 ) | ( x124 & ~n12196 ) | ( n12175 & ~n12196 ) ;
  assign n12501 = x124 & n12175 ;
  assign n12502 = ( ~n12180 & n12500 ) | ( ~n12180 & n12501 ) | ( n12500 & n12501 ) ;
  assign n12503 = ( n12180 & n12500 ) | ( n12180 & n12501 ) | ( n12500 & n12501 ) ;
  assign n12504 = ( n12180 & n12502 ) | ( n12180 & ~n12503 ) | ( n12502 & ~n12503 ) ;
  assign n12505 = ( x125 & n12181 ) | ( x125 & ~n12196 ) | ( n12181 & ~n12196 ) ;
  assign n12506 = x125 & n12181 ;
  assign n12507 = ( ~n12186 & n12505 ) | ( ~n12186 & n12506 ) | ( n12505 & n12506 ) ;
  assign n12508 = ( n12186 & n12505 ) | ( n12186 & n12506 ) | ( n12505 & n12506 ) ;
  assign n12509 = ( n12186 & n12507 ) | ( n12186 & ~n12508 ) | ( n12507 & ~n12508 ) ;
  assign n12510 = ( x126 & n12187 ) | ( x126 & ~n12196 ) | ( n12187 & ~n12196 ) ;
  assign n12511 = x126 & n12187 ;
  assign n12512 = ( ~n12192 & n12510 ) | ( ~n12192 & n12511 ) | ( n12510 & n12511 ) ;
  assign n12513 = ( n12192 & n12510 ) | ( n12192 & n12511 ) | ( n12510 & n12511 ) ;
  assign n12514 = ( n12192 & n12512 ) | ( n12192 & ~n12513 ) | ( n12512 & ~n12513 ) ;
  assign n12515 = ( x127 & n389 ) | ( x127 & n11445 ) | ( n389 & n11445 ) ;
  assign n12516 = ( n389 & n12193 ) | ( n389 & n12515 ) | ( n12193 & n12515 ) ;
  assign y0 = ~n12196 ;
  assign y1 = ~n11823 ;
  assign y2 = ~n11450 ;
  assign y3 = ~n11083 ;
  assign y4 = ~n10724 ;
  assign y5 = ~n10371 ;
  assign y6 = ~n10024 ;
  assign y7 = ~n9681 ;
  assign y8 = ~n9347 ;
  assign y9 = ~n9019 ;
  assign y10 = ~n8697 ;
  assign y11 = ~n8381 ;
  assign y12 = ~n8071 ;
  assign y13 = ~n7767 ;
  assign y14 = ~n7470 ;
  assign y15 = ~n7177 ;
  assign y16 = ~n6892 ;
  assign y17 = ~n6610 ;
  assign y18 = ~n6336 ;
  assign y19 = ~n6068 ;
  assign y20 = ~n5806 ;
  assign y21 = ~n5550 ;
  assign y22 = ~n5299 ;
  assign y23 = ~n5054 ;
  assign y24 = ~n4816 ;
  assign y25 = ~n4582 ;
  assign y26 = ~n4354 ;
  assign y27 = ~n4134 ;
  assign y28 = ~n3920 ;
  assign y29 = ~n3711 ;
  assign y30 = ~n3509 ;
  assign y31 = ~n3312 ;
  assign y32 = ~n3121 ;
  assign y33 = ~n2937 ;
  assign y34 = ~n2757 ;
  assign y35 = ~n2584 ;
  assign y36 = ~n2418 ;
  assign y37 = ~n2257 ;
  assign y38 = ~n2101 ;
  assign y39 = ~n1953 ;
  assign y40 = ~n1812 ;
  assign y41 = ~n1674 ;
  assign y42 = ~n1544 ;
  assign y43 = ~n1419 ;
  assign y44 = ~n1300 ;
  assign y45 = ~n1188 ;
  assign y46 = ~n1080 ;
  assign y47 = ~n979 ;
  assign y48 = ~n885 ;
  assign y49 = ~n797 ;
  assign y50 = ~n714 ;
  assign y51 = ~n638 ;
  assign y52 = ~n568 ;
  assign y53 = ~n503 ;
  assign y54 = ~n445 ;
  assign y55 = ~n393 ;
  assign y56 = ~n348 ;
  assign y57 = ~n305 ;
  assign y58 = ~n275 ;
  assign y59 = ~n248 ;
  assign y60 = ~n226 ;
  assign y61 = ~n205 ;
  assign y62 = ~n12197 ;
  assign y63 = ~n12200 ;
  assign y64 = n12204 ;
  assign y65 = n12209 ;
  assign y66 = n12214 ;
  assign y67 = n12219 ;
  assign y68 = n12224 ;
  assign y69 = n12229 ;
  assign y70 = n12234 ;
  assign y71 = n12239 ;
  assign y72 = n12244 ;
  assign y73 = n12249 ;
  assign y74 = n12254 ;
  assign y75 = n12259 ;
  assign y76 = n12264 ;
  assign y77 = n12269 ;
  assign y78 = n12274 ;
  assign y79 = n12279 ;
  assign y80 = n12284 ;
  assign y81 = n12289 ;
  assign y82 = n12294 ;
  assign y83 = n12299 ;
  assign y84 = n12304 ;
  assign y85 = n12309 ;
  assign y86 = n12314 ;
  assign y87 = n12319 ;
  assign y88 = n12324 ;
  assign y89 = n12329 ;
  assign y90 = n12334 ;
  assign y91 = n12339 ;
  assign y92 = n12344 ;
  assign y93 = n12349 ;
  assign y94 = n12354 ;
  assign y95 = n12359 ;
  assign y96 = n12364 ;
  assign y97 = n12369 ;
  assign y98 = n12374 ;
  assign y99 = n12379 ;
  assign y100 = n12384 ;
  assign y101 = n12389 ;
  assign y102 = n12394 ;
  assign y103 = n12399 ;
  assign y104 = n12404 ;
  assign y105 = n12409 ;
  assign y106 = n12414 ;
  assign y107 = n12419 ;
  assign y108 = n12424 ;
  assign y109 = n12429 ;
  assign y110 = n12434 ;
  assign y111 = n12439 ;
  assign y112 = n12444 ;
  assign y113 = n12449 ;
  assign y114 = n12454 ;
  assign y115 = n12459 ;
  assign y116 = n12464 ;
  assign y117 = n12469 ;
  assign y118 = n12474 ;
  assign y119 = n12479 ;
  assign y120 = n12484 ;
  assign y121 = n12489 ;
  assign y122 = n12494 ;
  assign y123 = n12499 ;
  assign y124 = n12504 ;
  assign y125 = n12509 ;
  assign y126 = n12514 ;
  assign y127 = n12516 ;
endmodule
